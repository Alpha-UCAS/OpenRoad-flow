module MyMem( // @[:@2236.2]
  input         clock, // @[:@2237.4]
  input         io_wen, // @[:@2239.4]
  input  [5:0]  io_addr, // @[:@2239.4]
  input  [31:0] io_wdata, // @[:@2239.4]
  output [31:0] io_rdata // @[:@2239.4]
);
  reg [31:0] mem [0:63]; // @[CaheCore.scala 16:24:@2241.4]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_15_data; // @[CaheCore.scala 16:24:@2241.4]
  wire [5:0] mem__T_15_addr; // @[CaheCore.scala 16:24:@2241.4]
  wire [31:0] mem__T_16_data; // @[CaheCore.scala 16:24:@2241.4]
  wire [5:0] mem__T_16_addr; // @[CaheCore.scala 16:24:@2241.4]
  wire  mem__T_16_mask; // @[CaheCore.scala 16:24:@2241.4]
  wire  mem__T_16_en; // @[CaheCore.scala 16:24:@2241.4]
  wire  _GEN_3; // @[CaheCore.scala 18:17:@2244.4]
  reg [5:0] mem__T_15_addr_pipe_0;
  reg [31:0] _RAND_1;
  assign mem__T_15_addr = mem__T_15_addr_pipe_0;
  assign mem__T_15_data = mem[mem__T_15_addr]; // @[CaheCore.scala 16:24:@2241.4]
  assign mem__T_16_data = io_wdata;
  assign mem__T_16_addr = io_addr;
  assign mem__T_16_mask = 1'h1;
  assign mem__T_16_en = io_wen;
  assign _GEN_3 = 1'h1; // @[CaheCore.scala 18:17:@2244.4]
  assign io_rdata = mem__T_15_data; // @[CaheCore.scala 17:12:@2243.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_15_addr_pipe_0 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_16_en & mem__T_16_mask) begin
      mem[mem__T_16_addr] <= mem__T_16_data; // @[CaheCore.scala 16:24:@2241.4]
    end
    if (_GEN_3) begin
      mem__T_15_addr_pipe_0 <= io_addr;
    end
  end
endmodule
module CaheCore( // @[:@2444.2]
  input         clock, // @[:@2445.4]
  input         reset, // @[:@2446.4]
  input         io_wen, // @[:@2447.4]
  input  [31:0] io_addr, // @[:@2447.4]
  input  [31:0] io_wdata_0, // @[:@2447.4]
  input  [31:0] io_wdata_1, // @[:@2447.4]
  input  [31:0] io_wdata_2, // @[:@2447.4]
  input  [31:0] io_wdata_3, // @[:@2447.4]
  input  [31:0] io_wdata_4, // @[:@2447.4]
  input  [31:0] io_wdata_5, // @[:@2447.4]
  input  [31:0] io_wdata_6, // @[:@2447.4]
  input  [31:0] io_wdata_7, // @[:@2447.4]
  input  [31:0] io_wdata_8, // @[:@2447.4]
  input  [31:0] io_wdata_9, // @[:@2447.4]
  input  [31:0] io_wdata_10, // @[:@2447.4]
  input  [31:0] io_wdata_11, // @[:@2447.4]
  input  [31:0] io_wdata_12, // @[:@2447.4]
  input  [31:0] io_wdata_13, // @[:@2447.4]
  input  [31:0] io_wdata_14, // @[:@2447.4]
  input  [31:0] io_wdata_15, // @[:@2447.4]
  input         io_wstatus, // @[:@2447.4]
  output [31:0] io_rdata, // @[:@2447.4]
  output        io_rvalid // @[:@2447.4]
);
  wire  MyMem_clock; // @[CaheCore.scala 34:43:@2449.4]
  wire  MyMem_io_wen; // @[CaheCore.scala 34:43:@2449.4]
  wire [5:0] MyMem_io_addr; // @[CaheCore.scala 34:43:@2449.4]
  wire [31:0] MyMem_io_wdata; // @[CaheCore.scala 34:43:@2449.4]
  wire [31:0] MyMem_io_rdata; // @[CaheCore.scala 34:43:@2449.4]
  wire  MyMem_1_clock; // @[CaheCore.scala 34:43:@2452.4]
  wire  MyMem_1_io_wen; // @[CaheCore.scala 34:43:@2452.4]
  wire [5:0] MyMem_1_io_addr; // @[CaheCore.scala 34:43:@2452.4]
  wire [31:0] MyMem_1_io_wdata; // @[CaheCore.scala 34:43:@2452.4]
  wire [31:0] MyMem_1_io_rdata; // @[CaheCore.scala 34:43:@2452.4]
  wire  MyMem_2_clock; // @[CaheCore.scala 34:43:@2455.4]
  wire  MyMem_2_io_wen; // @[CaheCore.scala 34:43:@2455.4]
  wire [5:0] MyMem_2_io_addr; // @[CaheCore.scala 34:43:@2455.4]
  wire [31:0] MyMem_2_io_wdata; // @[CaheCore.scala 34:43:@2455.4]
  wire [31:0] MyMem_2_io_rdata; // @[CaheCore.scala 34:43:@2455.4]
  wire  MyMem_3_clock; // @[CaheCore.scala 34:43:@2458.4]
  wire  MyMem_3_io_wen; // @[CaheCore.scala 34:43:@2458.4]
  wire [5:0] MyMem_3_io_addr; // @[CaheCore.scala 34:43:@2458.4]
  wire [31:0] MyMem_3_io_wdata; // @[CaheCore.scala 34:43:@2458.4]
  wire [31:0] MyMem_3_io_rdata; // @[CaheCore.scala 34:43:@2458.4]
  wire  MyMem_4_clock; // @[CaheCore.scala 34:43:@2461.4]
  wire  MyMem_4_io_wen; // @[CaheCore.scala 34:43:@2461.4]
  wire [5:0] MyMem_4_io_addr; // @[CaheCore.scala 34:43:@2461.4]
  wire [31:0] MyMem_4_io_wdata; // @[CaheCore.scala 34:43:@2461.4]
  wire [31:0] MyMem_4_io_rdata; // @[CaheCore.scala 34:43:@2461.4]
  wire  MyMem_5_clock; // @[CaheCore.scala 34:43:@2464.4]
  wire  MyMem_5_io_wen; // @[CaheCore.scala 34:43:@2464.4]
  wire [5:0] MyMem_5_io_addr; // @[CaheCore.scala 34:43:@2464.4]
  wire [31:0] MyMem_5_io_wdata; // @[CaheCore.scala 34:43:@2464.4]
  wire [31:0] MyMem_5_io_rdata; // @[CaheCore.scala 34:43:@2464.4]
  wire  MyMem_6_clock; // @[CaheCore.scala 34:43:@2467.4]
  wire  MyMem_6_io_wen; // @[CaheCore.scala 34:43:@2467.4]
  wire [5:0] MyMem_6_io_addr; // @[CaheCore.scala 34:43:@2467.4]
  wire [31:0] MyMem_6_io_wdata; // @[CaheCore.scala 34:43:@2467.4]
  wire [31:0] MyMem_6_io_rdata; // @[CaheCore.scala 34:43:@2467.4]
  wire  MyMem_7_clock; // @[CaheCore.scala 34:43:@2470.4]
  wire  MyMem_7_io_wen; // @[CaheCore.scala 34:43:@2470.4]
  wire [5:0] MyMem_7_io_addr; // @[CaheCore.scala 34:43:@2470.4]
  wire [31:0] MyMem_7_io_wdata; // @[CaheCore.scala 34:43:@2470.4]
  wire [31:0] MyMem_7_io_rdata; // @[CaheCore.scala 34:43:@2470.4]
  wire  MyMem_8_clock; // @[CaheCore.scala 34:43:@2473.4]
  wire  MyMem_8_io_wen; // @[CaheCore.scala 34:43:@2473.4]
  wire [5:0] MyMem_8_io_addr; // @[CaheCore.scala 34:43:@2473.4]
  wire [31:0] MyMem_8_io_wdata; // @[CaheCore.scala 34:43:@2473.4]
  wire [31:0] MyMem_8_io_rdata; // @[CaheCore.scala 34:43:@2473.4]
  wire  MyMem_9_clock; // @[CaheCore.scala 34:43:@2476.4]
  wire  MyMem_9_io_wen; // @[CaheCore.scala 34:43:@2476.4]
  wire [5:0] MyMem_9_io_addr; // @[CaheCore.scala 34:43:@2476.4]
  wire [31:0] MyMem_9_io_wdata; // @[CaheCore.scala 34:43:@2476.4]
  wire [31:0] MyMem_9_io_rdata; // @[CaheCore.scala 34:43:@2476.4]
  wire  MyMem_10_clock; // @[CaheCore.scala 34:43:@2479.4]
  wire  MyMem_10_io_wen; // @[CaheCore.scala 34:43:@2479.4]
  wire [5:0] MyMem_10_io_addr; // @[CaheCore.scala 34:43:@2479.4]
  wire [31:0] MyMem_10_io_wdata; // @[CaheCore.scala 34:43:@2479.4]
  wire [31:0] MyMem_10_io_rdata; // @[CaheCore.scala 34:43:@2479.4]
  wire  MyMem_11_clock; // @[CaheCore.scala 34:43:@2482.4]
  wire  MyMem_11_io_wen; // @[CaheCore.scala 34:43:@2482.4]
  wire [5:0] MyMem_11_io_addr; // @[CaheCore.scala 34:43:@2482.4]
  wire [31:0] MyMem_11_io_wdata; // @[CaheCore.scala 34:43:@2482.4]
  wire [31:0] MyMem_11_io_rdata; // @[CaheCore.scala 34:43:@2482.4]
  wire  MyMem_12_clock; // @[CaheCore.scala 34:43:@2485.4]
  wire  MyMem_12_io_wen; // @[CaheCore.scala 34:43:@2485.4]
  wire [5:0] MyMem_12_io_addr; // @[CaheCore.scala 34:43:@2485.4]
  wire [31:0] MyMem_12_io_wdata; // @[CaheCore.scala 34:43:@2485.4]
  wire [31:0] MyMem_12_io_rdata; // @[CaheCore.scala 34:43:@2485.4]
  wire  MyMem_13_clock; // @[CaheCore.scala 34:43:@2488.4]
  wire  MyMem_13_io_wen; // @[CaheCore.scala 34:43:@2488.4]
  wire [5:0] MyMem_13_io_addr; // @[CaheCore.scala 34:43:@2488.4]
  wire [31:0] MyMem_13_io_wdata; // @[CaheCore.scala 34:43:@2488.4]
  wire [31:0] MyMem_13_io_rdata; // @[CaheCore.scala 34:43:@2488.4]
  wire  MyMem_14_clock; // @[CaheCore.scala 34:43:@2491.4]
  wire  MyMem_14_io_wen; // @[CaheCore.scala 34:43:@2491.4]
  wire [5:0] MyMem_14_io_addr; // @[CaheCore.scala 34:43:@2491.4]
  wire [31:0] MyMem_14_io_wdata; // @[CaheCore.scala 34:43:@2491.4]
  wire [31:0] MyMem_14_io_rdata; // @[CaheCore.scala 34:43:@2491.4]
  wire  MyMem_15_clock; // @[CaheCore.scala 34:43:@2494.4]
  wire  MyMem_15_io_wen; // @[CaheCore.scala 34:43:@2494.4]
  wire [5:0] MyMem_15_io_addr; // @[CaheCore.scala 34:43:@2494.4]
  wire [31:0] MyMem_15_io_wdata; // @[CaheCore.scala 34:43:@2494.4]
  wire [31:0] MyMem_15_io_rdata; // @[CaheCore.scala 34:43:@2494.4]
  reg [19:0] tag_RAM [0:63]; // @[CaheCore.scala 35:30:@2497.4]
  reg [31:0] _RAND_0;
  wire [19:0] tag_RAM_rtag_data; // @[CaheCore.scala 35:30:@2497.4]
  wire [5:0] tag_RAM_rtag_addr; // @[CaheCore.scala 35:30:@2497.4]
  wire [19:0] tag_RAM__T_550_data; // @[CaheCore.scala 35:30:@2497.4]
  wire [5:0] tag_RAM__T_550_addr; // @[CaheCore.scala 35:30:@2497.4]
  wire  tag_RAM__T_550_mask; // @[CaheCore.scala 35:30:@2497.4]
  wire  tag_RAM__T_550_en; // @[CaheCore.scala 35:30:@2497.4]
  reg  statusVec_0; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_1;
  reg  statusVec_1; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_2;
  reg  statusVec_2; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_3;
  reg  statusVec_3; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_4;
  reg  statusVec_4; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_5;
  reg  statusVec_5; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_6;
  reg  statusVec_6; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_7;
  reg  statusVec_7; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_8;
  reg  statusVec_8; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_9;
  reg  statusVec_9; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_10;
  reg  statusVec_10; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_11;
  reg  statusVec_11; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_12;
  reg  statusVec_12; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_13;
  reg  statusVec_13; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_14;
  reg  statusVec_14; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_15;
  reg  statusVec_15; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_16;
  reg  statusVec_16; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_17;
  reg  statusVec_17; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_18;
  reg  statusVec_18; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_19;
  reg  statusVec_19; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_20;
  reg  statusVec_20; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_21;
  reg  statusVec_21; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_22;
  reg  statusVec_22; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_23;
  reg  statusVec_23; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_24;
  reg  statusVec_24; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_25;
  reg  statusVec_25; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_26;
  reg  statusVec_26; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_27;
  reg  statusVec_27; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_28;
  reg  statusVec_28; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_29;
  reg  statusVec_29; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_30;
  reg  statusVec_30; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_31;
  reg  statusVec_31; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_32;
  reg  statusVec_32; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_33;
  reg  statusVec_33; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_34;
  reg  statusVec_34; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_35;
  reg  statusVec_35; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_36;
  reg  statusVec_36; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_37;
  reg  statusVec_37; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_38;
  reg  statusVec_38; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_39;
  reg  statusVec_39; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_40;
  reg  statusVec_40; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_41;
  reg  statusVec_41; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_42;
  reg  statusVec_42; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_43;
  reg  statusVec_43; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_44;
  reg  statusVec_44; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_45;
  reg  statusVec_45; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_46;
  reg  statusVec_46; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_47;
  reg  statusVec_47; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_48;
  reg  statusVec_48; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_49;
  reg  statusVec_49; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_50;
  reg  statusVec_50; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_51;
  reg  statusVec_51; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_52;
  reg  statusVec_52; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_53;
  reg  statusVec_53; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_54;
  reg  statusVec_54; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_55;
  reg  statusVec_55; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_56;
  reg  statusVec_56; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_57;
  reg  statusVec_57; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_58;
  reg  statusVec_58; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_59;
  reg  statusVec_59; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_60;
  reg  statusVec_60; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_61;
  reg  statusVec_61; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_62;
  reg  statusVec_62; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_63;
  reg  statusVec_63; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_64;
  reg [3:0] line_idx; // @[CaheCore.scala 37:26:@2565.4]
  reg [31:0] _RAND_65;
  wire [5:0] off_idx; // @[CaheCore.scala 40:25:@2568.4]
  reg  rstatus; // @[CaheCore.scala 52:24:@2635.4]
  reg [31:0] _RAND_66;
  wire  _GEN_1; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_2; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_3; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_4; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_5; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_6; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_7; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_8; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_9; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_10; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_11; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_12; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_13; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_14; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_15; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_16; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_17; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_18; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_19; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_20; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_21; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_22; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_23; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_24; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_25; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_26; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_27; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_28; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_29; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_30; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_31; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_32; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_33; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_34; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_35; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_36; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_37; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_38; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_39; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_40; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_41; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_42; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_43; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_44; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_45; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_46; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_47; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_48; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_49; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_50; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_51; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_52; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_53; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_54; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_55; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_56; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_57; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_58; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_59; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_60; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_61; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_62; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_67; // @[CaheCore.scala 54:16:@2637.4]
  wire  _GEN_69; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_70; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_71; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_72; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_73; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_74; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_75; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_76; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_77; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_78; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_79; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_80; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_81; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_82; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_83; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_84; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_85; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_86; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_87; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_88; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_89; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_90; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_91; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_92; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_93; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_94; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_95; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_96; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_97; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_98; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_99; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_100; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_101; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_102; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_103; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_104; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_105; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_106; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_107; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_108; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_109; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_110; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_111; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_112; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_113; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_114; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_115; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_116; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_117; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_118; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_119; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_120; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_121; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_122; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_123; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_124; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_125; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_126; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_127; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_128; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_129; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_130; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_131; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_132; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_133; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_134; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_135; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_136; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_137; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_138; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_139; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_140; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_141; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_142; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_143; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_144; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_145; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_146; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_147; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_148; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_149; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_150; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_151; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_152; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_153; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_154; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_155; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_156; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_157; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_158; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_159; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_160; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_161; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_162; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_163; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_164; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_165; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_166; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_167; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_168; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_169; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_170; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_171; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_172; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_173; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_174; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_175; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_176; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_177; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_178; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_179; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_180; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_181; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_182; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_183; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_184; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_185; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_186; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_187; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_188; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_189; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_190; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_191; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_192; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_193; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_194; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_195; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_196; // @[CaheCore.scala 55:16:@2642.4]
  reg [19:0] tag; // @[CaheCore.scala 57:23:@2645.4]
  reg [31:0] _RAND_67;
  wire [31:0] rdata_0; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2573.4]
  wire [31:0] rdata_1; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2577.4]
  wire [31:0] _GEN_198; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_2; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2581.4]
  wire [31:0] _GEN_199; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_3; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2585.4]
  wire [31:0] _GEN_200; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_4; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2589.4]
  wire [31:0] _GEN_201; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_5; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2593.4]
  wire [31:0] _GEN_202; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_6; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2597.4]
  wire [31:0] _GEN_203; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_7; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2601.4]
  wire [31:0] _GEN_204; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_8; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2605.4]
  wire [31:0] _GEN_205; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_9; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2609.4]
  wire [31:0] _GEN_206; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_10; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2613.4]
  wire [31:0] _GEN_207; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_11; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2617.4]
  wire [31:0] _GEN_208; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_12; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2621.4]
  wire [31:0] _GEN_209; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_13; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2625.4]
  wire [31:0] _GEN_210; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_14; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2629.4]
  wire [31:0] _GEN_211; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_15; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2633.4]
  wire  _T_560; // @[CaheCore.scala 59:21:@2650.4]
  reg [5:0] tag_RAM_rtag_addr_pipe_0;
  reg [31:0] _RAND_68;
  MyMem MyMem ( // @[CaheCore.scala 34:43:@2449.4]
    .clock(MyMem_clock),
    .io_wen(MyMem_io_wen),
    .io_addr(MyMem_io_addr),
    .io_wdata(MyMem_io_wdata),
    .io_rdata(MyMem_io_rdata)
  );
  MyMem MyMem_1 ( // @[CaheCore.scala 34:43:@2452.4]
    .clock(MyMem_1_clock),
    .io_wen(MyMem_1_io_wen),
    .io_addr(MyMem_1_io_addr),
    .io_wdata(MyMem_1_io_wdata),
    .io_rdata(MyMem_1_io_rdata)
  );
  MyMem MyMem_2 ( // @[CaheCore.scala 34:43:@2455.4]
    .clock(MyMem_2_clock),
    .io_wen(MyMem_2_io_wen),
    .io_addr(MyMem_2_io_addr),
    .io_wdata(MyMem_2_io_wdata),
    .io_rdata(MyMem_2_io_rdata)
  );
  MyMem MyMem_3 ( // @[CaheCore.scala 34:43:@2458.4]
    .clock(MyMem_3_clock),
    .io_wen(MyMem_3_io_wen),
    .io_addr(MyMem_3_io_addr),
    .io_wdata(MyMem_3_io_wdata),
    .io_rdata(MyMem_3_io_rdata)
  );
  MyMem MyMem_4 ( // @[CaheCore.scala 34:43:@2461.4]
    .clock(MyMem_4_clock),
    .io_wen(MyMem_4_io_wen),
    .io_addr(MyMem_4_io_addr),
    .io_wdata(MyMem_4_io_wdata),
    .io_rdata(MyMem_4_io_rdata)
  );
  MyMem MyMem_5 ( // @[CaheCore.scala 34:43:@2464.4]
    .clock(MyMem_5_clock),
    .io_wen(MyMem_5_io_wen),
    .io_addr(MyMem_5_io_addr),
    .io_wdata(MyMem_5_io_wdata),
    .io_rdata(MyMem_5_io_rdata)
  );
  MyMem MyMem_6 ( // @[CaheCore.scala 34:43:@2467.4]
    .clock(MyMem_6_clock),
    .io_wen(MyMem_6_io_wen),
    .io_addr(MyMem_6_io_addr),
    .io_wdata(MyMem_6_io_wdata),
    .io_rdata(MyMem_6_io_rdata)
  );
  MyMem MyMem_7 ( // @[CaheCore.scala 34:43:@2470.4]
    .clock(MyMem_7_clock),
    .io_wen(MyMem_7_io_wen),
    .io_addr(MyMem_7_io_addr),
    .io_wdata(MyMem_7_io_wdata),
    .io_rdata(MyMem_7_io_rdata)
  );
  MyMem MyMem_8 ( // @[CaheCore.scala 34:43:@2473.4]
    .clock(MyMem_8_clock),
    .io_wen(MyMem_8_io_wen),
    .io_addr(MyMem_8_io_addr),
    .io_wdata(MyMem_8_io_wdata),
    .io_rdata(MyMem_8_io_rdata)
  );
  MyMem MyMem_9 ( // @[CaheCore.scala 34:43:@2476.4]
    .clock(MyMem_9_clock),
    .io_wen(MyMem_9_io_wen),
    .io_addr(MyMem_9_io_addr),
    .io_wdata(MyMem_9_io_wdata),
    .io_rdata(MyMem_9_io_rdata)
  );
  MyMem MyMem_10 ( // @[CaheCore.scala 34:43:@2479.4]
    .clock(MyMem_10_clock),
    .io_wen(MyMem_10_io_wen),
    .io_addr(MyMem_10_io_addr),
    .io_wdata(MyMem_10_io_wdata),
    .io_rdata(MyMem_10_io_rdata)
  );
  MyMem MyMem_11 ( // @[CaheCore.scala 34:43:@2482.4]
    .clock(MyMem_11_clock),
    .io_wen(MyMem_11_io_wen),
    .io_addr(MyMem_11_io_addr),
    .io_wdata(MyMem_11_io_wdata),
    .io_rdata(MyMem_11_io_rdata)
  );
  MyMem MyMem_12 ( // @[CaheCore.scala 34:43:@2485.4]
    .clock(MyMem_12_clock),
    .io_wen(MyMem_12_io_wen),
    .io_addr(MyMem_12_io_addr),
    .io_wdata(MyMem_12_io_wdata),
    .io_rdata(MyMem_12_io_rdata)
  );
  MyMem MyMem_13 ( // @[CaheCore.scala 34:43:@2488.4]
    .clock(MyMem_13_clock),
    .io_wen(MyMem_13_io_wen),
    .io_addr(MyMem_13_io_addr),
    .io_wdata(MyMem_13_io_wdata),
    .io_rdata(MyMem_13_io_rdata)
  );
  MyMem MyMem_14 ( // @[CaheCore.scala 34:43:@2491.4]
    .clock(MyMem_14_clock),
    .io_wen(MyMem_14_io_wen),
    .io_addr(MyMem_14_io_addr),
    .io_wdata(MyMem_14_io_wdata),
    .io_rdata(MyMem_14_io_rdata)
  );
  MyMem MyMem_15 ( // @[CaheCore.scala 34:43:@2494.4]
    .clock(MyMem_15_clock),
    .io_wen(MyMem_15_io_wen),
    .io_addr(MyMem_15_io_addr),
    .io_wdata(MyMem_15_io_wdata),
    .io_rdata(MyMem_15_io_rdata)
  );
  assign tag_RAM_rtag_addr = tag_RAM_rtag_addr_pipe_0;
  assign tag_RAM_rtag_data = tag_RAM[tag_RAM_rtag_addr]; // @[CaheCore.scala 35:30:@2497.4]
  assign tag_RAM__T_550_data = io_addr[31:12];
  assign tag_RAM__T_550_addr = io_addr[11:6];
  assign tag_RAM__T_550_mask = 1'h1;
  assign tag_RAM__T_550_en = io_wen;
  assign off_idx = io_addr[11:6]; // @[CaheCore.scala 40:25:@2568.4]
  assign _GEN_1 = 6'h1 == off_idx ? statusVec_1 : statusVec_0; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_2 = 6'h2 == off_idx ? statusVec_2 : _GEN_1; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_3 = 6'h3 == off_idx ? statusVec_3 : _GEN_2; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_4 = 6'h4 == off_idx ? statusVec_4 : _GEN_3; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_5 = 6'h5 == off_idx ? statusVec_5 : _GEN_4; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_6 = 6'h6 == off_idx ? statusVec_6 : _GEN_5; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_7 = 6'h7 == off_idx ? statusVec_7 : _GEN_6; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_8 = 6'h8 == off_idx ? statusVec_8 : _GEN_7; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_9 = 6'h9 == off_idx ? statusVec_9 : _GEN_8; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_10 = 6'ha == off_idx ? statusVec_10 : _GEN_9; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_11 = 6'hb == off_idx ? statusVec_11 : _GEN_10; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_12 = 6'hc == off_idx ? statusVec_12 : _GEN_11; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_13 = 6'hd == off_idx ? statusVec_13 : _GEN_12; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_14 = 6'he == off_idx ? statusVec_14 : _GEN_13; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_15 = 6'hf == off_idx ? statusVec_15 : _GEN_14; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_16 = 6'h10 == off_idx ? statusVec_16 : _GEN_15; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_17 = 6'h11 == off_idx ? statusVec_17 : _GEN_16; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_18 = 6'h12 == off_idx ? statusVec_18 : _GEN_17; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_19 = 6'h13 == off_idx ? statusVec_19 : _GEN_18; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_20 = 6'h14 == off_idx ? statusVec_20 : _GEN_19; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_21 = 6'h15 == off_idx ? statusVec_21 : _GEN_20; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_22 = 6'h16 == off_idx ? statusVec_22 : _GEN_21; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_23 = 6'h17 == off_idx ? statusVec_23 : _GEN_22; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_24 = 6'h18 == off_idx ? statusVec_24 : _GEN_23; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_25 = 6'h19 == off_idx ? statusVec_25 : _GEN_24; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_26 = 6'h1a == off_idx ? statusVec_26 : _GEN_25; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_27 = 6'h1b == off_idx ? statusVec_27 : _GEN_26; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_28 = 6'h1c == off_idx ? statusVec_28 : _GEN_27; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_29 = 6'h1d == off_idx ? statusVec_29 : _GEN_28; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_30 = 6'h1e == off_idx ? statusVec_30 : _GEN_29; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_31 = 6'h1f == off_idx ? statusVec_31 : _GEN_30; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_32 = 6'h20 == off_idx ? statusVec_32 : _GEN_31; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_33 = 6'h21 == off_idx ? statusVec_33 : _GEN_32; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_34 = 6'h22 == off_idx ? statusVec_34 : _GEN_33; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_35 = 6'h23 == off_idx ? statusVec_35 : _GEN_34; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_36 = 6'h24 == off_idx ? statusVec_36 : _GEN_35; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_37 = 6'h25 == off_idx ? statusVec_37 : _GEN_36; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_38 = 6'h26 == off_idx ? statusVec_38 : _GEN_37; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_39 = 6'h27 == off_idx ? statusVec_39 : _GEN_38; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_40 = 6'h28 == off_idx ? statusVec_40 : _GEN_39; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_41 = 6'h29 == off_idx ? statusVec_41 : _GEN_40; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_42 = 6'h2a == off_idx ? statusVec_42 : _GEN_41; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_43 = 6'h2b == off_idx ? statusVec_43 : _GEN_42; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_44 = 6'h2c == off_idx ? statusVec_44 : _GEN_43; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_45 = 6'h2d == off_idx ? statusVec_45 : _GEN_44; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_46 = 6'h2e == off_idx ? statusVec_46 : _GEN_45; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_47 = 6'h2f == off_idx ? statusVec_47 : _GEN_46; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_48 = 6'h30 == off_idx ? statusVec_48 : _GEN_47; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_49 = 6'h31 == off_idx ? statusVec_49 : _GEN_48; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_50 = 6'h32 == off_idx ? statusVec_50 : _GEN_49; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_51 = 6'h33 == off_idx ? statusVec_51 : _GEN_50; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_52 = 6'h34 == off_idx ? statusVec_52 : _GEN_51; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_53 = 6'h35 == off_idx ? statusVec_53 : _GEN_52; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_54 = 6'h36 == off_idx ? statusVec_54 : _GEN_53; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_55 = 6'h37 == off_idx ? statusVec_55 : _GEN_54; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_56 = 6'h38 == off_idx ? statusVec_56 : _GEN_55; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_57 = 6'h39 == off_idx ? statusVec_57 : _GEN_56; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_58 = 6'h3a == off_idx ? statusVec_58 : _GEN_57; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_59 = 6'h3b == off_idx ? statusVec_59 : _GEN_58; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_60 = 6'h3c == off_idx ? statusVec_60 : _GEN_59; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_61 = 6'h3d == off_idx ? statusVec_61 : _GEN_60; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_62 = 6'h3e == off_idx ? statusVec_62 : _GEN_61; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_67 = 1'h1; // @[CaheCore.scala 54:16:@2637.4]
  assign _GEN_69 = 6'h0 == off_idx ? io_wstatus : statusVec_0; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_70 = 6'h1 == off_idx ? io_wstatus : statusVec_1; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_71 = 6'h2 == off_idx ? io_wstatus : statusVec_2; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_72 = 6'h3 == off_idx ? io_wstatus : statusVec_3; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_73 = 6'h4 == off_idx ? io_wstatus : statusVec_4; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_74 = 6'h5 == off_idx ? io_wstatus : statusVec_5; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_75 = 6'h6 == off_idx ? io_wstatus : statusVec_6; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_76 = 6'h7 == off_idx ? io_wstatus : statusVec_7; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_77 = 6'h8 == off_idx ? io_wstatus : statusVec_8; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_78 = 6'h9 == off_idx ? io_wstatus : statusVec_9; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_79 = 6'ha == off_idx ? io_wstatus : statusVec_10; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_80 = 6'hb == off_idx ? io_wstatus : statusVec_11; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_81 = 6'hc == off_idx ? io_wstatus : statusVec_12; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_82 = 6'hd == off_idx ? io_wstatus : statusVec_13; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_83 = 6'he == off_idx ? io_wstatus : statusVec_14; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_84 = 6'hf == off_idx ? io_wstatus : statusVec_15; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_85 = 6'h10 == off_idx ? io_wstatus : statusVec_16; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_86 = 6'h11 == off_idx ? io_wstatus : statusVec_17; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_87 = 6'h12 == off_idx ? io_wstatus : statusVec_18; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_88 = 6'h13 == off_idx ? io_wstatus : statusVec_19; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_89 = 6'h14 == off_idx ? io_wstatus : statusVec_20; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_90 = 6'h15 == off_idx ? io_wstatus : statusVec_21; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_91 = 6'h16 == off_idx ? io_wstatus : statusVec_22; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_92 = 6'h17 == off_idx ? io_wstatus : statusVec_23; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_93 = 6'h18 == off_idx ? io_wstatus : statusVec_24; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_94 = 6'h19 == off_idx ? io_wstatus : statusVec_25; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_95 = 6'h1a == off_idx ? io_wstatus : statusVec_26; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_96 = 6'h1b == off_idx ? io_wstatus : statusVec_27; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_97 = 6'h1c == off_idx ? io_wstatus : statusVec_28; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_98 = 6'h1d == off_idx ? io_wstatus : statusVec_29; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_99 = 6'h1e == off_idx ? io_wstatus : statusVec_30; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_100 = 6'h1f == off_idx ? io_wstatus : statusVec_31; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_101 = 6'h20 == off_idx ? io_wstatus : statusVec_32; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_102 = 6'h21 == off_idx ? io_wstatus : statusVec_33; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_103 = 6'h22 == off_idx ? io_wstatus : statusVec_34; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_104 = 6'h23 == off_idx ? io_wstatus : statusVec_35; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_105 = 6'h24 == off_idx ? io_wstatus : statusVec_36; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_106 = 6'h25 == off_idx ? io_wstatus : statusVec_37; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_107 = 6'h26 == off_idx ? io_wstatus : statusVec_38; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_108 = 6'h27 == off_idx ? io_wstatus : statusVec_39; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_109 = 6'h28 == off_idx ? io_wstatus : statusVec_40; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_110 = 6'h29 == off_idx ? io_wstatus : statusVec_41; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_111 = 6'h2a == off_idx ? io_wstatus : statusVec_42; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_112 = 6'h2b == off_idx ? io_wstatus : statusVec_43; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_113 = 6'h2c == off_idx ? io_wstatus : statusVec_44; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_114 = 6'h2d == off_idx ? io_wstatus : statusVec_45; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_115 = 6'h2e == off_idx ? io_wstatus : statusVec_46; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_116 = 6'h2f == off_idx ? io_wstatus : statusVec_47; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_117 = 6'h30 == off_idx ? io_wstatus : statusVec_48; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_118 = 6'h31 == off_idx ? io_wstatus : statusVec_49; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_119 = 6'h32 == off_idx ? io_wstatus : statusVec_50; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_120 = 6'h33 == off_idx ? io_wstatus : statusVec_51; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_121 = 6'h34 == off_idx ? io_wstatus : statusVec_52; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_122 = 6'h35 == off_idx ? io_wstatus : statusVec_53; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_123 = 6'h36 == off_idx ? io_wstatus : statusVec_54; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_124 = 6'h37 == off_idx ? io_wstatus : statusVec_55; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_125 = 6'h38 == off_idx ? io_wstatus : statusVec_56; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_126 = 6'h39 == off_idx ? io_wstatus : statusVec_57; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_127 = 6'h3a == off_idx ? io_wstatus : statusVec_58; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_128 = 6'h3b == off_idx ? io_wstatus : statusVec_59; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_129 = 6'h3c == off_idx ? io_wstatus : statusVec_60; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_130 = 6'h3d == off_idx ? io_wstatus : statusVec_61; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_131 = 6'h3e == off_idx ? io_wstatus : statusVec_62; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_132 = 6'h3f == off_idx ? io_wstatus : statusVec_63; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_133 = io_wen ? _GEN_69 : statusVec_0; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_134 = io_wen ? _GEN_70 : statusVec_1; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_135 = io_wen ? _GEN_71 : statusVec_2; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_136 = io_wen ? _GEN_72 : statusVec_3; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_137 = io_wen ? _GEN_73 : statusVec_4; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_138 = io_wen ? _GEN_74 : statusVec_5; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_139 = io_wen ? _GEN_75 : statusVec_6; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_140 = io_wen ? _GEN_76 : statusVec_7; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_141 = io_wen ? _GEN_77 : statusVec_8; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_142 = io_wen ? _GEN_78 : statusVec_9; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_143 = io_wen ? _GEN_79 : statusVec_10; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_144 = io_wen ? _GEN_80 : statusVec_11; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_145 = io_wen ? _GEN_81 : statusVec_12; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_146 = io_wen ? _GEN_82 : statusVec_13; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_147 = io_wen ? _GEN_83 : statusVec_14; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_148 = io_wen ? _GEN_84 : statusVec_15; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_149 = io_wen ? _GEN_85 : statusVec_16; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_150 = io_wen ? _GEN_86 : statusVec_17; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_151 = io_wen ? _GEN_87 : statusVec_18; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_152 = io_wen ? _GEN_88 : statusVec_19; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_153 = io_wen ? _GEN_89 : statusVec_20; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_154 = io_wen ? _GEN_90 : statusVec_21; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_155 = io_wen ? _GEN_91 : statusVec_22; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_156 = io_wen ? _GEN_92 : statusVec_23; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_157 = io_wen ? _GEN_93 : statusVec_24; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_158 = io_wen ? _GEN_94 : statusVec_25; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_159 = io_wen ? _GEN_95 : statusVec_26; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_160 = io_wen ? _GEN_96 : statusVec_27; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_161 = io_wen ? _GEN_97 : statusVec_28; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_162 = io_wen ? _GEN_98 : statusVec_29; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_163 = io_wen ? _GEN_99 : statusVec_30; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_164 = io_wen ? _GEN_100 : statusVec_31; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_165 = io_wen ? _GEN_101 : statusVec_32; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_166 = io_wen ? _GEN_102 : statusVec_33; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_167 = io_wen ? _GEN_103 : statusVec_34; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_168 = io_wen ? _GEN_104 : statusVec_35; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_169 = io_wen ? _GEN_105 : statusVec_36; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_170 = io_wen ? _GEN_106 : statusVec_37; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_171 = io_wen ? _GEN_107 : statusVec_38; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_172 = io_wen ? _GEN_108 : statusVec_39; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_173 = io_wen ? _GEN_109 : statusVec_40; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_174 = io_wen ? _GEN_110 : statusVec_41; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_175 = io_wen ? _GEN_111 : statusVec_42; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_176 = io_wen ? _GEN_112 : statusVec_43; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_177 = io_wen ? _GEN_113 : statusVec_44; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_178 = io_wen ? _GEN_114 : statusVec_45; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_179 = io_wen ? _GEN_115 : statusVec_46; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_180 = io_wen ? _GEN_116 : statusVec_47; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_181 = io_wen ? _GEN_117 : statusVec_48; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_182 = io_wen ? _GEN_118 : statusVec_49; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_183 = io_wen ? _GEN_119 : statusVec_50; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_184 = io_wen ? _GEN_120 : statusVec_51; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_185 = io_wen ? _GEN_121 : statusVec_52; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_186 = io_wen ? _GEN_122 : statusVec_53; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_187 = io_wen ? _GEN_123 : statusVec_54; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_188 = io_wen ? _GEN_124 : statusVec_55; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_189 = io_wen ? _GEN_125 : statusVec_56; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_190 = io_wen ? _GEN_126 : statusVec_57; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_191 = io_wen ? _GEN_127 : statusVec_58; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_192 = io_wen ? _GEN_128 : statusVec_59; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_193 = io_wen ? _GEN_129 : statusVec_60; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_194 = io_wen ? _GEN_130 : statusVec_61; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_195 = io_wen ? _GEN_131 : statusVec_62; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_196 = io_wen ? _GEN_132 : statusVec_63; // @[CaheCore.scala 55:16:@2642.4]
  assign rdata_0 = MyMem_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2573.4]
  assign rdata_1 = MyMem_1_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2577.4]
  assign _GEN_198 = 4'h1 == line_idx ? rdata_1 : rdata_0; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_2 = MyMem_2_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2581.4]
  assign _GEN_199 = 4'h2 == line_idx ? rdata_2 : _GEN_198; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_3 = MyMem_3_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2585.4]
  assign _GEN_200 = 4'h3 == line_idx ? rdata_3 : _GEN_199; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_4 = MyMem_4_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2589.4]
  assign _GEN_201 = 4'h4 == line_idx ? rdata_4 : _GEN_200; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_5 = MyMem_5_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2593.4]
  assign _GEN_202 = 4'h5 == line_idx ? rdata_5 : _GEN_201; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_6 = MyMem_6_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2597.4]
  assign _GEN_203 = 4'h6 == line_idx ? rdata_6 : _GEN_202; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_7 = MyMem_7_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2601.4]
  assign _GEN_204 = 4'h7 == line_idx ? rdata_7 : _GEN_203; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_8 = MyMem_8_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2605.4]
  assign _GEN_205 = 4'h8 == line_idx ? rdata_8 : _GEN_204; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_9 = MyMem_9_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2609.4]
  assign _GEN_206 = 4'h9 == line_idx ? rdata_9 : _GEN_205; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_10 = MyMem_10_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2613.4]
  assign _GEN_207 = 4'ha == line_idx ? rdata_10 : _GEN_206; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_11 = MyMem_11_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2617.4]
  assign _GEN_208 = 4'hb == line_idx ? rdata_11 : _GEN_207; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_12 = MyMem_12_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2621.4]
  assign _GEN_209 = 4'hc == line_idx ? rdata_12 : _GEN_208; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_13 = MyMem_13_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2625.4]
  assign _GEN_210 = 4'hd == line_idx ? rdata_13 : _GEN_209; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_14 = MyMem_14_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2629.4]
  assign _GEN_211 = 4'he == line_idx ? rdata_14 : _GEN_210; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_15 = MyMem_15_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2633.4]
  assign _T_560 = tag_RAM_rtag_data == tag; // @[CaheCore.scala 59:21:@2650.4]
  assign io_rdata = 4'hf == line_idx ? rdata_15 : _GEN_211; // @[CaheCore.scala 58:13:@2649.4]
  assign io_rvalid = _T_560 & rstatus; // @[CaheCore.scala 59:13:@2652.4]
  assign MyMem_clock = clock; // @[:@2450.4]
  assign MyMem_io_wen = io_wen; // @[CaheCore.scala 46:24:@2571.4]
  assign MyMem_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2570.4]
  assign MyMem_io_wdata = io_wdata_0; // @[CaheCore.scala 47:24:@2572.4]
  assign MyMem_1_clock = clock; // @[:@2453.4]
  assign MyMem_1_io_wen = io_wen; // @[CaheCore.scala 46:24:@2575.4]
  assign MyMem_1_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2574.4]
  assign MyMem_1_io_wdata = io_wdata_1; // @[CaheCore.scala 47:24:@2576.4]
  assign MyMem_2_clock = clock; // @[:@2456.4]
  assign MyMem_2_io_wen = io_wen; // @[CaheCore.scala 46:24:@2579.4]
  assign MyMem_2_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2578.4]
  assign MyMem_2_io_wdata = io_wdata_2; // @[CaheCore.scala 47:24:@2580.4]
  assign MyMem_3_clock = clock; // @[:@2459.4]
  assign MyMem_3_io_wen = io_wen; // @[CaheCore.scala 46:24:@2583.4]
  assign MyMem_3_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2582.4]
  assign MyMem_3_io_wdata = io_wdata_3; // @[CaheCore.scala 47:24:@2584.4]
  assign MyMem_4_clock = clock; // @[:@2462.4]
  assign MyMem_4_io_wen = io_wen; // @[CaheCore.scala 46:24:@2587.4]
  assign MyMem_4_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2586.4]
  assign MyMem_4_io_wdata = io_wdata_4; // @[CaheCore.scala 47:24:@2588.4]
  assign MyMem_5_clock = clock; // @[:@2465.4]
  assign MyMem_5_io_wen = io_wen; // @[CaheCore.scala 46:24:@2591.4]
  assign MyMem_5_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2590.4]
  assign MyMem_5_io_wdata = io_wdata_5; // @[CaheCore.scala 47:24:@2592.4]
  assign MyMem_6_clock = clock; // @[:@2468.4]
  assign MyMem_6_io_wen = io_wen; // @[CaheCore.scala 46:24:@2595.4]
  assign MyMem_6_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2594.4]
  assign MyMem_6_io_wdata = io_wdata_6; // @[CaheCore.scala 47:24:@2596.4]
  assign MyMem_7_clock = clock; // @[:@2471.4]
  assign MyMem_7_io_wen = io_wen; // @[CaheCore.scala 46:24:@2599.4]
  assign MyMem_7_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2598.4]
  assign MyMem_7_io_wdata = io_wdata_7; // @[CaheCore.scala 47:24:@2600.4]
  assign MyMem_8_clock = clock; // @[:@2474.4]
  assign MyMem_8_io_wen = io_wen; // @[CaheCore.scala 46:24:@2603.4]
  assign MyMem_8_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2602.4]
  assign MyMem_8_io_wdata = io_wdata_8; // @[CaheCore.scala 47:24:@2604.4]
  assign MyMem_9_clock = clock; // @[:@2477.4]
  assign MyMem_9_io_wen = io_wen; // @[CaheCore.scala 46:24:@2607.4]
  assign MyMem_9_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2606.4]
  assign MyMem_9_io_wdata = io_wdata_9; // @[CaheCore.scala 47:24:@2608.4]
  assign MyMem_10_clock = clock; // @[:@2480.4]
  assign MyMem_10_io_wen = io_wen; // @[CaheCore.scala 46:24:@2611.4]
  assign MyMem_10_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2610.4]
  assign MyMem_10_io_wdata = io_wdata_10; // @[CaheCore.scala 47:24:@2612.4]
  assign MyMem_11_clock = clock; // @[:@2483.4]
  assign MyMem_11_io_wen = io_wen; // @[CaheCore.scala 46:24:@2615.4]
  assign MyMem_11_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2614.4]
  assign MyMem_11_io_wdata = io_wdata_11; // @[CaheCore.scala 47:24:@2616.4]
  assign MyMem_12_clock = clock; // @[:@2486.4]
  assign MyMem_12_io_wen = io_wen; // @[CaheCore.scala 46:24:@2619.4]
  assign MyMem_12_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2618.4]
  assign MyMem_12_io_wdata = io_wdata_12; // @[CaheCore.scala 47:24:@2620.4]
  assign MyMem_13_clock = clock; // @[:@2489.4]
  assign MyMem_13_io_wen = io_wen; // @[CaheCore.scala 46:24:@2623.4]
  assign MyMem_13_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2622.4]
  assign MyMem_13_io_wdata = io_wdata_13; // @[CaheCore.scala 47:24:@2624.4]
  assign MyMem_14_clock = clock; // @[:@2492.4]
  assign MyMem_14_io_wen = io_wen; // @[CaheCore.scala 46:24:@2627.4]
  assign MyMem_14_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2626.4]
  assign MyMem_14_io_wdata = io_wdata_14; // @[CaheCore.scala 47:24:@2628.4]
  assign MyMem_15_clock = clock; // @[:@2495.4]
  assign MyMem_15_io_wen = io_wen; // @[CaheCore.scala 46:24:@2631.4]
  assign MyMem_15_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2630.4]
  assign MyMem_15_io_wdata = io_wdata_15; // @[CaheCore.scala 47:24:@2632.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_RAM[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  statusVec_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  statusVec_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  statusVec_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  statusVec_3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  statusVec_4 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  statusVec_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  statusVec_6 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  statusVec_7 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  statusVec_8 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  statusVec_9 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  statusVec_10 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  statusVec_11 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  statusVec_12 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  statusVec_13 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  statusVec_14 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  statusVec_15 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  statusVec_16 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  statusVec_17 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  statusVec_18 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  statusVec_19 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  statusVec_20 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  statusVec_21 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  statusVec_22 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  statusVec_23 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  statusVec_24 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  statusVec_25 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  statusVec_26 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  statusVec_27 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  statusVec_28 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  statusVec_29 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  statusVec_30 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  statusVec_31 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  statusVec_32 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  statusVec_33 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  statusVec_34 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  statusVec_35 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  statusVec_36 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  statusVec_37 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  statusVec_38 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  statusVec_39 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  statusVec_40 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  statusVec_41 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  statusVec_42 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  statusVec_43 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  statusVec_44 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  statusVec_45 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  statusVec_46 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  statusVec_47 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  statusVec_48 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  statusVec_49 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  statusVec_50 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  statusVec_51 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  statusVec_52 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  statusVec_53 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  statusVec_54 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  statusVec_55 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  statusVec_56 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  statusVec_57 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  statusVec_58 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  statusVec_59 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  statusVec_60 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  statusVec_61 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  statusVec_62 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  statusVec_63 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  line_idx = _RAND_65[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  rstatus = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tag = _RAND_67[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tag_RAM_rtag_addr_pipe_0 = _RAND_68[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tag_RAM__T_550_en & tag_RAM__T_550_mask) begin
      tag_RAM[tag_RAM__T_550_addr] <= tag_RAM__T_550_data; // @[CaheCore.scala 35:30:@2497.4]
    end
    if (reset) begin
      statusVec_0 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h0 == off_idx) begin
          statusVec_0 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_1 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1 == off_idx) begin
          statusVec_1 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_2 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2 == off_idx) begin
          statusVec_2 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_3 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3 == off_idx) begin
          statusVec_3 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_4 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h4 == off_idx) begin
          statusVec_4 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_5 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h5 == off_idx) begin
          statusVec_5 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_6 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h6 == off_idx) begin
          statusVec_6 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_7 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h7 == off_idx) begin
          statusVec_7 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_8 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h8 == off_idx) begin
          statusVec_8 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_9 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h9 == off_idx) begin
          statusVec_9 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_10 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'ha == off_idx) begin
          statusVec_10 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_11 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hb == off_idx) begin
          statusVec_11 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_12 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hc == off_idx) begin
          statusVec_12 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_13 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hd == off_idx) begin
          statusVec_13 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_14 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'he == off_idx) begin
          statusVec_14 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_15 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hf == off_idx) begin
          statusVec_15 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_16 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h10 == off_idx) begin
          statusVec_16 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_17 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h11 == off_idx) begin
          statusVec_17 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_18 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h12 == off_idx) begin
          statusVec_18 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_19 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h13 == off_idx) begin
          statusVec_19 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_20 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h14 == off_idx) begin
          statusVec_20 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_21 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h15 == off_idx) begin
          statusVec_21 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_22 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h16 == off_idx) begin
          statusVec_22 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_23 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h17 == off_idx) begin
          statusVec_23 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_24 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h18 == off_idx) begin
          statusVec_24 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_25 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h19 == off_idx) begin
          statusVec_25 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_26 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1a == off_idx) begin
          statusVec_26 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_27 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1b == off_idx) begin
          statusVec_27 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_28 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1c == off_idx) begin
          statusVec_28 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_29 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1d == off_idx) begin
          statusVec_29 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_30 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1e == off_idx) begin
          statusVec_30 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_31 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1f == off_idx) begin
          statusVec_31 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_32 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h20 == off_idx) begin
          statusVec_32 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_33 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h21 == off_idx) begin
          statusVec_33 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_34 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h22 == off_idx) begin
          statusVec_34 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_35 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h23 == off_idx) begin
          statusVec_35 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_36 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h24 == off_idx) begin
          statusVec_36 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_37 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h25 == off_idx) begin
          statusVec_37 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_38 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h26 == off_idx) begin
          statusVec_38 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_39 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h27 == off_idx) begin
          statusVec_39 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_40 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h28 == off_idx) begin
          statusVec_40 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_41 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h29 == off_idx) begin
          statusVec_41 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_42 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2a == off_idx) begin
          statusVec_42 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_43 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2b == off_idx) begin
          statusVec_43 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_44 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2c == off_idx) begin
          statusVec_44 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_45 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2d == off_idx) begin
          statusVec_45 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_46 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2e == off_idx) begin
          statusVec_46 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_47 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2f == off_idx) begin
          statusVec_47 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_48 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h30 == off_idx) begin
          statusVec_48 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_49 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h31 == off_idx) begin
          statusVec_49 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_50 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h32 == off_idx) begin
          statusVec_50 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_51 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h33 == off_idx) begin
          statusVec_51 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_52 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h34 == off_idx) begin
          statusVec_52 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_53 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h35 == off_idx) begin
          statusVec_53 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_54 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h36 == off_idx) begin
          statusVec_54 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_55 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h37 == off_idx) begin
          statusVec_55 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_56 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h38 == off_idx) begin
          statusVec_56 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_57 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h39 == off_idx) begin
          statusVec_57 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_58 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3a == off_idx) begin
          statusVec_58 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_59 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3b == off_idx) begin
          statusVec_59 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_60 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3c == off_idx) begin
          statusVec_60 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_61 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3d == off_idx) begin
          statusVec_61 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_62 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3e == off_idx) begin
          statusVec_62 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_63 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3f == off_idx) begin
          statusVec_63 <= io_wstatus;
        end
      end
    end
    line_idx <= io_addr[5:2];
    if (6'h3f == off_idx) begin
      rstatus <= statusVec_63;
    end else begin
      if (6'h3e == off_idx) begin
        rstatus <= statusVec_62;
      end else begin
        if (6'h3d == off_idx) begin
          rstatus <= statusVec_61;
        end else begin
          if (6'h3c == off_idx) begin
            rstatus <= statusVec_60;
          end else begin
            if (6'h3b == off_idx) begin
              rstatus <= statusVec_59;
            end else begin
              if (6'h3a == off_idx) begin
                rstatus <= statusVec_58;
              end else begin
                if (6'h39 == off_idx) begin
                  rstatus <= statusVec_57;
                end else begin
                  if (6'h38 == off_idx) begin
                    rstatus <= statusVec_56;
                  end else begin
                    if (6'h37 == off_idx) begin
                      rstatus <= statusVec_55;
                    end else begin
                      if (6'h36 == off_idx) begin
                        rstatus <= statusVec_54;
                      end else begin
                        if (6'h35 == off_idx) begin
                          rstatus <= statusVec_53;
                        end else begin
                          if (6'h34 == off_idx) begin
                            rstatus <= statusVec_52;
                          end else begin
                            if (6'h33 == off_idx) begin
                              rstatus <= statusVec_51;
                            end else begin
                              if (6'h32 == off_idx) begin
                                rstatus <= statusVec_50;
                              end else begin
                                if (6'h31 == off_idx) begin
                                  rstatus <= statusVec_49;
                                end else begin
                                  if (6'h30 == off_idx) begin
                                    rstatus <= statusVec_48;
                                  end else begin
                                    if (6'h2f == off_idx) begin
                                      rstatus <= statusVec_47;
                                    end else begin
                                      if (6'h2e == off_idx) begin
                                        rstatus <= statusVec_46;
                                      end else begin
                                        if (6'h2d == off_idx) begin
                                          rstatus <= statusVec_45;
                                        end else begin
                                          if (6'h2c == off_idx) begin
                                            rstatus <= statusVec_44;
                                          end else begin
                                            if (6'h2b == off_idx) begin
                                              rstatus <= statusVec_43;
                                            end else begin
                                              if (6'h2a == off_idx) begin
                                                rstatus <= statusVec_42;
                                              end else begin
                                                if (6'h29 == off_idx) begin
                                                  rstatus <= statusVec_41;
                                                end else begin
                                                  if (6'h28 == off_idx) begin
                                                    rstatus <= statusVec_40;
                                                  end else begin
                                                    if (6'h27 == off_idx) begin
                                                      rstatus <= statusVec_39;
                                                    end else begin
                                                      if (6'h26 == off_idx) begin
                                                        rstatus <= statusVec_38;
                                                      end else begin
                                                        if (6'h25 == off_idx) begin
                                                          rstatus <= statusVec_37;
                                                        end else begin
                                                          if (6'h24 == off_idx) begin
                                                            rstatus <= statusVec_36;
                                                          end else begin
                                                            if (6'h23 == off_idx) begin
                                                              rstatus <= statusVec_35;
                                                            end else begin
                                                              if (6'h22 == off_idx) begin
                                                                rstatus <= statusVec_34;
                                                              end else begin
                                                                if (6'h21 == off_idx) begin
                                                                  rstatus <= statusVec_33;
                                                                end else begin
                                                                  if (6'h20 == off_idx) begin
                                                                    rstatus <= statusVec_32;
                                                                  end else begin
                                                                    if (6'h1f == off_idx) begin
                                                                      rstatus <= statusVec_31;
                                                                    end else begin
                                                                      if (6'h1e == off_idx) begin
                                                                        rstatus <= statusVec_30;
                                                                      end else begin
                                                                        if (6'h1d == off_idx) begin
                                                                          rstatus <= statusVec_29;
                                                                        end else begin
                                                                          if (6'h1c == off_idx) begin
                                                                            rstatus <= statusVec_28;
                                                                          end else begin
                                                                            if (6'h1b == off_idx) begin
                                                                              rstatus <= statusVec_27;
                                                                            end else begin
                                                                              if (6'h1a == off_idx) begin
                                                                                rstatus <= statusVec_26;
                                                                              end else begin
                                                                                if (6'h19 == off_idx) begin
                                                                                  rstatus <= statusVec_25;
                                                                                end else begin
                                                                                  if (6'h18 == off_idx) begin
                                                                                    rstatus <= statusVec_24;
                                                                                  end else begin
                                                                                    if (6'h17 == off_idx) begin
                                                                                      rstatus <= statusVec_23;
                                                                                    end else begin
                                                                                      if (6'h16 == off_idx) begin
                                                                                        rstatus <= statusVec_22;
                                                                                      end else begin
                                                                                        if (6'h15 == off_idx) begin
                                                                                          rstatus <= statusVec_21;
                                                                                        end else begin
                                                                                          if (6'h14 == off_idx) begin
                                                                                            rstatus <= statusVec_20;
                                                                                          end else begin
                                                                                            if (6'h13 == off_idx) begin
                                                                                              rstatus <= statusVec_19;
                                                                                            end else begin
                                                                                              if (6'h12 == off_idx) begin
                                                                                                rstatus <= statusVec_18;
                                                                                              end else begin
                                                                                                if (6'h11 == off_idx) begin
                                                                                                  rstatus <= statusVec_17;
                                                                                                end else begin
                                                                                                  if (6'h10 == off_idx) begin
                                                                                                    rstatus <= statusVec_16;
                                                                                                  end else begin
                                                                                                    if (6'hf == off_idx) begin
                                                                                                      rstatus <= statusVec_15;
                                                                                                    end else begin
                                                                                                      if (6'he == off_idx) begin
                                                                                                        rstatus <= statusVec_14;
                                                                                                      end else begin
                                                                                                        if (6'hd == off_idx) begin
                                                                                                          rstatus <= statusVec_13;
                                                                                                        end else begin
                                                                                                          if (6'hc == off_idx) begin
                                                                                                            rstatus <= statusVec_12;
                                                                                                          end else begin
                                                                                                            if (6'hb == off_idx) begin
                                                                                                              rstatus <= statusVec_11;
                                                                                                            end else begin
                                                                                                              if (6'ha == off_idx) begin
                                                                                                                rstatus <= statusVec_10;
                                                                                                              end else begin
                                                                                                                if (6'h9 == off_idx) begin
                                                                                                                  rstatus <= statusVec_9;
                                                                                                                end else begin
                                                                                                                  if (6'h8 == off_idx) begin
                                                                                                                    rstatus <= statusVec_8;
                                                                                                                  end else begin
                                                                                                                    if (6'h7 == off_idx) begin
                                                                                                                      rstatus <= statusVec_7;
                                                                                                                    end else begin
                                                                                                                      if (6'h6 == off_idx) begin
                                                                                                                        rstatus <= statusVec_6;
                                                                                                                      end else begin
                                                                                                                        if (6'h5 == off_idx) begin
                                                                                                                          rstatus <= statusVec_5;
                                                                                                                        end else begin
                                                                                                                          if (6'h4 == off_idx) begin
                                                                                                                            rstatus <= statusVec_4;
                                                                                                                          end else begin
                                                                                                                            if (6'h3 == off_idx) begin
                                                                                                                              rstatus <= statusVec_3;
                                                                                                                            end else begin
                                                                                                                              if (6'h2 == off_idx) begin
                                                                                                                                rstatus <= statusVec_2;
                                                                                                                              end else begin
                                                                                                                                if (6'h1 == off_idx) begin
                                                                                                                                  rstatus <= statusVec_1;
                                                                                                                                end else begin
                                                                                                                                  rstatus <= statusVec_0;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    tag <= io_addr[31:12];
    if (_GEN_67) begin
      tag_RAM_rtag_addr_pipe_0 <= off_idx;
    end
  end
endmodule
module Icache( // @[:@2654.2]
  input         clock, // @[:@2655.4]
  input         reset, // @[:@2656.4]
  input         io_core_pc_valid, // @[:@2657.4]
  input  [31:0] io_core_pc_bits, // @[:@2657.4]
  output        io_core_inst_valid, // @[:@2657.4]
  output [31:0] io_core_inst_bits, // @[:@2657.4]
  output        io_core_ready, // @[:@2657.4]
  input  [31:0] io_axi_r_data, // @[:@2657.4]
  input         io_axi_r_valid, // @[:@2657.4]
  input         io_axi_r_last, // @[:@2657.4]
  input         io_axi_ar_ready, // @[:@2657.4]
  output        io_axi_ar_valid, // @[:@2657.4]
  output [31:0] io_axi_ar_addr // @[:@2657.4]
);
  wire  icache_clock; // @[Icache.scala 66:22:@2677.4]
  wire  icache_reset; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_wen; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_addr; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_0; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_1; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_2; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_3; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_4; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_5; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_6; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_7; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_8; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_9; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_10; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_11; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_12; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_13; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_14; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_15; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_wstatus; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_rdata; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_rvalid; // @[Icache.scala 66:22:@2677.4]
  reg  pc_valid; // @[Icache.scala 56:25:@2667.4]
  reg [31:0] _RAND_0;
  reg [31:0] pc; // @[Icache.scala 57:15:@2668.4]
  reg [31:0] _RAND_1;
  wire  pc_accept; // @[Icache.scala 58:39:@2669.4]
  reg [1:0] state; // @[Icache.scala 62:22:@2674.4]
  reg [31:0] _RAND_2;
  reg [31:0] wb_buffer_0; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_3;
  reg [31:0] wb_buffer_1; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_4;
  reg [31:0] wb_buffer_2; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_5;
  reg [31:0] wb_buffer_3; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_6;
  reg [31:0] wb_buffer_4; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_7;
  reg [31:0] wb_buffer_5; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_8;
  reg [31:0] wb_buffer_6; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_9;
  reg [31:0] wb_buffer_7; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_10;
  reg [31:0] wb_buffer_8; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_11;
  reg [31:0] wb_buffer_9; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_12;
  reg [31:0] wb_buffer_10; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_13;
  reg [31:0] wb_buffer_11; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_14;
  reg [31:0] wb_buffer_12; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_15;
  reg [31:0] wb_buffer_13; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_16;
  reg [31:0] wb_buffer_14; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_17;
  reg [31:0] wb_buffer_15; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_18;
  reg [25:0] wb_addr; // @[Icache.scala 65:20:@2676.4]
  reg [31:0] _RAND_19;
  wire  _T_78; // @[Icache.scala 67:30:@2680.4]
  wire [31:0] _T_81; // @[Cat.scala 30:58:@2683.4]
  wire  cache_hit; // @[Icache.scala 73:33:@2705.4]
  wire [25:0] _T_84; // @[Icache.scala 74:26:@2706.4]
  wire  line_hit; // @[Icache.scala 74:59:@2707.4]
  wire  _T_86; // @[Icache.scala 75:36:@2708.4]
  wire  miss; // @[Icache.scala 75:33:@2709.4]
  wire  _T_87; // @[Icache.scala 76:39:@2710.4]
  wire  _T_89; // @[Icache.scala 76:54:@2711.4]
  wire  _T_90; // @[Icache.scala 76:51:@2712.4]
  wire  pc_miss; // @[Icache.scala 76:29:@2713.4]
  wire  _T_91; // @[Icache.scala 79:50:@2714.4]
  wire  _T_92; // @[Icache.scala 79:41:@2715.4]
  wire  _T_95; // @[Icache.scala 79:62:@2717.4]
  reg  _T_99; // @[Icache.scala 27:27:@2719.4]
  reg [31:0] _RAND_20;
  wire  _GEN_1; // @[Icache.scala 29:20:@2724.6]
  wire  _GEN_2; // @[Icache.scala 28:17:@2720.4]
  wire  pc_double_miss; // @[Icache.scala 30:8:@2727.4]
  reg  _T_104; // @[Icache.scala 27:27:@2728.4]
  reg [31:0] _RAND_21;
  wire  _GEN_3; // @[Icache.scala 29:20:@2733.6]
  wire  _GEN_4; // @[Icache.scala 28:17:@2729.4]
  wire  _T_112; // @[Conditional.scala 37:30:@2743.4]
  wire [1:0] _GEN_5; // @[Icache.scala 86:22:@2745.6]
  wire  _T_113; // @[Conditional.scala 37:30:@2753.6]
  wire  _T_114; // @[Icache.scala 90:19:@2755.8]
  wire [1:0] _GEN_6; // @[Icache.scala 90:30:@2756.8]
  wire  _T_115; // @[Conditional.scala 37:30:@2764.8]
  wire [1:0] _GEN_7; // @[Icache.scala 94:29:@2766.10]
  wire [1:0] _GEN_8; // @[Conditional.scala 39:67:@2765.8]
  wire [1:0] _GEN_9; // @[Conditional.scala 39:67:@2754.6]
  wire [1:0] _GEN_10; // @[Conditional.scala 40:58:@2744.4]
  wire  _T_117; // @[Icache.scala 99:31:@2774.4]
  wire  _T_119; // @[Icache.scala 100:31:@2776.4]
  wire  _T_120; // @[Icache.scala 99:43:@2777.4]
  reg [3:0] cnt; // @[Icache.scala 103:20:@2782.4]
  reg [31:0] _RAND_22;
  reg  wb_buf_valid_0; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_23;
  reg  wb_buf_valid_1; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_24;
  reg  wb_buf_valid_2; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_25;
  reg  wb_buf_valid_3; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_26;
  reg  wb_buf_valid_4; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_27;
  reg  wb_buf_valid_5; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_28;
  reg  wb_buf_valid_6; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_29;
  reg  wb_buf_valid_7; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_30;
  reg  wb_buf_valid_8; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_31;
  reg  wb_buf_valid_9; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_32;
  reg  wb_buf_valid_10; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_33;
  reg  wb_buf_valid_11; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_34;
  reg  wb_buf_valid_12; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_35;
  reg  wb_buf_valid_13; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_36;
  reg  wb_buf_valid_14; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_37;
  reg  wb_buf_valid_15; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_38;
  wire [4:0] _T_268; // @[Icache.scala 110:18:@2820.8]
  wire [3:0] _T_269; // @[Icache.scala 110:18:@2821.8]
  wire  _GEN_12; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_13; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_14; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_15; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_16; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_17; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_18; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_19; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_20; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_21; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_22; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_23; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_24; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_25; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_26; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_27; // @[Icache.scala 111:25:@2823.8]
  wire [3:0] _GEN_28; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_29; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_30; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_31; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_32; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_33; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_34; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_35; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_36; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_37; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_38; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_39; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_40; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_41; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_42; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_43; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_44; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_45; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_46; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_47; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_48; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_49; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_50; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_51; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_52; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_53; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_54; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_55; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_56; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_57; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_58; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_59; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_60; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_62; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_63; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_64; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_65; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_66; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_67; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_68; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_69; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_70; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_71; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_72; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_73; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_74; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_75; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_76; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_77; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_78; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_79; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_80; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_81; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_82; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_83; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_84; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_85; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_86; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_87; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_88; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_89; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_90; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_91; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_92; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_93; // @[Icache.scala 105:31:@2802.4]
  wire [3:0] _GEN_94; // @[Icache.scala 105:31:@2802.4]
  wire [31:0] _GEN_95; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_96; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_97; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_98; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_99; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_100; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_101; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_102; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_103; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_104; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_105; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_106; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_107; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_108; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_109; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_110; // @[Icache.scala 118:34:@2834.6]
  wire  _T_283; // @[Icache.scala 121:27:@2837.4]
  wire  _T_284; // @[Icache.scala 121:39:@2838.4]
  wire  _T_287; // @[Icache.scala 121:52:@2841.4]
  wire  wait_inst_back; // @[Icache.scala 122:39:@2844.4]
  wire [3:0] line_idx; // @[Icache.scala 125:23:@2845.4]
  wire [31:0] _GEN_128; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_129; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_130; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_131; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_132; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_133; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_134; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_135; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_136; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_137; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_138; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_139; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_140; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_141; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_142; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] buffer_inst; // @[Icache.scala 126:24:@2846.4]
  wire  _GEN_144; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_145; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_146; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_147; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_148; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_149; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_150; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_151; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_152; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_153; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_154; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_155; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_156; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_157; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_158; // @[Icache.scala 127:78:@2847.4]
  wire  _T_294; // @[Icache.scala 127:78:@2847.4]
  reg  _T_297; // @[Icache.scala 36:27:@2848.4]
  reg [31:0] _RAND_39;
  wire  _GEN_159; // @[Icache.scala 38:20:@2853.6]
  wire  _GEN_160; // @[Icache.scala 37:17:@2849.4]
  wire  _T_300; // @[Icache.scala 39:9:@2856.4]
  wire  _T_301; // @[Icache.scala 39:22:@2857.4]
  wire  buf_inst_valid; // @[Icache.scala 127:91:@2858.4]
  CaheCore icache ( // @[Icache.scala 66:22:@2677.4]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_wen(icache_io_wen),
    .io_addr(icache_io_addr),
    .io_wdata_0(icache_io_wdata_0),
    .io_wdata_1(icache_io_wdata_1),
    .io_wdata_2(icache_io_wdata_2),
    .io_wdata_3(icache_io_wdata_3),
    .io_wdata_4(icache_io_wdata_4),
    .io_wdata_5(icache_io_wdata_5),
    .io_wdata_6(icache_io_wdata_6),
    .io_wdata_7(icache_io_wdata_7),
    .io_wdata_8(icache_io_wdata_8),
    .io_wdata_9(icache_io_wdata_9),
    .io_wdata_10(icache_io_wdata_10),
    .io_wdata_11(icache_io_wdata_11),
    .io_wdata_12(icache_io_wdata_12),
    .io_wdata_13(icache_io_wdata_13),
    .io_wdata_14(icache_io_wdata_14),
    .io_wdata_15(icache_io_wdata_15),
    .io_wstatus(icache_io_wstatus),
    .io_rdata(icache_io_rdata),
    .io_rvalid(icache_io_rvalid)
  );
  assign pc_accept = io_core_ready & io_core_pc_valid; // @[Icache.scala 58:39:@2669.4]
  assign _T_78 = state == 2'h2; // @[Icache.scala 67:30:@2680.4]
  assign _T_81 = {wb_addr,6'h0}; // @[Cat.scala 30:58:@2683.4]
  assign cache_hit = pc_valid & icache_io_rvalid; // @[Icache.scala 73:33:@2705.4]
  assign _T_84 = pc[31:6]; // @[Icache.scala 74:26:@2706.4]
  assign line_hit = _T_84 == wb_addr; // @[Icache.scala 74:59:@2707.4]
  assign _T_86 = icache_io_rvalid == 1'h0; // @[Icache.scala 75:36:@2708.4]
  assign miss = pc_valid & _T_86; // @[Icache.scala 75:33:@2709.4]
  assign _T_87 = state == 2'h0; // @[Icache.scala 76:39:@2710.4]
  assign _T_89 = line_hit == 1'h0; // @[Icache.scala 76:54:@2711.4]
  assign _T_90 = _T_87 | _T_89; // @[Icache.scala 76:51:@2712.4]
  assign pc_miss = miss & _T_90; // @[Icache.scala 76:29:@2713.4]
  assign _T_91 = state != 2'h0; // @[Icache.scala 79:50:@2714.4]
  assign _T_92 = miss & _T_91; // @[Icache.scala 79:41:@2715.4]
  assign _T_95 = _T_92 & _T_89; // @[Icache.scala 79:62:@2717.4]
  assign _GEN_1 = _T_95 ? 1'h1 : _T_99; // @[Icache.scala 29:20:@2724.6]
  assign _GEN_2 = _T_78 ? 1'h0 : _GEN_1; // @[Icache.scala 28:17:@2720.4]
  assign pc_double_miss = _T_95 | _T_99; // @[Icache.scala 30:8:@2727.4]
  assign _GEN_3 = pc_miss ? 1'h1 : _T_104; // @[Icache.scala 29:20:@2733.6]
  assign _GEN_4 = io_axi_ar_ready ? 1'h0 : _GEN_3; // @[Icache.scala 28:17:@2729.4]
  assign _T_112 = 2'h0 == state; // @[Conditional.scala 37:30:@2743.4]
  assign _GEN_5 = pc_miss ? 2'h1 : 2'h0; // @[Icache.scala 86:22:@2745.6]
  assign _T_113 = 2'h1 == state; // @[Conditional.scala 37:30:@2753.6]
  assign _T_114 = io_axi_r_last & io_axi_r_valid; // @[Icache.scala 90:19:@2755.8]
  assign _GEN_6 = _T_114 ? 2'h2 : 2'h1; // @[Icache.scala 90:30:@2756.8]
  assign _T_115 = 2'h2 == state; // @[Conditional.scala 37:30:@2764.8]
  assign _GEN_7 = pc_double_miss ? 2'h1 : 2'h0; // @[Icache.scala 94:29:@2766.10]
  assign _GEN_8 = _T_115 ? _GEN_7 : state; // @[Conditional.scala 39:67:@2765.8]
  assign _GEN_9 = _T_113 ? _GEN_6 : _GEN_8; // @[Conditional.scala 39:67:@2754.6]
  assign _GEN_10 = _T_112 ? _GEN_5 : _GEN_9; // @[Conditional.scala 40:58:@2744.4]
  assign _T_117 = _T_87 & pc_miss; // @[Icache.scala 99:31:@2774.4]
  assign _T_119 = _T_78 & pc_double_miss; // @[Icache.scala 100:31:@2776.4]
  assign _T_120 = _T_117 | _T_119; // @[Icache.scala 99:43:@2777.4]
  assign _T_268 = cnt + 4'h1; // @[Icache.scala 110:18:@2820.8]
  assign _T_269 = cnt + 4'h1; // @[Icache.scala 110:18:@2821.8]
  assign _GEN_12 = 4'h0 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_13 = 4'h1 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_14 = 4'h2 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_15 = 4'h3 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_16 = 4'h4 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_17 = 4'h5 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_18 = 4'h6 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_19 = 4'h7 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_20 = 4'h8 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_21 = 4'h9 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_22 = 4'ha == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_23 = 4'hb == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_24 = 4'hc == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_25 = 4'hd == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_26 = 4'he == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_27 = 4'hf == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_28 = io_axi_r_valid ? _T_269 : cnt; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_29 = io_axi_r_valid ? _GEN_12 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_30 = io_axi_r_valid ? _GEN_13 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_31 = io_axi_r_valid ? _GEN_14 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_32 = io_axi_r_valid ? _GEN_15 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_33 = io_axi_r_valid ? _GEN_16 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_34 = io_axi_r_valid ? _GEN_17 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_35 = io_axi_r_valid ? _GEN_18 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_36 = io_axi_r_valid ? _GEN_19 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_37 = io_axi_r_valid ? _GEN_20 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_38 = io_axi_r_valid ? _GEN_21 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_39 = io_axi_r_valid ? _GEN_22 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_40 = io_axi_r_valid ? _GEN_23 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_41 = io_axi_r_valid ? _GEN_24 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_42 = io_axi_r_valid ? _GEN_25 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_43 = io_axi_r_valid ? _GEN_26 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_44 = io_axi_r_valid ? _GEN_27 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_45 = 4'h0 == cnt ? 1'h1 : wb_buf_valid_0; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_46 = 4'h1 == cnt ? 1'h1 : wb_buf_valid_1; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_47 = 4'h2 == cnt ? 1'h1 : wb_buf_valid_2; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_48 = 4'h3 == cnt ? 1'h1 : wb_buf_valid_3; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_49 = 4'h4 == cnt ? 1'h1 : wb_buf_valid_4; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_50 = 4'h5 == cnt ? 1'h1 : wb_buf_valid_5; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_51 = 4'h6 == cnt ? 1'h1 : wb_buf_valid_6; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_52 = 4'h7 == cnt ? 1'h1 : wb_buf_valid_7; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_53 = 4'h8 == cnt ? 1'h1 : wb_buf_valid_8; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_54 = 4'h9 == cnt ? 1'h1 : wb_buf_valid_9; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_55 = 4'ha == cnt ? 1'h1 : wb_buf_valid_10; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_56 = 4'hb == cnt ? 1'h1 : wb_buf_valid_11; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_57 = 4'hc == cnt ? 1'h1 : wb_buf_valid_12; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_58 = 4'hd == cnt ? 1'h1 : wb_buf_valid_13; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_59 = 4'he == cnt ? 1'h1 : wb_buf_valid_14; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_60 = 4'hf == cnt ? 1'h1 : wb_buf_valid_15; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_62 = io_axi_r_valid ? _GEN_45 : wb_buf_valid_0; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_63 = io_axi_r_valid ? _GEN_46 : wb_buf_valid_1; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_64 = io_axi_r_valid ? _GEN_47 : wb_buf_valid_2; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_65 = io_axi_r_valid ? _GEN_48 : wb_buf_valid_3; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_66 = io_axi_r_valid ? _GEN_49 : wb_buf_valid_4; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_67 = io_axi_r_valid ? _GEN_50 : wb_buf_valid_5; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_68 = io_axi_r_valid ? _GEN_51 : wb_buf_valid_6; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_69 = io_axi_r_valid ? _GEN_52 : wb_buf_valid_7; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_70 = io_axi_r_valid ? _GEN_53 : wb_buf_valid_8; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_71 = io_axi_r_valid ? _GEN_54 : wb_buf_valid_9; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_72 = io_axi_r_valid ? _GEN_55 : wb_buf_valid_10; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_73 = io_axi_r_valid ? _GEN_56 : wb_buf_valid_11; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_74 = io_axi_r_valid ? _GEN_57 : wb_buf_valid_12; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_75 = io_axi_r_valid ? _GEN_58 : wb_buf_valid_13; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_76 = io_axi_r_valid ? _GEN_59 : wb_buf_valid_14; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_77 = io_axi_r_valid ? _GEN_60 : wb_buf_valid_15; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_78 = _T_78 ? _GEN_29 : _GEN_62; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_79 = _T_78 ? _GEN_30 : _GEN_63; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_80 = _T_78 ? _GEN_31 : _GEN_64; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_81 = _T_78 ? _GEN_32 : _GEN_65; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_82 = _T_78 ? _GEN_33 : _GEN_66; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_83 = _T_78 ? _GEN_34 : _GEN_67; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_84 = _T_78 ? _GEN_35 : _GEN_68; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_85 = _T_78 ? _GEN_36 : _GEN_69; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_86 = _T_78 ? _GEN_37 : _GEN_70; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_87 = _T_78 ? _GEN_38 : _GEN_71; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_88 = _T_78 ? _GEN_39 : _GEN_72; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_89 = _T_78 ? _GEN_40 : _GEN_73; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_90 = _T_78 ? _GEN_41 : _GEN_74; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_91 = _T_78 ? _GEN_42 : _GEN_75; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_92 = _T_78 ? _GEN_43 : _GEN_76; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_93 = _T_78 ? _GEN_44 : _GEN_77; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_94 = _T_78 ? _GEN_28 : _GEN_28; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_95 = 4'h0 == cnt ? io_axi_r_data : wb_buffer_0; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_96 = 4'h1 == cnt ? io_axi_r_data : wb_buffer_1; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_97 = 4'h2 == cnt ? io_axi_r_data : wb_buffer_2; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_98 = 4'h3 == cnt ? io_axi_r_data : wb_buffer_3; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_99 = 4'h4 == cnt ? io_axi_r_data : wb_buffer_4; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_100 = 4'h5 == cnt ? io_axi_r_data : wb_buffer_5; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_101 = 4'h6 == cnt ? io_axi_r_data : wb_buffer_6; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_102 = 4'h7 == cnt ? io_axi_r_data : wb_buffer_7; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_103 = 4'h8 == cnt ? io_axi_r_data : wb_buffer_8; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_104 = 4'h9 == cnt ? io_axi_r_data : wb_buffer_9; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_105 = 4'ha == cnt ? io_axi_r_data : wb_buffer_10; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_106 = 4'hb == cnt ? io_axi_r_data : wb_buffer_11; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_107 = 4'hc == cnt ? io_axi_r_data : wb_buffer_12; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_108 = 4'hd == cnt ? io_axi_r_data : wb_buffer_13; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_109 = 4'he == cnt ? io_axi_r_data : wb_buffer_14; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_110 = 4'hf == cnt ? io_axi_r_data : wb_buffer_15; // @[Icache.scala 118:34:@2834.6]
  assign _T_283 = _T_91 & pc_valid; // @[Icache.scala 121:27:@2837.4]
  assign _T_284 = _T_283 & line_hit; // @[Icache.scala 121:39:@2838.4]
  assign _T_287 = _T_284 | _T_117; // @[Icache.scala 121:52:@2841.4]
  assign wait_inst_back = _T_287 | _T_119; // @[Icache.scala 122:39:@2844.4]
  assign line_idx = pc[5:2]; // @[Icache.scala 125:23:@2845.4]
  assign _GEN_128 = 4'h1 == line_idx ? wb_buffer_1 : wb_buffer_0; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_129 = 4'h2 == line_idx ? wb_buffer_2 : _GEN_128; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_130 = 4'h3 == line_idx ? wb_buffer_3 : _GEN_129; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_131 = 4'h4 == line_idx ? wb_buffer_4 : _GEN_130; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_132 = 4'h5 == line_idx ? wb_buffer_5 : _GEN_131; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_133 = 4'h6 == line_idx ? wb_buffer_6 : _GEN_132; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_134 = 4'h7 == line_idx ? wb_buffer_7 : _GEN_133; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_135 = 4'h8 == line_idx ? wb_buffer_8 : _GEN_134; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_136 = 4'h9 == line_idx ? wb_buffer_9 : _GEN_135; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_137 = 4'ha == line_idx ? wb_buffer_10 : _GEN_136; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_138 = 4'hb == line_idx ? wb_buffer_11 : _GEN_137; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_139 = 4'hc == line_idx ? wb_buffer_12 : _GEN_138; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_140 = 4'hd == line_idx ? wb_buffer_13 : _GEN_139; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_141 = 4'he == line_idx ? wb_buffer_14 : _GEN_140; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_142 = 4'hf == line_idx ? wb_buffer_15 : _GEN_141; // @[Icache.scala 126:24:@2846.4]
  assign buffer_inst = line_hit ? _GEN_142 : icache_io_rdata; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_144 = 4'h1 == line_idx ? wb_buf_valid_1 : wb_buf_valid_0; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_145 = 4'h2 == line_idx ? wb_buf_valid_2 : _GEN_144; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_146 = 4'h3 == line_idx ? wb_buf_valid_3 : _GEN_145; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_147 = 4'h4 == line_idx ? wb_buf_valid_4 : _GEN_146; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_148 = 4'h5 == line_idx ? wb_buf_valid_5 : _GEN_147; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_149 = 4'h6 == line_idx ? wb_buf_valid_6 : _GEN_148; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_150 = 4'h7 == line_idx ? wb_buf_valid_7 : _GEN_149; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_151 = 4'h8 == line_idx ? wb_buf_valid_8 : _GEN_150; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_152 = 4'h9 == line_idx ? wb_buf_valid_9 : _GEN_151; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_153 = 4'ha == line_idx ? wb_buf_valid_10 : _GEN_152; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_154 = 4'hb == line_idx ? wb_buf_valid_11 : _GEN_153; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_155 = 4'hc == line_idx ? wb_buf_valid_12 : _GEN_154; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_156 = 4'hd == line_idx ? wb_buf_valid_13 : _GEN_155; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_157 = 4'he == line_idx ? wb_buf_valid_14 : _GEN_156; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_158 = 4'hf == line_idx ? wb_buf_valid_15 : _GEN_157; // @[Icache.scala 127:78:@2847.4]
  assign _T_294 = _GEN_158 & line_hit; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_159 = wait_inst_back ? 1'h1 : _T_297; // @[Icache.scala 38:20:@2853.6]
  assign _GEN_160 = _T_294 ? 1'h0 : _GEN_159; // @[Icache.scala 37:17:@2849.4]
  assign _T_300 = wait_inst_back | _T_297; // @[Icache.scala 39:9:@2856.4]
  assign _T_301 = _T_300 & _T_294; // @[Icache.scala 39:22:@2857.4]
  assign buf_inst_valid = _T_301 | cache_hit; // @[Icache.scala 127:91:@2858.4]
  assign io_core_inst_valid = _T_87 ? cache_hit : buf_inst_valid; // @[Icache.scala 128:22:@2861.4]
  assign io_core_inst_bits = _T_87 ? icache_io_rdata : buffer_inst; // @[Icache.scala 129:22:@2864.4]
  assign io_core_ready = state != 2'h2; // @[Icache.scala 82:19:@2742.4]
  assign io_axi_ar_valid = pc_miss | _T_104; // @[Icache.scala 80:19:@2737.4]
  assign io_axi_ar_addr = {_T_84,6'h0}; // @[Icache.scala 81:19:@2740.4]
  assign icache_clock = clock; // @[:@2678.4]
  assign icache_reset = reset; // @[:@2679.4]
  assign icache_io_wen = state == 2'h2; // @[Icache.scala 67:21:@2681.4]
  assign icache_io_addr = _T_78 ? _T_81 : io_core_pc_bits; // @[Icache.scala 68:21:@2685.4]
  assign icache_io_wdata_0 = wb_buffer_0; // @[Icache.scala 69:21:@2686.4]
  assign icache_io_wdata_1 = wb_buffer_1; // @[Icache.scala 69:21:@2687.4]
  assign icache_io_wdata_2 = wb_buffer_2; // @[Icache.scala 69:21:@2688.4]
  assign icache_io_wdata_3 = wb_buffer_3; // @[Icache.scala 69:21:@2689.4]
  assign icache_io_wdata_4 = wb_buffer_4; // @[Icache.scala 69:21:@2690.4]
  assign icache_io_wdata_5 = wb_buffer_5; // @[Icache.scala 69:21:@2691.4]
  assign icache_io_wdata_6 = wb_buffer_6; // @[Icache.scala 69:21:@2692.4]
  assign icache_io_wdata_7 = wb_buffer_7; // @[Icache.scala 69:21:@2693.4]
  assign icache_io_wdata_8 = wb_buffer_8; // @[Icache.scala 69:21:@2694.4]
  assign icache_io_wdata_9 = wb_buffer_9; // @[Icache.scala 69:21:@2695.4]
  assign icache_io_wdata_10 = wb_buffer_10; // @[Icache.scala 69:21:@2696.4]
  assign icache_io_wdata_11 = wb_buffer_11; // @[Icache.scala 69:21:@2697.4]
  assign icache_io_wdata_12 = wb_buffer_12; // @[Icache.scala 69:21:@2698.4]
  assign icache_io_wdata_13 = wb_buffer_13; // @[Icache.scala 69:21:@2699.4]
  assign icache_io_wdata_14 = wb_buffer_14; // @[Icache.scala 69:21:@2700.4]
  assign icache_io_wdata_15 = wb_buffer_15; // @[Icache.scala 69:21:@2701.4]
  assign icache_io_wstatus = state == 2'h2; // @[Icache.scala 70:21:@2703.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wb_buffer_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  wb_buffer_1 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  wb_buffer_2 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  wb_buffer_3 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wb_buffer_4 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wb_buffer_5 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wb_buffer_6 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wb_buffer_7 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wb_buffer_8 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wb_buffer_9 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wb_buffer_10 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wb_buffer_11 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wb_buffer_12 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wb_buffer_13 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wb_buffer_14 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wb_buffer_15 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wb_addr = _RAND_19[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_99 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_104 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  cnt = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  wb_buf_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wb_buf_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  wb_buf_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  wb_buf_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  wb_buf_valid_4 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  wb_buf_valid_5 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  wb_buf_valid_6 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  wb_buf_valid_7 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  wb_buf_valid_8 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  wb_buf_valid_9 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_buf_valid_10 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wb_buf_valid_11 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wb_buf_valid_12 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wb_buf_valid_13 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wb_buf_valid_14 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wb_buf_valid_15 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_297 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc_valid <= 1'h0;
    end else begin
      pc_valid <= pc_accept;
    end
    if (pc_accept) begin
      pc <= io_core_pc_bits;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_112) begin
        if (pc_miss) begin
          state <= 2'h1;
        end else begin
          state <= 2'h0;
        end
      end else begin
        if (_T_113) begin
          if (_T_114) begin
            state <= 2'h2;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_115) begin
            if (pc_double_miss) begin
              state <= 2'h1;
            end else begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    if (io_axi_r_valid) begin
      if (4'h0 == cnt) begin
        wb_buffer_0 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h1 == cnt) begin
        wb_buffer_1 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h2 == cnt) begin
        wb_buffer_2 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h3 == cnt) begin
        wb_buffer_3 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h4 == cnt) begin
        wb_buffer_4 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h5 == cnt) begin
        wb_buffer_5 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h6 == cnt) begin
        wb_buffer_6 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h7 == cnt) begin
        wb_buffer_7 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h8 == cnt) begin
        wb_buffer_8 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h9 == cnt) begin
        wb_buffer_9 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'ha == cnt) begin
        wb_buffer_10 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hb == cnt) begin
        wb_buffer_11 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hc == cnt) begin
        wb_buffer_12 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hd == cnt) begin
        wb_buffer_13 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'he == cnt) begin
        wb_buffer_14 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hf == cnt) begin
        wb_buffer_15 <= io_axi_r_data;
      end
    end
    if (_T_120) begin
      wb_addr <= _T_84;
    end
    if (reset) begin
      _T_99 <= 1'h0;
    end else begin
      if (_T_78) begin
        _T_99 <= 1'h0;
      end else begin
        if (_T_95) begin
          _T_99 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_104 <= 1'h0;
    end else begin
      if (io_axi_ar_ready) begin
        _T_104 <= 1'h0;
      end else begin
        if (pc_miss) begin
          _T_104 <= 1'h1;
        end
      end
    end
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          cnt <= _T_269;
        end
      end else begin
        if (io_axi_r_valid) begin
          cnt <= _T_269;
        end
      end
    end
    if (reset) begin
      wb_buf_valid_0 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_0 <= _GEN_12;
        end else begin
          wb_buf_valid_0 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h0 == cnt) begin
            wb_buf_valid_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_1 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_1 <= _GEN_13;
        end else begin
          wb_buf_valid_1 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h1 == cnt) begin
            wb_buf_valid_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_2 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_2 <= _GEN_14;
        end else begin
          wb_buf_valid_2 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h2 == cnt) begin
            wb_buf_valid_2 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_3 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_3 <= _GEN_15;
        end else begin
          wb_buf_valid_3 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h3 == cnt) begin
            wb_buf_valid_3 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_4 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_4 <= _GEN_16;
        end else begin
          wb_buf_valid_4 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h4 == cnt) begin
            wb_buf_valid_4 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_5 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_5 <= _GEN_17;
        end else begin
          wb_buf_valid_5 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h5 == cnt) begin
            wb_buf_valid_5 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_6 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_6 <= _GEN_18;
        end else begin
          wb_buf_valid_6 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h6 == cnt) begin
            wb_buf_valid_6 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_7 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_7 <= _GEN_19;
        end else begin
          wb_buf_valid_7 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h7 == cnt) begin
            wb_buf_valid_7 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_8 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_8 <= _GEN_20;
        end else begin
          wb_buf_valid_8 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h8 == cnt) begin
            wb_buf_valid_8 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_9 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_9 <= _GEN_21;
        end else begin
          wb_buf_valid_9 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h9 == cnt) begin
            wb_buf_valid_9 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_10 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_10 <= _GEN_22;
        end else begin
          wb_buf_valid_10 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'ha == cnt) begin
            wb_buf_valid_10 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_11 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_11 <= _GEN_23;
        end else begin
          wb_buf_valid_11 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hb == cnt) begin
            wb_buf_valid_11 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_12 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_12 <= _GEN_24;
        end else begin
          wb_buf_valid_12 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hc == cnt) begin
            wb_buf_valid_12 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_13 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_13 <= _GEN_25;
        end else begin
          wb_buf_valid_13 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hd == cnt) begin
            wb_buf_valid_13 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_14 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_14 <= _GEN_26;
        end else begin
          wb_buf_valid_14 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'he == cnt) begin
            wb_buf_valid_14 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_15 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_15 <= _GEN_27;
        end else begin
          wb_buf_valid_15 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hf == cnt) begin
            wb_buf_valid_15 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_297 <= 1'h0;
    end else begin
      if (_T_294) begin
        _T_297 <= 1'h0;
      end else begin
        if (wait_inst_back) begin
          _T_297 <= 1'h1;
        end
      end
    end
  end
endmodule