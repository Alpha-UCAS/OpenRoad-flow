module RAS( // @[:@709.2]
  input         clock, // @[:@710.4]
  input         reset, // @[:@711.4]
  input         io_push_valid, // @[:@712.4]
  input  [31:0] io_push_bits, // @[:@712.4]
  input         io_pop, // @[:@712.4]
  output [31:0] io_peek // @[:@712.4]
);
  reg [31:0] stack [0:7]; // @[RAS.scala 13:18:@714.4]
  reg [31:0] _RAND_0;
  wire [31:0] stack__T_23_data; // @[RAS.scala 13:18:@714.4]
  wire [2:0] stack__T_23_addr; // @[RAS.scala 13:18:@714.4]
  wire [31:0] stack__T_24_data; // @[RAS.scala 13:18:@714.4]
  wire [2:0] stack__T_24_addr; // @[RAS.scala 13:18:@714.4]
  wire  stack__T_24_mask; // @[RAS.scala 13:18:@714.4]
  wire  stack__T_24_en; // @[RAS.scala 13:18:@714.4]
  wire [31:0] stack__T_25_data; // @[RAS.scala 13:18:@714.4]
  wire [2:0] stack__T_25_addr; // @[RAS.scala 13:18:@714.4]
  wire  stack__T_25_mask; // @[RAS.scala 13:18:@714.4]
  wire  stack__T_25_en; // @[RAS.scala 13:18:@714.4]
  reg [2:0] pos; // @[RAS.scala 14:22:@715.4]
  reg [31:0] _RAND_1;
  reg [2:0] next; // @[RAS.scala 15:22:@716.4]
  reg [31:0] _RAND_2;
  wire  _GEN_7; // @[RAS.scala 19:18:@720.6]
  wire  _T_27; // @[RAS.scala 26:26:@729.4]
  wire  _T_28; // @[RAS.scala 26:23:@730.4]
  wire [3:0] _T_30; // @[RAS.scala 27:18:@732.6]
  wire [2:0] _T_31; // @[RAS.scala 27:18:@733.6]
  wire [3:0] _T_33; // @[RAS.scala 28:18:@735.6]
  wire [2:0] _T_34; // @[RAS.scala 28:18:@736.6]
  wire [3:0] _T_36; // @[RAS.scala 31:18:@741.8]
  wire [3:0] _T_37; // @[RAS.scala 31:18:@742.8]
  wire [2:0] _T_38; // @[RAS.scala 31:18:@743.8]
  wire [3:0] _T_40; // @[RAS.scala 32:18:@745.8]
  wire [3:0] _T_41; // @[RAS.scala 32:18:@746.8]
  wire [2:0] _T_42; // @[RAS.scala 32:18:@747.8]
  wire [2:0] _GEN_20; // @[RAS.scala 29:22:@740.6]
  wire [2:0] _GEN_21; // @[RAS.scala 29:22:@740.6]
  wire [2:0] _GEN_22; // @[RAS.scala 26:35:@731.4]
  wire [2:0] _GEN_23; // @[RAS.scala 26:35:@731.4]
  assign stack__T_23_addr = pos;
  assign stack__T_23_data = stack[stack__T_23_addr]; // @[RAS.scala 13:18:@714.4]
  assign stack__T_24_data = io_push_bits;
  assign stack__T_24_addr = pos;
  assign stack__T_24_mask = 1'h1;
  assign stack__T_24_en = io_push_valid ? io_pop : 1'h0;
  assign stack__T_25_data = io_push_bits;
  assign stack__T_25_addr = next;
  assign stack__T_25_mask = 1'h1;
  assign stack__T_25_en = io_push_valid ? _GEN_7 : 1'h0;
  assign _GEN_7 = io_pop ? 1'h0 : 1'h1; // @[RAS.scala 19:18:@720.6]
  assign _T_27 = io_pop == 1'h0; // @[RAS.scala 26:26:@729.4]
  assign _T_28 = io_push_valid & _T_27; // @[RAS.scala 26:23:@730.4]
  assign _T_30 = pos + 3'h1; // @[RAS.scala 27:18:@732.6]
  assign _T_31 = pos + 3'h1; // @[RAS.scala 27:18:@733.6]
  assign _T_33 = next + 3'h1; // @[RAS.scala 28:18:@735.6]
  assign _T_34 = next + 3'h1; // @[RAS.scala 28:18:@736.6]
  assign _T_36 = pos - 3'h1; // @[RAS.scala 31:18:@741.8]
  assign _T_37 = $unsigned(_T_36); // @[RAS.scala 31:18:@742.8]
  assign _T_38 = _T_37[2:0]; // @[RAS.scala 31:18:@743.8]
  assign _T_40 = next - 3'h1; // @[RAS.scala 32:18:@745.8]
  assign _T_41 = $unsigned(_T_40); // @[RAS.scala 32:18:@746.8]
  assign _T_42 = _T_41[2:0]; // @[RAS.scala 32:18:@747.8]
  assign _GEN_20 = io_pop ? _T_38 : pos; // @[RAS.scala 29:22:@740.6]
  assign _GEN_21 = io_pop ? _T_42 : next; // @[RAS.scala 29:22:@740.6]
  assign _GEN_22 = _T_28 ? _T_31 : _GEN_20; // @[RAS.scala 26:35:@731.4]
  assign _GEN_23 = _T_28 ? _T_34 : _GEN_21; // @[RAS.scala 26:35:@731.4]
  assign io_peek = stack__T_23_data; // @[RAS.scala 16:11:@718.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 8; initvar = initvar+1)
    stack[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pos = _RAND_1[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  next = _RAND_2[2:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(stack__T_24_en & stack__T_24_mask) begin
      stack[stack__T_24_addr] <= stack__T_24_data; // @[RAS.scala 13:18:@714.4]
    end
    if(stack__T_25_en & stack__T_25_mask) begin
      stack[stack__T_25_addr] <= stack__T_25_data; // @[RAS.scala 13:18:@714.4]
    end
    if (reset) begin
      pos <= 3'h7;
    end else begin
      if (_T_28) begin
        pos <= _T_31;
      end else begin
        if (io_pop) begin
          pos <= _T_38;
        end
      end
    end
    if (reset) begin
      next <= 3'h0;
    end else begin
      if (_T_28) begin
        next <= _T_34;
      end else begin
        if (io_pop) begin
          next <= _T_42;
        end
      end
    end
  end
endmodule
module BTB( // @[:@751.2]
  input         clock, // @[:@752.4]
  input         reset, // @[:@753.4]
  input         io_if_pc_valid, // @[:@754.4]
  input  [31:0] io_if_pc_bits, // @[:@754.4]
  output        io_predict_0_redirect, // @[:@754.4]
  output [9:0]  io_predict_0_history, // @[:@754.4]
  output        io_predict_0_diff, // @[:@754.4]
  output [31:0] io_predict_0_tgt, // @[:@754.4]
  output        io_predict_1_redirect, // @[:@754.4]
  output [9:0]  io_predict_1_history, // @[:@754.4]
  output        io_predict_1_diff, // @[:@754.4]
  output [31:0] io_predict_1_tgt, // @[:@754.4]
  output        io_split, // @[:@754.4]
  input         io_branch, // @[:@754.4]
  input         io_ras_pop, // @[:@754.4]
  input         io_ras_push_valid, // @[:@754.4]
  input  [31:0] io_ras_push_bits, // @[:@754.4]
  input         io_fb_pc_valid, // @[:@754.4]
  input  [31:0] io_fb_pc_bits, // @[:@754.4]
  input  [1:0]  io_fb_type, // @[:@754.4]
  input         io_feedBack_redirect, // @[:@754.4]
  input  [9:0]  io_feedBack_history, // @[:@754.4]
  input         io_feedBack_diff, // @[:@754.4]
  input  [31:0] io_feedBack_tgt, // @[:@754.4]
  input         io_feedBack_valid, // @[:@754.4]
  input  [31:0] io_cyc // @[:@754.4]
);
  reg [1:0] bht [0:1023]; // @[BTB.scala 77:16:@757.4]
  reg [31:0] _RAND_0;
  wire [1:0] bht__T_1239_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_1239_addr; // @[BTB.scala 77:16:@757.4]
  wire [1:0] bht__T_2316_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_2316_addr; // @[BTB.scala 77:16:@757.4]
  wire [1:0] bht__T_2923_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_2923_addr; // @[BTB.scala 77:16:@757.4]
  wire [1:0] bht__T_3298_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_3298_addr; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3298_mask; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3298_en; // @[BTB.scala 77:16:@757.4]
  wire [1:0] bht__T_3316_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_3316_addr; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3316_mask; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3316_en; // @[BTB.scala 77:16:@757.4]
  wire [1:0] bht__T_3327_data; // @[BTB.scala 77:16:@757.4]
  wire [9:0] bht__T_3327_addr; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3327_mask; // @[BTB.scala 77:16:@757.4]
  wire  bht__T_3327_en; // @[BTB.scala 77:16:@757.4]
  reg  arb [0:1023]; // @[BTB.scala 78:16:@758.4]
  reg [31:0] _RAND_1;
  wire  arb__T_1238_data; // @[BTB.scala 78:16:@758.4]
  wire [9:0] arb__T_1238_addr; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_2315_data; // @[BTB.scala 78:16:@758.4]
  wire [9:0] arb__T_2315_addr; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3280_data; // @[BTB.scala 78:16:@758.4]
  wire [9:0] arb__T_3280_addr; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3335_data; // @[BTB.scala 78:16:@758.4]
  wire [9:0] arb__T_3335_addr; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3335_mask; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3335_en; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3337_data; // @[BTB.scala 78:16:@758.4]
  wire [9:0] arb__T_3337_addr; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3337_mask; // @[BTB.scala 78:16:@758.4]
  wire  arb__T_3337_en; // @[BTB.scala 78:16:@758.4]
  wire  RAS_clock; // @[BTB.scala 79:19:@759.4]
  wire  RAS_reset; // @[BTB.scala 79:19:@759.4]
  wire  RAS_io_push_valid; // @[BTB.scala 79:19:@759.4]
  wire [31:0] RAS_io_push_bits; // @[BTB.scala 79:19:@759.4]
  wire  RAS_io_pop; // @[BTB.scala 79:19:@759.4]
  wire [31:0] RAS_io_peek; // @[BTB.scala 79:19:@759.4]
  reg [9:0] gb_history; // @[BTB.scala 76:27:@756.4]
  reg [31:0] _RAND_2;
  reg  btb_valid_0; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_3;
  reg  btb_valid_1; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_4;
  reg  btb_valid_2; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_5;
  reg  btb_valid_3; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_6;
  reg  btb_valid_4; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_7;
  reg  btb_valid_5; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_8;
  reg  btb_valid_6; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_9;
  reg  btb_valid_7; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_10;
  reg  btb_valid_8; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_11;
  reg  btb_valid_9; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_12;
  reg  btb_valid_10; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_13;
  reg  btb_valid_11; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_14;
  reg  btb_valid_12; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_15;
  reg  btb_valid_13; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_16;
  reg  btb_valid_14; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_17;
  reg  btb_valid_15; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_18;
  reg  btb_valid_16; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_19;
  reg  btb_valid_17; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_20;
  reg  btb_valid_18; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_21;
  reg  btb_valid_19; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_22;
  reg  btb_valid_20; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_23;
  reg  btb_valid_21; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_24;
  reg  btb_valid_22; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_25;
  reg  btb_valid_23; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_26;
  reg  btb_valid_24; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_27;
  reg  btb_valid_25; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_28;
  reg  btb_valid_26; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_29;
  reg  btb_valid_27; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_30;
  reg  btb_valid_28; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_31;
  reg  btb_valid_29; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_32;
  reg  btb_valid_30; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_33;
  reg  btb_valid_31; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_34;
  reg  btb_valid_32; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_35;
  reg  btb_valid_33; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_36;
  reg  btb_valid_34; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_37;
  reg  btb_valid_35; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_38;
  reg  btb_valid_36; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_39;
  reg  btb_valid_37; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_40;
  reg  btb_valid_38; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_41;
  reg  btb_valid_39; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_42;
  reg  btb_valid_40; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_43;
  reg  btb_valid_41; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_44;
  reg  btb_valid_42; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_45;
  reg  btb_valid_43; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_46;
  reg  btb_valid_44; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_47;
  reg  btb_valid_45; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_48;
  reg  btb_valid_46; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_49;
  reg  btb_valid_47; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_50;
  reg  btb_valid_48; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_51;
  reg  btb_valid_49; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_52;
  reg  btb_valid_50; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_53;
  reg  btb_valid_51; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_54;
  reg  btb_valid_52; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_55;
  reg  btb_valid_53; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_56;
  reg  btb_valid_54; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_57;
  reg  btb_valid_55; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_58;
  reg  btb_valid_56; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_59;
  reg  btb_valid_57; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_60;
  reg  btb_valid_58; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_61;
  reg  btb_valid_59; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_62;
  reg  btb_valid_60; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_63;
  reg  btb_valid_61; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_64;
  reg  btb_valid_62; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_65;
  reg  btb_valid_63; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_66;
  reg [29:0] btb_pc_0; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_67;
  reg [29:0] btb_pc_1; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_68;
  reg [29:0] btb_pc_2; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_69;
  reg [29:0] btb_pc_3; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_70;
  reg [29:0] btb_pc_4; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_71;
  reg [29:0] btb_pc_5; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_72;
  reg [29:0] btb_pc_6; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_73;
  reg [29:0] btb_pc_7; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_74;
  reg [29:0] btb_pc_8; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_75;
  reg [29:0] btb_pc_9; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_76;
  reg [29:0] btb_pc_10; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_77;
  reg [29:0] btb_pc_11; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_78;
  reg [29:0] btb_pc_12; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_79;
  reg [29:0] btb_pc_13; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_80;
  reg [29:0] btb_pc_14; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_81;
  reg [29:0] btb_pc_15; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_82;
  reg [29:0] btb_pc_16; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_83;
  reg [29:0] btb_pc_17; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_84;
  reg [29:0] btb_pc_18; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_85;
  reg [29:0] btb_pc_19; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_86;
  reg [29:0] btb_pc_20; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_87;
  reg [29:0] btb_pc_21; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_88;
  reg [29:0] btb_pc_22; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_89;
  reg [29:0] btb_pc_23; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_90;
  reg [29:0] btb_pc_24; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_91;
  reg [29:0] btb_pc_25; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_92;
  reg [29:0] btb_pc_26; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_93;
  reg [29:0] btb_pc_27; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_94;
  reg [29:0] btb_pc_28; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_95;
  reg [29:0] btb_pc_29; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_96;
  reg [29:0] btb_pc_30; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_97;
  reg [29:0] btb_pc_31; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_98;
  reg [29:0] btb_pc_32; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_99;
  reg [29:0] btb_pc_33; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_100;
  reg [29:0] btb_pc_34; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_101;
  reg [29:0] btb_pc_35; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_102;
  reg [29:0] btb_pc_36; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_103;
  reg [29:0] btb_pc_37; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_104;
  reg [29:0] btb_pc_38; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_105;
  reg [29:0] btb_pc_39; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_106;
  reg [29:0] btb_pc_40; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_107;
  reg [29:0] btb_pc_41; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_108;
  reg [29:0] btb_pc_42; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_109;
  reg [29:0] btb_pc_43; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_110;
  reg [29:0] btb_pc_44; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_111;
  reg [29:0] btb_pc_45; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_112;
  reg [29:0] btb_pc_46; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_113;
  reg [29:0] btb_pc_47; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_114;
  reg [29:0] btb_pc_48; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_115;
  reg [29:0] btb_pc_49; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_116;
  reg [29:0] btb_pc_50; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_117;
  reg [29:0] btb_pc_51; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_118;
  reg [29:0] btb_pc_52; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_119;
  reg [29:0] btb_pc_53; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_120;
  reg [29:0] btb_pc_54; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_121;
  reg [29:0] btb_pc_55; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_122;
  reg [29:0] btb_pc_56; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_123;
  reg [29:0] btb_pc_57; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_124;
  reg [29:0] btb_pc_58; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_125;
  reg [29:0] btb_pc_59; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_126;
  reg [29:0] btb_pc_60; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_127;
  reg [29:0] btb_pc_61; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_128;
  reg [29:0] btb_pc_62; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_129;
  reg [29:0] btb_pc_63; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_130;
  reg [29:0] btb_tgt_0; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_131;
  reg [29:0] btb_tgt_1; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_132;
  reg [29:0] btb_tgt_2; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_133;
  reg [29:0] btb_tgt_3; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_134;
  reg [29:0] btb_tgt_4; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_135;
  reg [29:0] btb_tgt_5; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_136;
  reg [29:0] btb_tgt_6; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_137;
  reg [29:0] btb_tgt_7; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_138;
  reg [29:0] btb_tgt_8; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_139;
  reg [29:0] btb_tgt_9; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_140;
  reg [29:0] btb_tgt_10; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_141;
  reg [29:0] btb_tgt_11; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_142;
  reg [29:0] btb_tgt_12; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_143;
  reg [29:0] btb_tgt_13; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_144;
  reg [29:0] btb_tgt_14; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_145;
  reg [29:0] btb_tgt_15; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_146;
  reg [29:0] btb_tgt_16; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_147;
  reg [29:0] btb_tgt_17; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_148;
  reg [29:0] btb_tgt_18; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_149;
  reg [29:0] btb_tgt_19; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_150;
  reg [29:0] btb_tgt_20; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_151;
  reg [29:0] btb_tgt_21; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_152;
  reg [29:0] btb_tgt_22; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_153;
  reg [29:0] btb_tgt_23; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_154;
  reg [29:0] btb_tgt_24; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_155;
  reg [29:0] btb_tgt_25; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_156;
  reg [29:0] btb_tgt_26; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_157;
  reg [29:0] btb_tgt_27; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_158;
  reg [29:0] btb_tgt_28; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_159;
  reg [29:0] btb_tgt_29; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_160;
  reg [29:0] btb_tgt_30; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_161;
  reg [29:0] btb_tgt_31; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_162;
  reg [29:0] btb_tgt_32; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_163;
  reg [29:0] btb_tgt_33; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_164;
  reg [29:0] btb_tgt_34; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_165;
  reg [29:0] btb_tgt_35; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_166;
  reg [29:0] btb_tgt_36; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_167;
  reg [29:0] btb_tgt_37; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_168;
  reg [29:0] btb_tgt_38; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_169;
  reg [29:0] btb_tgt_39; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_170;
  reg [29:0] btb_tgt_40; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_171;
  reg [29:0] btb_tgt_41; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_172;
  reg [29:0] btb_tgt_42; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_173;
  reg [29:0] btb_tgt_43; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_174;
  reg [29:0] btb_tgt_44; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_175;
  reg [29:0] btb_tgt_45; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_176;
  reg [29:0] btb_tgt_46; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_177;
  reg [29:0] btb_tgt_47; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_178;
  reg [29:0] btb_tgt_48; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_179;
  reg [29:0] btb_tgt_49; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_180;
  reg [29:0] btb_tgt_50; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_181;
  reg [29:0] btb_tgt_51; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_182;
  reg [29:0] btb_tgt_52; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_183;
  reg [29:0] btb_tgt_53; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_184;
  reg [29:0] btb_tgt_54; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_185;
  reg [29:0] btb_tgt_55; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_186;
  reg [29:0] btb_tgt_56; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_187;
  reg [29:0] btb_tgt_57; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_188;
  reg [29:0] btb_tgt_58; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_189;
  reg [29:0] btb_tgt_59; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_190;
  reg [29:0] btb_tgt_60; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_191;
  reg [29:0] btb_tgt_61; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_192;
  reg [29:0] btb_tgt_62; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_193;
  reg [29:0] btb_tgt_63; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_194;
  reg [1:0] btb_bj_type_0; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_195;
  reg [1:0] btb_bj_type_1; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_196;
  reg [1:0] btb_bj_type_2; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_197;
  reg [1:0] btb_bj_type_3; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_198;
  reg [1:0] btb_bj_type_4; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_199;
  reg [1:0] btb_bj_type_5; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_200;
  reg [1:0] btb_bj_type_6; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_201;
  reg [1:0] btb_bj_type_7; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_202;
  reg [1:0] btb_bj_type_8; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_203;
  reg [1:0] btb_bj_type_9; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_204;
  reg [1:0] btb_bj_type_10; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_205;
  reg [1:0] btb_bj_type_11; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_206;
  reg [1:0] btb_bj_type_12; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_207;
  reg [1:0] btb_bj_type_13; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_208;
  reg [1:0] btb_bj_type_14; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_209;
  reg [1:0] btb_bj_type_15; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_210;
  reg [1:0] btb_bj_type_16; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_211;
  reg [1:0] btb_bj_type_17; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_212;
  reg [1:0] btb_bj_type_18; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_213;
  reg [1:0] btb_bj_type_19; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_214;
  reg [1:0] btb_bj_type_20; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_215;
  reg [1:0] btb_bj_type_21; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_216;
  reg [1:0] btb_bj_type_22; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_217;
  reg [1:0] btb_bj_type_23; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_218;
  reg [1:0] btb_bj_type_24; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_219;
  reg [1:0] btb_bj_type_25; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_220;
  reg [1:0] btb_bj_type_26; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_221;
  reg [1:0] btb_bj_type_27; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_222;
  reg [1:0] btb_bj_type_28; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_223;
  reg [1:0] btb_bj_type_29; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_224;
  reg [1:0] btb_bj_type_30; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_225;
  reg [1:0] btb_bj_type_31; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_226;
  reg [1:0] btb_bj_type_32; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_227;
  reg [1:0] btb_bj_type_33; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_228;
  reg [1:0] btb_bj_type_34; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_229;
  reg [1:0] btb_bj_type_35; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_230;
  reg [1:0] btb_bj_type_36; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_231;
  reg [1:0] btb_bj_type_37; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_232;
  reg [1:0] btb_bj_type_38; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_233;
  reg [1:0] btb_bj_type_39; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_234;
  reg [1:0] btb_bj_type_40; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_235;
  reg [1:0] btb_bj_type_41; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_236;
  reg [1:0] btb_bj_type_42; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_237;
  reg [1:0] btb_bj_type_43; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_238;
  reg [1:0] btb_bj_type_44; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_239;
  reg [1:0] btb_bj_type_45; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_240;
  reg [1:0] btb_bj_type_46; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_241;
  reg [1:0] btb_bj_type_47; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_242;
  reg [1:0] btb_bj_type_48; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_243;
  reg [1:0] btb_bj_type_49; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_244;
  reg [1:0] btb_bj_type_50; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_245;
  reg [1:0] btb_bj_type_51; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_246;
  reg [1:0] btb_bj_type_52; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_247;
  reg [1:0] btb_bj_type_53; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_248;
  reg [1:0] btb_bj_type_54; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_249;
  reg [1:0] btb_bj_type_55; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_250;
  reg [1:0] btb_bj_type_56; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_251;
  reg [1:0] btb_bj_type_57; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_252;
  reg [1:0] btb_bj_type_58; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_253;
  reg [1:0] btb_bj_type_59; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_254;
  reg [1:0] btb_bj_type_60; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_255;
  reg [1:0] btb_bj_type_61; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_256;
  reg [1:0] btb_bj_type_62; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_257;
  reg [1:0] btb_bj_type_63; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_258;
  reg [1:0] btb_h_count_0; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_259;
  reg [1:0] btb_h_count_1; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_260;
  reg [1:0] btb_h_count_2; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_261;
  reg [1:0] btb_h_count_3; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_262;
  reg [1:0] btb_h_count_4; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_263;
  reg [1:0] btb_h_count_5; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_264;
  reg [1:0] btb_h_count_6; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_265;
  reg [1:0] btb_h_count_7; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_266;
  reg [1:0] btb_h_count_8; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_267;
  reg [1:0] btb_h_count_9; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_268;
  reg [1:0] btb_h_count_10; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_269;
  reg [1:0] btb_h_count_11; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_270;
  reg [1:0] btb_h_count_12; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_271;
  reg [1:0] btb_h_count_13; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_272;
  reg [1:0] btb_h_count_14; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_273;
  reg [1:0] btb_h_count_15; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_274;
  reg [1:0] btb_h_count_16; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_275;
  reg [1:0] btb_h_count_17; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_276;
  reg [1:0] btb_h_count_18; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_277;
  reg [1:0] btb_h_count_19; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_278;
  reg [1:0] btb_h_count_20; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_279;
  reg [1:0] btb_h_count_21; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_280;
  reg [1:0] btb_h_count_22; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_281;
  reg [1:0] btb_h_count_23; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_282;
  reg [1:0] btb_h_count_24; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_283;
  reg [1:0] btb_h_count_25; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_284;
  reg [1:0] btb_h_count_26; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_285;
  reg [1:0] btb_h_count_27; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_286;
  reg [1:0] btb_h_count_28; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_287;
  reg [1:0] btb_h_count_29; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_288;
  reg [1:0] btb_h_count_30; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_289;
  reg [1:0] btb_h_count_31; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_290;
  reg [1:0] btb_h_count_32; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_291;
  reg [1:0] btb_h_count_33; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_292;
  reg [1:0] btb_h_count_34; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_293;
  reg [1:0] btb_h_count_35; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_294;
  reg [1:0] btb_h_count_36; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_295;
  reg [1:0] btb_h_count_37; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_296;
  reg [1:0] btb_h_count_38; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_297;
  reg [1:0] btb_h_count_39; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_298;
  reg [1:0] btb_h_count_40; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_299;
  reg [1:0] btb_h_count_41; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_300;
  reg [1:0] btb_h_count_42; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_301;
  reg [1:0] btb_h_count_43; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_302;
  reg [1:0] btb_h_count_44; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_303;
  reg [1:0] btb_h_count_45; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_304;
  reg [1:0] btb_h_count_46; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_305;
  reg [1:0] btb_h_count_47; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_306;
  reg [1:0] btb_h_count_48; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_307;
  reg [1:0] btb_h_count_49; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_308;
  reg [1:0] btb_h_count_50; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_309;
  reg [1:0] btb_h_count_51; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_310;
  reg [1:0] btb_h_count_52; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_311;
  reg [1:0] btb_h_count_53; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_312;
  reg [1:0] btb_h_count_54; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_313;
  reg [1:0] btb_h_count_55; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_314;
  reg [1:0] btb_h_count_56; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_315;
  reg [1:0] btb_h_count_57; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_316;
  reg [1:0] btb_h_count_58; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_317;
  reg [1:0] btb_h_count_59; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_318;
  reg [1:0] btb_h_count_60; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_319;
  reg [1:0] btb_h_count_61; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_320;
  reg [1:0] btb_h_count_62; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_321;
  reg [1:0] btb_h_count_63; // @[BTB.scala 82:20:@1086.4]
  reg [31:0] _RAND_322;
  wire [28:0] _T_175; // @[BTB.scala 99:43:@1088.4]
  wire [29:0] _T_178; // @[Cat.scala 30:58:@1089.4]
  wire [31:0] predict_0_cont_tgt; // @[Cat.scala 30:58:@1090.4]
  wire [32:0] _T_181; // @[BTB.scala 100:46:@1092.4]
  wire [31:0] predict_1_cont_tgt; // @[BTB.scala 100:46:@1093.4]
  wire  _T_183; // @[BTB.scala 101:55:@1095.4]
  wire  _T_186; // @[BTB.scala 101:41:@1097.4]
  wire [29:0] if_pc_0; // @[Cat.scala 30:58:@1102.4]
  wire  _T_198; // @[BTB.scala 105:47:@1104.4]
  wire  _T_199; // @[BTB.scala 105:47:@1105.4]
  wire  _T_200; // @[BTB.scala 105:47:@1106.4]
  wire  _T_201; // @[BTB.scala 105:47:@1107.4]
  wire  _T_202; // @[BTB.scala 105:47:@1108.4]
  wire  _T_203; // @[BTB.scala 105:47:@1109.4]
  wire  _T_204; // @[BTB.scala 105:47:@1110.4]
  wire  _T_205; // @[BTB.scala 105:47:@1111.4]
  wire  _T_206; // @[BTB.scala 105:47:@1112.4]
  wire  _T_207; // @[BTB.scala 105:47:@1113.4]
  wire  _T_208; // @[BTB.scala 105:47:@1114.4]
  wire  _T_209; // @[BTB.scala 105:47:@1115.4]
  wire  _T_210; // @[BTB.scala 105:47:@1116.4]
  wire  _T_211; // @[BTB.scala 105:47:@1117.4]
  wire  _T_212; // @[BTB.scala 105:47:@1118.4]
  wire  _T_213; // @[BTB.scala 105:47:@1119.4]
  wire  _T_214; // @[BTB.scala 105:47:@1120.4]
  wire  _T_215; // @[BTB.scala 105:47:@1121.4]
  wire  _T_216; // @[BTB.scala 105:47:@1122.4]
  wire  _T_217; // @[BTB.scala 105:47:@1123.4]
  wire  _T_218; // @[BTB.scala 105:47:@1124.4]
  wire  _T_219; // @[BTB.scala 105:47:@1125.4]
  wire  _T_220; // @[BTB.scala 105:47:@1126.4]
  wire  _T_221; // @[BTB.scala 105:47:@1127.4]
  wire  _T_222; // @[BTB.scala 105:47:@1128.4]
  wire  _T_223; // @[BTB.scala 105:47:@1129.4]
  wire  _T_224; // @[BTB.scala 105:47:@1130.4]
  wire  _T_225; // @[BTB.scala 105:47:@1131.4]
  wire  _T_226; // @[BTB.scala 105:47:@1132.4]
  wire  _T_227; // @[BTB.scala 105:47:@1133.4]
  wire  _T_228; // @[BTB.scala 105:47:@1134.4]
  wire  _T_229; // @[BTB.scala 105:47:@1135.4]
  wire  _T_230; // @[BTB.scala 105:47:@1136.4]
  wire  _T_231; // @[BTB.scala 105:47:@1137.4]
  wire  _T_232; // @[BTB.scala 105:47:@1138.4]
  wire  _T_233; // @[BTB.scala 105:47:@1139.4]
  wire  _T_234; // @[BTB.scala 105:47:@1140.4]
  wire  _T_235; // @[BTB.scala 105:47:@1141.4]
  wire  _T_236; // @[BTB.scala 105:47:@1142.4]
  wire  _T_237; // @[BTB.scala 105:47:@1143.4]
  wire  _T_238; // @[BTB.scala 105:47:@1144.4]
  wire  _T_239; // @[BTB.scala 105:47:@1145.4]
  wire  _T_240; // @[BTB.scala 105:47:@1146.4]
  wire  _T_241; // @[BTB.scala 105:47:@1147.4]
  wire  _T_242; // @[BTB.scala 105:47:@1148.4]
  wire  _T_243; // @[BTB.scala 105:47:@1149.4]
  wire  _T_244; // @[BTB.scala 105:47:@1150.4]
  wire  _T_245; // @[BTB.scala 105:47:@1151.4]
  wire  _T_246; // @[BTB.scala 105:47:@1152.4]
  wire  _T_247; // @[BTB.scala 105:47:@1153.4]
  wire  _T_248; // @[BTB.scala 105:47:@1154.4]
  wire  _T_249; // @[BTB.scala 105:47:@1155.4]
  wire  _T_250; // @[BTB.scala 105:47:@1156.4]
  wire  _T_251; // @[BTB.scala 105:47:@1157.4]
  wire  _T_252; // @[BTB.scala 105:47:@1158.4]
  wire  _T_253; // @[BTB.scala 105:47:@1159.4]
  wire  _T_254; // @[BTB.scala 105:47:@1160.4]
  wire  _T_255; // @[BTB.scala 105:47:@1161.4]
  wire  _T_256; // @[BTB.scala 105:47:@1162.4]
  wire  _T_257; // @[BTB.scala 105:47:@1163.4]
  wire  _T_258; // @[BTB.scala 105:47:@1164.4]
  wire  _T_259; // @[BTB.scala 105:47:@1165.4]
  wire  _T_260; // @[BTB.scala 105:47:@1166.4]
  wire  _T_261; // @[BTB.scala 105:47:@1167.4]
  wire [7:0] _T_338; // @[BTB.scala 105:62:@1239.4]
  wire [15:0] _T_346; // @[BTB.scala 105:62:@1247.4]
  wire [7:0] _T_353; // @[BTB.scala 105:62:@1254.4]
  wire [31:0] _T_362; // @[BTB.scala 105:62:@1263.4]
  wire [7:0] _T_369; // @[BTB.scala 105:62:@1270.4]
  wire [15:0] _T_377; // @[BTB.scala 105:62:@1278.4]
  wire [7:0] _T_384; // @[BTB.scala 105:62:@1285.4]
  wire [31:0] _T_393; // @[BTB.scala 105:62:@1294.4]
  wire [63:0] _T_394; // @[BTB.scala 105:62:@1295.4]
  wire [7:0] _T_401; // @[BTB.scala 105:81:@1302.4]
  wire [15:0] _T_409; // @[BTB.scala 105:81:@1310.4]
  wire [7:0] _T_416; // @[BTB.scala 105:81:@1317.4]
  wire [31:0] _T_425; // @[BTB.scala 105:81:@1326.4]
  wire [7:0] _T_432; // @[BTB.scala 105:81:@1333.4]
  wire [15:0] _T_440; // @[BTB.scala 105:81:@1341.4]
  wire [7:0] _T_447; // @[BTB.scala 105:81:@1348.4]
  wire [31:0] _T_456; // @[BTB.scala 105:81:@1357.4]
  wire [63:0] _T_457; // @[BTB.scala 105:81:@1358.4]
  wire [63:0] predict_0_lookup; // @[BTB.scala 105:69:@1359.4]
  wire  _T_459; // @[Mux.scala 21:36:@1361.4]
  wire  _T_460; // @[Mux.scala 21:36:@1362.4]
  wire  _T_461; // @[Mux.scala 21:36:@1363.4]
  wire  _T_462; // @[Mux.scala 21:36:@1364.4]
  wire  _T_463; // @[Mux.scala 21:36:@1365.4]
  wire  _T_464; // @[Mux.scala 21:36:@1366.4]
  wire  _T_465; // @[Mux.scala 21:36:@1367.4]
  wire  _T_466; // @[Mux.scala 21:36:@1368.4]
  wire  _T_467; // @[Mux.scala 21:36:@1369.4]
  wire  _T_468; // @[Mux.scala 21:36:@1370.4]
  wire  _T_469; // @[Mux.scala 21:36:@1371.4]
  wire  _T_470; // @[Mux.scala 21:36:@1372.4]
  wire  _T_471; // @[Mux.scala 21:36:@1373.4]
  wire  _T_472; // @[Mux.scala 21:36:@1374.4]
  wire  _T_473; // @[Mux.scala 21:36:@1375.4]
  wire  _T_474; // @[Mux.scala 21:36:@1376.4]
  wire  _T_475; // @[Mux.scala 21:36:@1377.4]
  wire  _T_476; // @[Mux.scala 21:36:@1378.4]
  wire  _T_477; // @[Mux.scala 21:36:@1379.4]
  wire  _T_478; // @[Mux.scala 21:36:@1380.4]
  wire  _T_479; // @[Mux.scala 21:36:@1381.4]
  wire  _T_480; // @[Mux.scala 21:36:@1382.4]
  wire  _T_481; // @[Mux.scala 21:36:@1383.4]
  wire  _T_482; // @[Mux.scala 21:36:@1384.4]
  wire  _T_483; // @[Mux.scala 21:36:@1385.4]
  wire  _T_484; // @[Mux.scala 21:36:@1386.4]
  wire  _T_485; // @[Mux.scala 21:36:@1387.4]
  wire  _T_486; // @[Mux.scala 21:36:@1388.4]
  wire  _T_487; // @[Mux.scala 21:36:@1389.4]
  wire  _T_488; // @[Mux.scala 21:36:@1390.4]
  wire  _T_489; // @[Mux.scala 21:36:@1391.4]
  wire  _T_490; // @[Mux.scala 21:36:@1392.4]
  wire  _T_491; // @[Mux.scala 21:36:@1393.4]
  wire  _T_492; // @[Mux.scala 21:36:@1394.4]
  wire  _T_493; // @[Mux.scala 21:36:@1395.4]
  wire  _T_494; // @[Mux.scala 21:36:@1396.4]
  wire  _T_495; // @[Mux.scala 21:36:@1397.4]
  wire  _T_496; // @[Mux.scala 21:36:@1398.4]
  wire  _T_497; // @[Mux.scala 21:36:@1399.4]
  wire  _T_498; // @[Mux.scala 21:36:@1400.4]
  wire  _T_499; // @[Mux.scala 21:36:@1401.4]
  wire  _T_500; // @[Mux.scala 21:36:@1402.4]
  wire  _T_501; // @[Mux.scala 21:36:@1403.4]
  wire  _T_502; // @[Mux.scala 21:36:@1404.4]
  wire  _T_503; // @[Mux.scala 21:36:@1405.4]
  wire  _T_504; // @[Mux.scala 21:36:@1406.4]
  wire  _T_505; // @[Mux.scala 21:36:@1407.4]
  wire  _T_506; // @[Mux.scala 21:36:@1408.4]
  wire  _T_507; // @[Mux.scala 21:36:@1409.4]
  wire  _T_508; // @[Mux.scala 21:36:@1410.4]
  wire  _T_509; // @[Mux.scala 21:36:@1411.4]
  wire  _T_510; // @[Mux.scala 21:36:@1412.4]
  wire  _T_511; // @[Mux.scala 21:36:@1413.4]
  wire  _T_512; // @[Mux.scala 21:36:@1414.4]
  wire  _T_513; // @[Mux.scala 21:36:@1415.4]
  wire  _T_514; // @[Mux.scala 21:36:@1416.4]
  wire  _T_515; // @[Mux.scala 21:36:@1417.4]
  wire  _T_516; // @[Mux.scala 21:36:@1418.4]
  wire  _T_517; // @[Mux.scala 21:36:@1419.4]
  wire  _T_518; // @[Mux.scala 21:36:@1420.4]
  wire  _T_519; // @[Mux.scala 21:36:@1421.4]
  wire  _T_520; // @[Mux.scala 21:36:@1422.4]
  wire  _T_521; // @[Mux.scala 21:36:@1423.4]
  wire  _T_522; // @[Mux.scala 21:36:@1424.4]
  wire [29:0] _T_525; // @[Mux.scala 19:72:@1425.4]
  wire [29:0] _T_527; // @[Mux.scala 19:72:@1426.4]
  wire [29:0] _T_529; // @[Mux.scala 19:72:@1427.4]
  wire [29:0] _T_531; // @[Mux.scala 19:72:@1428.4]
  wire [29:0] _T_533; // @[Mux.scala 19:72:@1429.4]
  wire [29:0] _T_535; // @[Mux.scala 19:72:@1430.4]
  wire [29:0] _T_537; // @[Mux.scala 19:72:@1431.4]
  wire [29:0] _T_539; // @[Mux.scala 19:72:@1432.4]
  wire [29:0] _T_541; // @[Mux.scala 19:72:@1433.4]
  wire [29:0] _T_543; // @[Mux.scala 19:72:@1434.4]
  wire [29:0] _T_545; // @[Mux.scala 19:72:@1435.4]
  wire [29:0] _T_547; // @[Mux.scala 19:72:@1436.4]
  wire [29:0] _T_549; // @[Mux.scala 19:72:@1437.4]
  wire [29:0] _T_551; // @[Mux.scala 19:72:@1438.4]
  wire [29:0] _T_553; // @[Mux.scala 19:72:@1439.4]
  wire [29:0] _T_555; // @[Mux.scala 19:72:@1440.4]
  wire [29:0] _T_557; // @[Mux.scala 19:72:@1441.4]
  wire [29:0] _T_559; // @[Mux.scala 19:72:@1442.4]
  wire [29:0] _T_561; // @[Mux.scala 19:72:@1443.4]
  wire [29:0] _T_563; // @[Mux.scala 19:72:@1444.4]
  wire [29:0] _T_565; // @[Mux.scala 19:72:@1445.4]
  wire [29:0] _T_567; // @[Mux.scala 19:72:@1446.4]
  wire [29:0] _T_569; // @[Mux.scala 19:72:@1447.4]
  wire [29:0] _T_571; // @[Mux.scala 19:72:@1448.4]
  wire [29:0] _T_573; // @[Mux.scala 19:72:@1449.4]
  wire [29:0] _T_575; // @[Mux.scala 19:72:@1450.4]
  wire [29:0] _T_577; // @[Mux.scala 19:72:@1451.4]
  wire [29:0] _T_579; // @[Mux.scala 19:72:@1452.4]
  wire [29:0] _T_581; // @[Mux.scala 19:72:@1453.4]
  wire [29:0] _T_583; // @[Mux.scala 19:72:@1454.4]
  wire [29:0] _T_585; // @[Mux.scala 19:72:@1455.4]
  wire [29:0] _T_587; // @[Mux.scala 19:72:@1456.4]
  wire [29:0] _T_589; // @[Mux.scala 19:72:@1457.4]
  wire [29:0] _T_591; // @[Mux.scala 19:72:@1458.4]
  wire [29:0] _T_593; // @[Mux.scala 19:72:@1459.4]
  wire [29:0] _T_595; // @[Mux.scala 19:72:@1460.4]
  wire [29:0] _T_597; // @[Mux.scala 19:72:@1461.4]
  wire [29:0] _T_599; // @[Mux.scala 19:72:@1462.4]
  wire [29:0] _T_601; // @[Mux.scala 19:72:@1463.4]
  wire [29:0] _T_603; // @[Mux.scala 19:72:@1464.4]
  wire [29:0] _T_605; // @[Mux.scala 19:72:@1465.4]
  wire [29:0] _T_607; // @[Mux.scala 19:72:@1466.4]
  wire [29:0] _T_609; // @[Mux.scala 19:72:@1467.4]
  wire [29:0] _T_611; // @[Mux.scala 19:72:@1468.4]
  wire [29:0] _T_613; // @[Mux.scala 19:72:@1469.4]
  wire [29:0] _T_615; // @[Mux.scala 19:72:@1470.4]
  wire [29:0] _T_617; // @[Mux.scala 19:72:@1471.4]
  wire [29:0] _T_619; // @[Mux.scala 19:72:@1472.4]
  wire [29:0] _T_621; // @[Mux.scala 19:72:@1473.4]
  wire [29:0] _T_623; // @[Mux.scala 19:72:@1474.4]
  wire [29:0] _T_625; // @[Mux.scala 19:72:@1475.4]
  wire [29:0] _T_627; // @[Mux.scala 19:72:@1476.4]
  wire [29:0] _T_629; // @[Mux.scala 19:72:@1477.4]
  wire [29:0] _T_631; // @[Mux.scala 19:72:@1478.4]
  wire [29:0] _T_633; // @[Mux.scala 19:72:@1479.4]
  wire [29:0] _T_635; // @[Mux.scala 19:72:@1480.4]
  wire [29:0] _T_637; // @[Mux.scala 19:72:@1481.4]
  wire [29:0] _T_639; // @[Mux.scala 19:72:@1482.4]
  wire [29:0] _T_641; // @[Mux.scala 19:72:@1483.4]
  wire [29:0] _T_643; // @[Mux.scala 19:72:@1484.4]
  wire [29:0] _T_645; // @[Mux.scala 19:72:@1485.4]
  wire [29:0] _T_647; // @[Mux.scala 19:72:@1486.4]
  wire [29:0] _T_649; // @[Mux.scala 19:72:@1487.4]
  wire [29:0] _T_651; // @[Mux.scala 19:72:@1488.4]
  wire [29:0] _T_652; // @[Mux.scala 19:72:@1489.4]
  wire [29:0] _T_653; // @[Mux.scala 19:72:@1490.4]
  wire [29:0] _T_654; // @[Mux.scala 19:72:@1491.4]
  wire [29:0] _T_655; // @[Mux.scala 19:72:@1492.4]
  wire [29:0] _T_656; // @[Mux.scala 19:72:@1493.4]
  wire [29:0] _T_657; // @[Mux.scala 19:72:@1494.4]
  wire [29:0] _T_658; // @[Mux.scala 19:72:@1495.4]
  wire [29:0] _T_659; // @[Mux.scala 19:72:@1496.4]
  wire [29:0] _T_660; // @[Mux.scala 19:72:@1497.4]
  wire [29:0] _T_661; // @[Mux.scala 19:72:@1498.4]
  wire [29:0] _T_662; // @[Mux.scala 19:72:@1499.4]
  wire [29:0] _T_663; // @[Mux.scala 19:72:@1500.4]
  wire [29:0] _T_664; // @[Mux.scala 19:72:@1501.4]
  wire [29:0] _T_665; // @[Mux.scala 19:72:@1502.4]
  wire [29:0] _T_666; // @[Mux.scala 19:72:@1503.4]
  wire [29:0] _T_667; // @[Mux.scala 19:72:@1504.4]
  wire [29:0] _T_668; // @[Mux.scala 19:72:@1505.4]
  wire [29:0] _T_669; // @[Mux.scala 19:72:@1506.4]
  wire [29:0] _T_670; // @[Mux.scala 19:72:@1507.4]
  wire [29:0] _T_671; // @[Mux.scala 19:72:@1508.4]
  wire [29:0] _T_672; // @[Mux.scala 19:72:@1509.4]
  wire [29:0] _T_673; // @[Mux.scala 19:72:@1510.4]
  wire [29:0] _T_674; // @[Mux.scala 19:72:@1511.4]
  wire [29:0] _T_675; // @[Mux.scala 19:72:@1512.4]
  wire [29:0] _T_676; // @[Mux.scala 19:72:@1513.4]
  wire [29:0] _T_677; // @[Mux.scala 19:72:@1514.4]
  wire [29:0] _T_678; // @[Mux.scala 19:72:@1515.4]
  wire [29:0] _T_679; // @[Mux.scala 19:72:@1516.4]
  wire [29:0] _T_680; // @[Mux.scala 19:72:@1517.4]
  wire [29:0] _T_681; // @[Mux.scala 19:72:@1518.4]
  wire [29:0] _T_682; // @[Mux.scala 19:72:@1519.4]
  wire [29:0] _T_683; // @[Mux.scala 19:72:@1520.4]
  wire [29:0] _T_684; // @[Mux.scala 19:72:@1521.4]
  wire [29:0] _T_685; // @[Mux.scala 19:72:@1522.4]
  wire [29:0] _T_686; // @[Mux.scala 19:72:@1523.4]
  wire [29:0] _T_687; // @[Mux.scala 19:72:@1524.4]
  wire [29:0] _T_688; // @[Mux.scala 19:72:@1525.4]
  wire [29:0] _T_689; // @[Mux.scala 19:72:@1526.4]
  wire [29:0] _T_690; // @[Mux.scala 19:72:@1527.4]
  wire [29:0] _T_691; // @[Mux.scala 19:72:@1528.4]
  wire [29:0] _T_692; // @[Mux.scala 19:72:@1529.4]
  wire [29:0] _T_693; // @[Mux.scala 19:72:@1530.4]
  wire [29:0] _T_694; // @[Mux.scala 19:72:@1531.4]
  wire [29:0] _T_695; // @[Mux.scala 19:72:@1532.4]
  wire [29:0] _T_696; // @[Mux.scala 19:72:@1533.4]
  wire [29:0] _T_697; // @[Mux.scala 19:72:@1534.4]
  wire [29:0] _T_698; // @[Mux.scala 19:72:@1535.4]
  wire [29:0] _T_699; // @[Mux.scala 19:72:@1536.4]
  wire [29:0] _T_700; // @[Mux.scala 19:72:@1537.4]
  wire [29:0] _T_701; // @[Mux.scala 19:72:@1538.4]
  wire [29:0] _T_702; // @[Mux.scala 19:72:@1539.4]
  wire [29:0] _T_703; // @[Mux.scala 19:72:@1540.4]
  wire [29:0] _T_704; // @[Mux.scala 19:72:@1541.4]
  wire [29:0] _T_705; // @[Mux.scala 19:72:@1542.4]
  wire [29:0] _T_706; // @[Mux.scala 19:72:@1543.4]
  wire [29:0] _T_707; // @[Mux.scala 19:72:@1544.4]
  wire [29:0] _T_708; // @[Mux.scala 19:72:@1545.4]
  wire [29:0] _T_709; // @[Mux.scala 19:72:@1546.4]
  wire [29:0] _T_710; // @[Mux.scala 19:72:@1547.4]
  wire [29:0] _T_711; // @[Mux.scala 19:72:@1548.4]
  wire [29:0] _T_712; // @[Mux.scala 19:72:@1549.4]
  wire [29:0] _T_713; // @[Mux.scala 19:72:@1550.4]
  wire [29:0] _T_714; // @[Mux.scala 19:72:@1551.4]
  wire [31:0] predict_0_jump_tgt; // @[Cat.scala 30:58:@1554.4]
  wire [1:0] _T_785; // @[Mux.scala 19:72:@1620.4]
  wire [1:0] _T_787; // @[Mux.scala 19:72:@1621.4]
  wire [1:0] _T_789; // @[Mux.scala 19:72:@1622.4]
  wire [1:0] _T_791; // @[Mux.scala 19:72:@1623.4]
  wire [1:0] _T_793; // @[Mux.scala 19:72:@1624.4]
  wire [1:0] _T_795; // @[Mux.scala 19:72:@1625.4]
  wire [1:0] _T_797; // @[Mux.scala 19:72:@1626.4]
  wire [1:0] _T_799; // @[Mux.scala 19:72:@1627.4]
  wire [1:0] _T_801; // @[Mux.scala 19:72:@1628.4]
  wire [1:0] _T_803; // @[Mux.scala 19:72:@1629.4]
  wire [1:0] _T_805; // @[Mux.scala 19:72:@1630.4]
  wire [1:0] _T_807; // @[Mux.scala 19:72:@1631.4]
  wire [1:0] _T_809; // @[Mux.scala 19:72:@1632.4]
  wire [1:0] _T_811; // @[Mux.scala 19:72:@1633.4]
  wire [1:0] _T_813; // @[Mux.scala 19:72:@1634.4]
  wire [1:0] _T_815; // @[Mux.scala 19:72:@1635.4]
  wire [1:0] _T_817; // @[Mux.scala 19:72:@1636.4]
  wire [1:0] _T_819; // @[Mux.scala 19:72:@1637.4]
  wire [1:0] _T_821; // @[Mux.scala 19:72:@1638.4]
  wire [1:0] _T_823; // @[Mux.scala 19:72:@1639.4]
  wire [1:0] _T_825; // @[Mux.scala 19:72:@1640.4]
  wire [1:0] _T_827; // @[Mux.scala 19:72:@1641.4]
  wire [1:0] _T_829; // @[Mux.scala 19:72:@1642.4]
  wire [1:0] _T_831; // @[Mux.scala 19:72:@1643.4]
  wire [1:0] _T_833; // @[Mux.scala 19:72:@1644.4]
  wire [1:0] _T_835; // @[Mux.scala 19:72:@1645.4]
  wire [1:0] _T_837; // @[Mux.scala 19:72:@1646.4]
  wire [1:0] _T_839; // @[Mux.scala 19:72:@1647.4]
  wire [1:0] _T_841; // @[Mux.scala 19:72:@1648.4]
  wire [1:0] _T_843; // @[Mux.scala 19:72:@1649.4]
  wire [1:0] _T_845; // @[Mux.scala 19:72:@1650.4]
  wire [1:0] _T_847; // @[Mux.scala 19:72:@1651.4]
  wire [1:0] _T_849; // @[Mux.scala 19:72:@1652.4]
  wire [1:0] _T_851; // @[Mux.scala 19:72:@1653.4]
  wire [1:0] _T_853; // @[Mux.scala 19:72:@1654.4]
  wire [1:0] _T_855; // @[Mux.scala 19:72:@1655.4]
  wire [1:0] _T_857; // @[Mux.scala 19:72:@1656.4]
  wire [1:0] _T_859; // @[Mux.scala 19:72:@1657.4]
  wire [1:0] _T_861; // @[Mux.scala 19:72:@1658.4]
  wire [1:0] _T_863; // @[Mux.scala 19:72:@1659.4]
  wire [1:0] _T_865; // @[Mux.scala 19:72:@1660.4]
  wire [1:0] _T_867; // @[Mux.scala 19:72:@1661.4]
  wire [1:0] _T_869; // @[Mux.scala 19:72:@1662.4]
  wire [1:0] _T_871; // @[Mux.scala 19:72:@1663.4]
  wire [1:0] _T_873; // @[Mux.scala 19:72:@1664.4]
  wire [1:0] _T_875; // @[Mux.scala 19:72:@1665.4]
  wire [1:0] _T_877; // @[Mux.scala 19:72:@1666.4]
  wire [1:0] _T_879; // @[Mux.scala 19:72:@1667.4]
  wire [1:0] _T_881; // @[Mux.scala 19:72:@1668.4]
  wire [1:0] _T_883; // @[Mux.scala 19:72:@1669.4]
  wire [1:0] _T_885; // @[Mux.scala 19:72:@1670.4]
  wire [1:0] _T_887; // @[Mux.scala 19:72:@1671.4]
  wire [1:0] _T_889; // @[Mux.scala 19:72:@1672.4]
  wire [1:0] _T_891; // @[Mux.scala 19:72:@1673.4]
  wire [1:0] _T_893; // @[Mux.scala 19:72:@1674.4]
  wire [1:0] _T_895; // @[Mux.scala 19:72:@1675.4]
  wire [1:0] _T_897; // @[Mux.scala 19:72:@1676.4]
  wire [1:0] _T_899; // @[Mux.scala 19:72:@1677.4]
  wire [1:0] _T_901; // @[Mux.scala 19:72:@1678.4]
  wire [1:0] _T_903; // @[Mux.scala 19:72:@1679.4]
  wire [1:0] _T_905; // @[Mux.scala 19:72:@1680.4]
  wire [1:0] _T_907; // @[Mux.scala 19:72:@1681.4]
  wire [1:0] _T_909; // @[Mux.scala 19:72:@1682.4]
  wire [1:0] _T_911; // @[Mux.scala 19:72:@1683.4]
  wire [1:0] _T_912; // @[Mux.scala 19:72:@1684.4]
  wire [1:0] _T_913; // @[Mux.scala 19:72:@1685.4]
  wire [1:0] _T_914; // @[Mux.scala 19:72:@1686.4]
  wire [1:0] _T_915; // @[Mux.scala 19:72:@1687.4]
  wire [1:0] _T_916; // @[Mux.scala 19:72:@1688.4]
  wire [1:0] _T_917; // @[Mux.scala 19:72:@1689.4]
  wire [1:0] _T_918; // @[Mux.scala 19:72:@1690.4]
  wire [1:0] _T_919; // @[Mux.scala 19:72:@1691.4]
  wire [1:0] _T_920; // @[Mux.scala 19:72:@1692.4]
  wire [1:0] _T_921; // @[Mux.scala 19:72:@1693.4]
  wire [1:0] _T_922; // @[Mux.scala 19:72:@1694.4]
  wire [1:0] _T_923; // @[Mux.scala 19:72:@1695.4]
  wire [1:0] _T_924; // @[Mux.scala 19:72:@1696.4]
  wire [1:0] _T_925; // @[Mux.scala 19:72:@1697.4]
  wire [1:0] _T_926; // @[Mux.scala 19:72:@1698.4]
  wire [1:0] _T_927; // @[Mux.scala 19:72:@1699.4]
  wire [1:0] _T_928; // @[Mux.scala 19:72:@1700.4]
  wire [1:0] _T_929; // @[Mux.scala 19:72:@1701.4]
  wire [1:0] _T_930; // @[Mux.scala 19:72:@1702.4]
  wire [1:0] _T_931; // @[Mux.scala 19:72:@1703.4]
  wire [1:0] _T_932; // @[Mux.scala 19:72:@1704.4]
  wire [1:0] _T_933; // @[Mux.scala 19:72:@1705.4]
  wire [1:0] _T_934; // @[Mux.scala 19:72:@1706.4]
  wire [1:0] _T_935; // @[Mux.scala 19:72:@1707.4]
  wire [1:0] _T_936; // @[Mux.scala 19:72:@1708.4]
  wire [1:0] _T_937; // @[Mux.scala 19:72:@1709.4]
  wire [1:0] _T_938; // @[Mux.scala 19:72:@1710.4]
  wire [1:0] _T_939; // @[Mux.scala 19:72:@1711.4]
  wire [1:0] _T_940; // @[Mux.scala 19:72:@1712.4]
  wire [1:0] _T_941; // @[Mux.scala 19:72:@1713.4]
  wire [1:0] _T_942; // @[Mux.scala 19:72:@1714.4]
  wire [1:0] _T_943; // @[Mux.scala 19:72:@1715.4]
  wire [1:0] _T_944; // @[Mux.scala 19:72:@1716.4]
  wire [1:0] _T_945; // @[Mux.scala 19:72:@1717.4]
  wire [1:0] _T_946; // @[Mux.scala 19:72:@1718.4]
  wire [1:0] _T_947; // @[Mux.scala 19:72:@1719.4]
  wire [1:0] _T_948; // @[Mux.scala 19:72:@1720.4]
  wire [1:0] _T_949; // @[Mux.scala 19:72:@1721.4]
  wire [1:0] _T_950; // @[Mux.scala 19:72:@1722.4]
  wire [1:0] _T_951; // @[Mux.scala 19:72:@1723.4]
  wire [1:0] _T_952; // @[Mux.scala 19:72:@1724.4]
  wire [1:0] _T_953; // @[Mux.scala 19:72:@1725.4]
  wire [1:0] _T_954; // @[Mux.scala 19:72:@1726.4]
  wire [1:0] _T_955; // @[Mux.scala 19:72:@1727.4]
  wire [1:0] _T_956; // @[Mux.scala 19:72:@1728.4]
  wire [1:0] _T_957; // @[Mux.scala 19:72:@1729.4]
  wire [1:0] _T_958; // @[Mux.scala 19:72:@1730.4]
  wire [1:0] _T_959; // @[Mux.scala 19:72:@1731.4]
  wire [1:0] _T_960; // @[Mux.scala 19:72:@1732.4]
  wire [1:0] _T_961; // @[Mux.scala 19:72:@1733.4]
  wire [1:0] _T_962; // @[Mux.scala 19:72:@1734.4]
  wire [1:0] _T_963; // @[Mux.scala 19:72:@1735.4]
  wire [1:0] _T_964; // @[Mux.scala 19:72:@1736.4]
  wire [1:0] _T_965; // @[Mux.scala 19:72:@1737.4]
  wire [1:0] _T_966; // @[Mux.scala 19:72:@1738.4]
  wire [1:0] _T_967; // @[Mux.scala 19:72:@1739.4]
  wire [1:0] _T_968; // @[Mux.scala 19:72:@1740.4]
  wire [1:0] _T_969; // @[Mux.scala 19:72:@1741.4]
  wire [1:0] _T_970; // @[Mux.scala 19:72:@1742.4]
  wire [1:0] _T_971; // @[Mux.scala 19:72:@1743.4]
  wire [1:0] _T_972; // @[Mux.scala 19:72:@1744.4]
  wire [1:0] _T_973; // @[Mux.scala 19:72:@1745.4]
  wire [1:0] predict_0_bj_type; // @[Mux.scala 19:72:@1746.4]
  wire [1:0] _T_1043; // @[Mux.scala 19:72:@1814.4]
  wire [1:0] _T_1045; // @[Mux.scala 19:72:@1815.4]
  wire [1:0] _T_1047; // @[Mux.scala 19:72:@1816.4]
  wire [1:0] _T_1049; // @[Mux.scala 19:72:@1817.4]
  wire [1:0] _T_1051; // @[Mux.scala 19:72:@1818.4]
  wire [1:0] _T_1053; // @[Mux.scala 19:72:@1819.4]
  wire [1:0] _T_1055; // @[Mux.scala 19:72:@1820.4]
  wire [1:0] _T_1057; // @[Mux.scala 19:72:@1821.4]
  wire [1:0] _T_1059; // @[Mux.scala 19:72:@1822.4]
  wire [1:0] _T_1061; // @[Mux.scala 19:72:@1823.4]
  wire [1:0] _T_1063; // @[Mux.scala 19:72:@1824.4]
  wire [1:0] _T_1065; // @[Mux.scala 19:72:@1825.4]
  wire [1:0] _T_1067; // @[Mux.scala 19:72:@1826.4]
  wire [1:0] _T_1069; // @[Mux.scala 19:72:@1827.4]
  wire [1:0] _T_1071; // @[Mux.scala 19:72:@1828.4]
  wire [1:0] _T_1073; // @[Mux.scala 19:72:@1829.4]
  wire [1:0] _T_1075; // @[Mux.scala 19:72:@1830.4]
  wire [1:0] _T_1077; // @[Mux.scala 19:72:@1831.4]
  wire [1:0] _T_1079; // @[Mux.scala 19:72:@1832.4]
  wire [1:0] _T_1081; // @[Mux.scala 19:72:@1833.4]
  wire [1:0] _T_1083; // @[Mux.scala 19:72:@1834.4]
  wire [1:0] _T_1085; // @[Mux.scala 19:72:@1835.4]
  wire [1:0] _T_1087; // @[Mux.scala 19:72:@1836.4]
  wire [1:0] _T_1089; // @[Mux.scala 19:72:@1837.4]
  wire [1:0] _T_1091; // @[Mux.scala 19:72:@1838.4]
  wire [1:0] _T_1093; // @[Mux.scala 19:72:@1839.4]
  wire [1:0] _T_1095; // @[Mux.scala 19:72:@1840.4]
  wire [1:0] _T_1097; // @[Mux.scala 19:72:@1841.4]
  wire [1:0] _T_1099; // @[Mux.scala 19:72:@1842.4]
  wire [1:0] _T_1101; // @[Mux.scala 19:72:@1843.4]
  wire [1:0] _T_1103; // @[Mux.scala 19:72:@1844.4]
  wire [1:0] _T_1105; // @[Mux.scala 19:72:@1845.4]
  wire [1:0] _T_1107; // @[Mux.scala 19:72:@1846.4]
  wire [1:0] _T_1109; // @[Mux.scala 19:72:@1847.4]
  wire [1:0] _T_1111; // @[Mux.scala 19:72:@1848.4]
  wire [1:0] _T_1113; // @[Mux.scala 19:72:@1849.4]
  wire [1:0] _T_1115; // @[Mux.scala 19:72:@1850.4]
  wire [1:0] _T_1117; // @[Mux.scala 19:72:@1851.4]
  wire [1:0] _T_1119; // @[Mux.scala 19:72:@1852.4]
  wire [1:0] _T_1121; // @[Mux.scala 19:72:@1853.4]
  wire [1:0] _T_1123; // @[Mux.scala 19:72:@1854.4]
  wire [1:0] _T_1125; // @[Mux.scala 19:72:@1855.4]
  wire [1:0] _T_1127; // @[Mux.scala 19:72:@1856.4]
  wire [1:0] _T_1129; // @[Mux.scala 19:72:@1857.4]
  wire [1:0] _T_1131; // @[Mux.scala 19:72:@1858.4]
  wire [1:0] _T_1133; // @[Mux.scala 19:72:@1859.4]
  wire [1:0] _T_1135; // @[Mux.scala 19:72:@1860.4]
  wire [1:0] _T_1137; // @[Mux.scala 19:72:@1861.4]
  wire [1:0] _T_1139; // @[Mux.scala 19:72:@1862.4]
  wire [1:0] _T_1141; // @[Mux.scala 19:72:@1863.4]
  wire [1:0] _T_1143; // @[Mux.scala 19:72:@1864.4]
  wire [1:0] _T_1145; // @[Mux.scala 19:72:@1865.4]
  wire [1:0] _T_1147; // @[Mux.scala 19:72:@1866.4]
  wire [1:0] _T_1149; // @[Mux.scala 19:72:@1867.4]
  wire [1:0] _T_1151; // @[Mux.scala 19:72:@1868.4]
  wire [1:0] _T_1153; // @[Mux.scala 19:72:@1869.4]
  wire [1:0] _T_1155; // @[Mux.scala 19:72:@1870.4]
  wire [1:0] _T_1157; // @[Mux.scala 19:72:@1871.4]
  wire [1:0] _T_1159; // @[Mux.scala 19:72:@1872.4]
  wire [1:0] _T_1161; // @[Mux.scala 19:72:@1873.4]
  wire [1:0] _T_1163; // @[Mux.scala 19:72:@1874.4]
  wire [1:0] _T_1165; // @[Mux.scala 19:72:@1875.4]
  wire [1:0] _T_1167; // @[Mux.scala 19:72:@1876.4]
  wire [1:0] _T_1169; // @[Mux.scala 19:72:@1877.4]
  wire [1:0] _T_1170; // @[Mux.scala 19:72:@1878.4]
  wire [1:0] _T_1171; // @[Mux.scala 19:72:@1879.4]
  wire [1:0] _T_1172; // @[Mux.scala 19:72:@1880.4]
  wire [1:0] _T_1173; // @[Mux.scala 19:72:@1881.4]
  wire [1:0] _T_1174; // @[Mux.scala 19:72:@1882.4]
  wire [1:0] _T_1175; // @[Mux.scala 19:72:@1883.4]
  wire [1:0] _T_1176; // @[Mux.scala 19:72:@1884.4]
  wire [1:0] _T_1177; // @[Mux.scala 19:72:@1885.4]
  wire [1:0] _T_1178; // @[Mux.scala 19:72:@1886.4]
  wire [1:0] _T_1179; // @[Mux.scala 19:72:@1887.4]
  wire [1:0] _T_1180; // @[Mux.scala 19:72:@1888.4]
  wire [1:0] _T_1181; // @[Mux.scala 19:72:@1889.4]
  wire [1:0] _T_1182; // @[Mux.scala 19:72:@1890.4]
  wire [1:0] _T_1183; // @[Mux.scala 19:72:@1891.4]
  wire [1:0] _T_1184; // @[Mux.scala 19:72:@1892.4]
  wire [1:0] _T_1185; // @[Mux.scala 19:72:@1893.4]
  wire [1:0] _T_1186; // @[Mux.scala 19:72:@1894.4]
  wire [1:0] _T_1187; // @[Mux.scala 19:72:@1895.4]
  wire [1:0] _T_1188; // @[Mux.scala 19:72:@1896.4]
  wire [1:0] _T_1189; // @[Mux.scala 19:72:@1897.4]
  wire [1:0] _T_1190; // @[Mux.scala 19:72:@1898.4]
  wire [1:0] _T_1191; // @[Mux.scala 19:72:@1899.4]
  wire [1:0] _T_1192; // @[Mux.scala 19:72:@1900.4]
  wire [1:0] _T_1193; // @[Mux.scala 19:72:@1901.4]
  wire [1:0] _T_1194; // @[Mux.scala 19:72:@1902.4]
  wire [1:0] _T_1195; // @[Mux.scala 19:72:@1903.4]
  wire [1:0] _T_1196; // @[Mux.scala 19:72:@1904.4]
  wire [1:0] _T_1197; // @[Mux.scala 19:72:@1905.4]
  wire [1:0] _T_1198; // @[Mux.scala 19:72:@1906.4]
  wire [1:0] _T_1199; // @[Mux.scala 19:72:@1907.4]
  wire [1:0] _T_1200; // @[Mux.scala 19:72:@1908.4]
  wire [1:0] _T_1201; // @[Mux.scala 19:72:@1909.4]
  wire [1:0] _T_1202; // @[Mux.scala 19:72:@1910.4]
  wire [1:0] _T_1203; // @[Mux.scala 19:72:@1911.4]
  wire [1:0] _T_1204; // @[Mux.scala 19:72:@1912.4]
  wire [1:0] _T_1205; // @[Mux.scala 19:72:@1913.4]
  wire [1:0] _T_1206; // @[Mux.scala 19:72:@1914.4]
  wire [1:0] _T_1207; // @[Mux.scala 19:72:@1915.4]
  wire [1:0] _T_1208; // @[Mux.scala 19:72:@1916.4]
  wire [1:0] _T_1209; // @[Mux.scala 19:72:@1917.4]
  wire [1:0] _T_1210; // @[Mux.scala 19:72:@1918.4]
  wire [1:0] _T_1211; // @[Mux.scala 19:72:@1919.4]
  wire [1:0] _T_1212; // @[Mux.scala 19:72:@1920.4]
  wire [1:0] _T_1213; // @[Mux.scala 19:72:@1921.4]
  wire [1:0] _T_1214; // @[Mux.scala 19:72:@1922.4]
  wire [1:0] _T_1215; // @[Mux.scala 19:72:@1923.4]
  wire [1:0] _T_1216; // @[Mux.scala 19:72:@1924.4]
  wire [1:0] _T_1217; // @[Mux.scala 19:72:@1925.4]
  wire [1:0] _T_1218; // @[Mux.scala 19:72:@1926.4]
  wire [1:0] _T_1219; // @[Mux.scala 19:72:@1927.4]
  wire [1:0] _T_1220; // @[Mux.scala 19:72:@1928.4]
  wire [1:0] _T_1221; // @[Mux.scala 19:72:@1929.4]
  wire [1:0] _T_1222; // @[Mux.scala 19:72:@1930.4]
  wire [1:0] _T_1223; // @[Mux.scala 19:72:@1931.4]
  wire [1:0] _T_1224; // @[Mux.scala 19:72:@1932.4]
  wire [1:0] _T_1225; // @[Mux.scala 19:72:@1933.4]
  wire [1:0] _T_1226; // @[Mux.scala 19:72:@1934.4]
  wire [1:0] _T_1227; // @[Mux.scala 19:72:@1935.4]
  wire [1:0] _T_1228; // @[Mux.scala 19:72:@1936.4]
  wire [1:0] _T_1229; // @[Mux.scala 19:72:@1937.4]
  wire [1:0] _T_1230; // @[Mux.scala 19:72:@1938.4]
  wire [1:0] _T_1231; // @[Mux.scala 19:72:@1939.4]
  wire [1:0] predict_0_h_count; // @[Mux.scala 19:72:@1940.4]
  wire [9:0] _T_1236; // @[BTB.scala 110:54:@1945.4]
  wire [9:0] predict_0_gshxor; // @[BTB.scala 110:44:@1946.4]
  wire [8:0] _T_1240; // @[BTB.scala 113:42:@1952.4]
  wire [1:0] predict_0_gshare; // @[BTB.scala 98:21:@1087.4 BTB.scala 112:25:@1951.4]
  wire  _T_1241; // @[BTB.scala 47:40:@1953.4]
  wire  _T_1242; // @[BTB.scala 47:52:@1954.4]
  wire  predict_0_select; // @[BTB.scala 98:21:@1087.4 BTB.scala 111:25:@1949.4]
  wire  _T_1243; // @[BTB.scala 47:25:@1955.4]
  wire [9:0] predict_0_history; // @[Cat.scala 30:58:@1956.4]
  wire  _T_1246; // @[BTB.scala 40:28:@1958.4]
  wire  _T_1250; // @[BTB.scala 49:42:@1961.4]
  wire  _T_1254; // @[BTB.scala 49:63:@1965.4]
  wire  _T_1255; // @[BTB.scala 49:30:@1966.4]
  wire  _T_1260; // @[BTB.scala 119:54:@1973.4]
  wire [31:0] _T_1270; // @[BTB.scala 120:34:@1981.4]
  wire  _T_1275; // @[BTB.scala 105:47:@1987.4]
  wire  _T_1276; // @[BTB.scala 105:47:@1988.4]
  wire  _T_1277; // @[BTB.scala 105:47:@1989.4]
  wire  _T_1278; // @[BTB.scala 105:47:@1990.4]
  wire  _T_1279; // @[BTB.scala 105:47:@1991.4]
  wire  _T_1280; // @[BTB.scala 105:47:@1992.4]
  wire  _T_1281; // @[BTB.scala 105:47:@1993.4]
  wire  _T_1282; // @[BTB.scala 105:47:@1994.4]
  wire  _T_1283; // @[BTB.scala 105:47:@1995.4]
  wire  _T_1284; // @[BTB.scala 105:47:@1996.4]
  wire  _T_1285; // @[BTB.scala 105:47:@1997.4]
  wire  _T_1286; // @[BTB.scala 105:47:@1998.4]
  wire  _T_1287; // @[BTB.scala 105:47:@1999.4]
  wire  _T_1288; // @[BTB.scala 105:47:@2000.4]
  wire  _T_1289; // @[BTB.scala 105:47:@2001.4]
  wire  _T_1290; // @[BTB.scala 105:47:@2002.4]
  wire  _T_1291; // @[BTB.scala 105:47:@2003.4]
  wire  _T_1292; // @[BTB.scala 105:47:@2004.4]
  wire  _T_1293; // @[BTB.scala 105:47:@2005.4]
  wire  _T_1294; // @[BTB.scala 105:47:@2006.4]
  wire  _T_1295; // @[BTB.scala 105:47:@2007.4]
  wire  _T_1296; // @[BTB.scala 105:47:@2008.4]
  wire  _T_1297; // @[BTB.scala 105:47:@2009.4]
  wire  _T_1298; // @[BTB.scala 105:47:@2010.4]
  wire  _T_1299; // @[BTB.scala 105:47:@2011.4]
  wire  _T_1300; // @[BTB.scala 105:47:@2012.4]
  wire  _T_1301; // @[BTB.scala 105:47:@2013.4]
  wire  _T_1302; // @[BTB.scala 105:47:@2014.4]
  wire  _T_1303; // @[BTB.scala 105:47:@2015.4]
  wire  _T_1304; // @[BTB.scala 105:47:@2016.4]
  wire  _T_1305; // @[BTB.scala 105:47:@2017.4]
  wire  _T_1306; // @[BTB.scala 105:47:@2018.4]
  wire  _T_1307; // @[BTB.scala 105:47:@2019.4]
  wire  _T_1308; // @[BTB.scala 105:47:@2020.4]
  wire  _T_1309; // @[BTB.scala 105:47:@2021.4]
  wire  _T_1310; // @[BTB.scala 105:47:@2022.4]
  wire  _T_1311; // @[BTB.scala 105:47:@2023.4]
  wire  _T_1312; // @[BTB.scala 105:47:@2024.4]
  wire  _T_1313; // @[BTB.scala 105:47:@2025.4]
  wire  _T_1314; // @[BTB.scala 105:47:@2026.4]
  wire  _T_1315; // @[BTB.scala 105:47:@2027.4]
  wire  _T_1316; // @[BTB.scala 105:47:@2028.4]
  wire  _T_1317; // @[BTB.scala 105:47:@2029.4]
  wire  _T_1318; // @[BTB.scala 105:47:@2030.4]
  wire  _T_1319; // @[BTB.scala 105:47:@2031.4]
  wire  _T_1320; // @[BTB.scala 105:47:@2032.4]
  wire  _T_1321; // @[BTB.scala 105:47:@2033.4]
  wire  _T_1322; // @[BTB.scala 105:47:@2034.4]
  wire  _T_1323; // @[BTB.scala 105:47:@2035.4]
  wire  _T_1324; // @[BTB.scala 105:47:@2036.4]
  wire  _T_1325; // @[BTB.scala 105:47:@2037.4]
  wire  _T_1326; // @[BTB.scala 105:47:@2038.4]
  wire  _T_1327; // @[BTB.scala 105:47:@2039.4]
  wire  _T_1328; // @[BTB.scala 105:47:@2040.4]
  wire  _T_1329; // @[BTB.scala 105:47:@2041.4]
  wire  _T_1330; // @[BTB.scala 105:47:@2042.4]
  wire  _T_1331; // @[BTB.scala 105:47:@2043.4]
  wire  _T_1332; // @[BTB.scala 105:47:@2044.4]
  wire  _T_1333; // @[BTB.scala 105:47:@2045.4]
  wire  _T_1334; // @[BTB.scala 105:47:@2046.4]
  wire  _T_1335; // @[BTB.scala 105:47:@2047.4]
  wire  _T_1336; // @[BTB.scala 105:47:@2048.4]
  wire  _T_1337; // @[BTB.scala 105:47:@2049.4]
  wire  _T_1338; // @[BTB.scala 105:47:@2050.4]
  wire [7:0] _T_1415; // @[BTB.scala 105:62:@2122.4]
  wire [15:0] _T_1423; // @[BTB.scala 105:62:@2130.4]
  wire [7:0] _T_1430; // @[BTB.scala 105:62:@2137.4]
  wire [31:0] _T_1439; // @[BTB.scala 105:62:@2146.4]
  wire [7:0] _T_1446; // @[BTB.scala 105:62:@2153.4]
  wire [15:0] _T_1454; // @[BTB.scala 105:62:@2161.4]
  wire [7:0] _T_1461; // @[BTB.scala 105:62:@2168.4]
  wire [31:0] _T_1470; // @[BTB.scala 105:62:@2177.4]
  wire [63:0] _T_1471; // @[BTB.scala 105:62:@2178.4]
  wire [63:0] predict_1_lookup; // @[BTB.scala 105:69:@2242.4]
  wire  _T_1536; // @[Mux.scala 21:36:@2244.4]
  wire  _T_1537; // @[Mux.scala 21:36:@2245.4]
  wire  _T_1538; // @[Mux.scala 21:36:@2246.4]
  wire  _T_1539; // @[Mux.scala 21:36:@2247.4]
  wire  _T_1540; // @[Mux.scala 21:36:@2248.4]
  wire  _T_1541; // @[Mux.scala 21:36:@2249.4]
  wire  _T_1542; // @[Mux.scala 21:36:@2250.4]
  wire  _T_1543; // @[Mux.scala 21:36:@2251.4]
  wire  _T_1544; // @[Mux.scala 21:36:@2252.4]
  wire  _T_1545; // @[Mux.scala 21:36:@2253.4]
  wire  _T_1546; // @[Mux.scala 21:36:@2254.4]
  wire  _T_1547; // @[Mux.scala 21:36:@2255.4]
  wire  _T_1548; // @[Mux.scala 21:36:@2256.4]
  wire  _T_1549; // @[Mux.scala 21:36:@2257.4]
  wire  _T_1550; // @[Mux.scala 21:36:@2258.4]
  wire  _T_1551; // @[Mux.scala 21:36:@2259.4]
  wire  _T_1552; // @[Mux.scala 21:36:@2260.4]
  wire  _T_1553; // @[Mux.scala 21:36:@2261.4]
  wire  _T_1554; // @[Mux.scala 21:36:@2262.4]
  wire  _T_1555; // @[Mux.scala 21:36:@2263.4]
  wire  _T_1556; // @[Mux.scala 21:36:@2264.4]
  wire  _T_1557; // @[Mux.scala 21:36:@2265.4]
  wire  _T_1558; // @[Mux.scala 21:36:@2266.4]
  wire  _T_1559; // @[Mux.scala 21:36:@2267.4]
  wire  _T_1560; // @[Mux.scala 21:36:@2268.4]
  wire  _T_1561; // @[Mux.scala 21:36:@2269.4]
  wire  _T_1562; // @[Mux.scala 21:36:@2270.4]
  wire  _T_1563; // @[Mux.scala 21:36:@2271.4]
  wire  _T_1564; // @[Mux.scala 21:36:@2272.4]
  wire  _T_1565; // @[Mux.scala 21:36:@2273.4]
  wire  _T_1566; // @[Mux.scala 21:36:@2274.4]
  wire  _T_1567; // @[Mux.scala 21:36:@2275.4]
  wire  _T_1568; // @[Mux.scala 21:36:@2276.4]
  wire  _T_1569; // @[Mux.scala 21:36:@2277.4]
  wire  _T_1570; // @[Mux.scala 21:36:@2278.4]
  wire  _T_1571; // @[Mux.scala 21:36:@2279.4]
  wire  _T_1572; // @[Mux.scala 21:36:@2280.4]
  wire  _T_1573; // @[Mux.scala 21:36:@2281.4]
  wire  _T_1574; // @[Mux.scala 21:36:@2282.4]
  wire  _T_1575; // @[Mux.scala 21:36:@2283.4]
  wire  _T_1576; // @[Mux.scala 21:36:@2284.4]
  wire  _T_1577; // @[Mux.scala 21:36:@2285.4]
  wire  _T_1578; // @[Mux.scala 21:36:@2286.4]
  wire  _T_1579; // @[Mux.scala 21:36:@2287.4]
  wire  _T_1580; // @[Mux.scala 21:36:@2288.4]
  wire  _T_1581; // @[Mux.scala 21:36:@2289.4]
  wire  _T_1582; // @[Mux.scala 21:36:@2290.4]
  wire  _T_1583; // @[Mux.scala 21:36:@2291.4]
  wire  _T_1584; // @[Mux.scala 21:36:@2292.4]
  wire  _T_1585; // @[Mux.scala 21:36:@2293.4]
  wire  _T_1586; // @[Mux.scala 21:36:@2294.4]
  wire  _T_1587; // @[Mux.scala 21:36:@2295.4]
  wire  _T_1588; // @[Mux.scala 21:36:@2296.4]
  wire  _T_1589; // @[Mux.scala 21:36:@2297.4]
  wire  _T_1590; // @[Mux.scala 21:36:@2298.4]
  wire  _T_1591; // @[Mux.scala 21:36:@2299.4]
  wire  _T_1592; // @[Mux.scala 21:36:@2300.4]
  wire  _T_1593; // @[Mux.scala 21:36:@2301.4]
  wire  _T_1594; // @[Mux.scala 21:36:@2302.4]
  wire  _T_1595; // @[Mux.scala 21:36:@2303.4]
  wire  _T_1596; // @[Mux.scala 21:36:@2304.4]
  wire  _T_1597; // @[Mux.scala 21:36:@2305.4]
  wire  _T_1598; // @[Mux.scala 21:36:@2306.4]
  wire  _T_1599; // @[Mux.scala 21:36:@2307.4]
  wire [29:0] _T_1602; // @[Mux.scala 19:72:@2308.4]
  wire [29:0] _T_1604; // @[Mux.scala 19:72:@2309.4]
  wire [29:0] _T_1606; // @[Mux.scala 19:72:@2310.4]
  wire [29:0] _T_1608; // @[Mux.scala 19:72:@2311.4]
  wire [29:0] _T_1610; // @[Mux.scala 19:72:@2312.4]
  wire [29:0] _T_1612; // @[Mux.scala 19:72:@2313.4]
  wire [29:0] _T_1614; // @[Mux.scala 19:72:@2314.4]
  wire [29:0] _T_1616; // @[Mux.scala 19:72:@2315.4]
  wire [29:0] _T_1618; // @[Mux.scala 19:72:@2316.4]
  wire [29:0] _T_1620; // @[Mux.scala 19:72:@2317.4]
  wire [29:0] _T_1622; // @[Mux.scala 19:72:@2318.4]
  wire [29:0] _T_1624; // @[Mux.scala 19:72:@2319.4]
  wire [29:0] _T_1626; // @[Mux.scala 19:72:@2320.4]
  wire [29:0] _T_1628; // @[Mux.scala 19:72:@2321.4]
  wire [29:0] _T_1630; // @[Mux.scala 19:72:@2322.4]
  wire [29:0] _T_1632; // @[Mux.scala 19:72:@2323.4]
  wire [29:0] _T_1634; // @[Mux.scala 19:72:@2324.4]
  wire [29:0] _T_1636; // @[Mux.scala 19:72:@2325.4]
  wire [29:0] _T_1638; // @[Mux.scala 19:72:@2326.4]
  wire [29:0] _T_1640; // @[Mux.scala 19:72:@2327.4]
  wire [29:0] _T_1642; // @[Mux.scala 19:72:@2328.4]
  wire [29:0] _T_1644; // @[Mux.scala 19:72:@2329.4]
  wire [29:0] _T_1646; // @[Mux.scala 19:72:@2330.4]
  wire [29:0] _T_1648; // @[Mux.scala 19:72:@2331.4]
  wire [29:0] _T_1650; // @[Mux.scala 19:72:@2332.4]
  wire [29:0] _T_1652; // @[Mux.scala 19:72:@2333.4]
  wire [29:0] _T_1654; // @[Mux.scala 19:72:@2334.4]
  wire [29:0] _T_1656; // @[Mux.scala 19:72:@2335.4]
  wire [29:0] _T_1658; // @[Mux.scala 19:72:@2336.4]
  wire [29:0] _T_1660; // @[Mux.scala 19:72:@2337.4]
  wire [29:0] _T_1662; // @[Mux.scala 19:72:@2338.4]
  wire [29:0] _T_1664; // @[Mux.scala 19:72:@2339.4]
  wire [29:0] _T_1666; // @[Mux.scala 19:72:@2340.4]
  wire [29:0] _T_1668; // @[Mux.scala 19:72:@2341.4]
  wire [29:0] _T_1670; // @[Mux.scala 19:72:@2342.4]
  wire [29:0] _T_1672; // @[Mux.scala 19:72:@2343.4]
  wire [29:0] _T_1674; // @[Mux.scala 19:72:@2344.4]
  wire [29:0] _T_1676; // @[Mux.scala 19:72:@2345.4]
  wire [29:0] _T_1678; // @[Mux.scala 19:72:@2346.4]
  wire [29:0] _T_1680; // @[Mux.scala 19:72:@2347.4]
  wire [29:0] _T_1682; // @[Mux.scala 19:72:@2348.4]
  wire [29:0] _T_1684; // @[Mux.scala 19:72:@2349.4]
  wire [29:0] _T_1686; // @[Mux.scala 19:72:@2350.4]
  wire [29:0] _T_1688; // @[Mux.scala 19:72:@2351.4]
  wire [29:0] _T_1690; // @[Mux.scala 19:72:@2352.4]
  wire [29:0] _T_1692; // @[Mux.scala 19:72:@2353.4]
  wire [29:0] _T_1694; // @[Mux.scala 19:72:@2354.4]
  wire [29:0] _T_1696; // @[Mux.scala 19:72:@2355.4]
  wire [29:0] _T_1698; // @[Mux.scala 19:72:@2356.4]
  wire [29:0] _T_1700; // @[Mux.scala 19:72:@2357.4]
  wire [29:0] _T_1702; // @[Mux.scala 19:72:@2358.4]
  wire [29:0] _T_1704; // @[Mux.scala 19:72:@2359.4]
  wire [29:0] _T_1706; // @[Mux.scala 19:72:@2360.4]
  wire [29:0] _T_1708; // @[Mux.scala 19:72:@2361.4]
  wire [29:0] _T_1710; // @[Mux.scala 19:72:@2362.4]
  wire [29:0] _T_1712; // @[Mux.scala 19:72:@2363.4]
  wire [29:0] _T_1714; // @[Mux.scala 19:72:@2364.4]
  wire [29:0] _T_1716; // @[Mux.scala 19:72:@2365.4]
  wire [29:0] _T_1718; // @[Mux.scala 19:72:@2366.4]
  wire [29:0] _T_1720; // @[Mux.scala 19:72:@2367.4]
  wire [29:0] _T_1722; // @[Mux.scala 19:72:@2368.4]
  wire [29:0] _T_1724; // @[Mux.scala 19:72:@2369.4]
  wire [29:0] _T_1726; // @[Mux.scala 19:72:@2370.4]
  wire [29:0] _T_1728; // @[Mux.scala 19:72:@2371.4]
  wire [29:0] _T_1729; // @[Mux.scala 19:72:@2372.4]
  wire [29:0] _T_1730; // @[Mux.scala 19:72:@2373.4]
  wire [29:0] _T_1731; // @[Mux.scala 19:72:@2374.4]
  wire [29:0] _T_1732; // @[Mux.scala 19:72:@2375.4]
  wire [29:0] _T_1733; // @[Mux.scala 19:72:@2376.4]
  wire [29:0] _T_1734; // @[Mux.scala 19:72:@2377.4]
  wire [29:0] _T_1735; // @[Mux.scala 19:72:@2378.4]
  wire [29:0] _T_1736; // @[Mux.scala 19:72:@2379.4]
  wire [29:0] _T_1737; // @[Mux.scala 19:72:@2380.4]
  wire [29:0] _T_1738; // @[Mux.scala 19:72:@2381.4]
  wire [29:0] _T_1739; // @[Mux.scala 19:72:@2382.4]
  wire [29:0] _T_1740; // @[Mux.scala 19:72:@2383.4]
  wire [29:0] _T_1741; // @[Mux.scala 19:72:@2384.4]
  wire [29:0] _T_1742; // @[Mux.scala 19:72:@2385.4]
  wire [29:0] _T_1743; // @[Mux.scala 19:72:@2386.4]
  wire [29:0] _T_1744; // @[Mux.scala 19:72:@2387.4]
  wire [29:0] _T_1745; // @[Mux.scala 19:72:@2388.4]
  wire [29:0] _T_1746; // @[Mux.scala 19:72:@2389.4]
  wire [29:0] _T_1747; // @[Mux.scala 19:72:@2390.4]
  wire [29:0] _T_1748; // @[Mux.scala 19:72:@2391.4]
  wire [29:0] _T_1749; // @[Mux.scala 19:72:@2392.4]
  wire [29:0] _T_1750; // @[Mux.scala 19:72:@2393.4]
  wire [29:0] _T_1751; // @[Mux.scala 19:72:@2394.4]
  wire [29:0] _T_1752; // @[Mux.scala 19:72:@2395.4]
  wire [29:0] _T_1753; // @[Mux.scala 19:72:@2396.4]
  wire [29:0] _T_1754; // @[Mux.scala 19:72:@2397.4]
  wire [29:0] _T_1755; // @[Mux.scala 19:72:@2398.4]
  wire [29:0] _T_1756; // @[Mux.scala 19:72:@2399.4]
  wire [29:0] _T_1757; // @[Mux.scala 19:72:@2400.4]
  wire [29:0] _T_1758; // @[Mux.scala 19:72:@2401.4]
  wire [29:0] _T_1759; // @[Mux.scala 19:72:@2402.4]
  wire [29:0] _T_1760; // @[Mux.scala 19:72:@2403.4]
  wire [29:0] _T_1761; // @[Mux.scala 19:72:@2404.4]
  wire [29:0] _T_1762; // @[Mux.scala 19:72:@2405.4]
  wire [29:0] _T_1763; // @[Mux.scala 19:72:@2406.4]
  wire [29:0] _T_1764; // @[Mux.scala 19:72:@2407.4]
  wire [29:0] _T_1765; // @[Mux.scala 19:72:@2408.4]
  wire [29:0] _T_1766; // @[Mux.scala 19:72:@2409.4]
  wire [29:0] _T_1767; // @[Mux.scala 19:72:@2410.4]
  wire [29:0] _T_1768; // @[Mux.scala 19:72:@2411.4]
  wire [29:0] _T_1769; // @[Mux.scala 19:72:@2412.4]
  wire [29:0] _T_1770; // @[Mux.scala 19:72:@2413.4]
  wire [29:0] _T_1771; // @[Mux.scala 19:72:@2414.4]
  wire [29:0] _T_1772; // @[Mux.scala 19:72:@2415.4]
  wire [29:0] _T_1773; // @[Mux.scala 19:72:@2416.4]
  wire [29:0] _T_1774; // @[Mux.scala 19:72:@2417.4]
  wire [29:0] _T_1775; // @[Mux.scala 19:72:@2418.4]
  wire [29:0] _T_1776; // @[Mux.scala 19:72:@2419.4]
  wire [29:0] _T_1777; // @[Mux.scala 19:72:@2420.4]
  wire [29:0] _T_1778; // @[Mux.scala 19:72:@2421.4]
  wire [29:0] _T_1779; // @[Mux.scala 19:72:@2422.4]
  wire [29:0] _T_1780; // @[Mux.scala 19:72:@2423.4]
  wire [29:0] _T_1781; // @[Mux.scala 19:72:@2424.4]
  wire [29:0] _T_1782; // @[Mux.scala 19:72:@2425.4]
  wire [29:0] _T_1783; // @[Mux.scala 19:72:@2426.4]
  wire [29:0] _T_1784; // @[Mux.scala 19:72:@2427.4]
  wire [29:0] _T_1785; // @[Mux.scala 19:72:@2428.4]
  wire [29:0] _T_1786; // @[Mux.scala 19:72:@2429.4]
  wire [29:0] _T_1787; // @[Mux.scala 19:72:@2430.4]
  wire [29:0] _T_1788; // @[Mux.scala 19:72:@2431.4]
  wire [29:0] _T_1789; // @[Mux.scala 19:72:@2432.4]
  wire [29:0] _T_1790; // @[Mux.scala 19:72:@2433.4]
  wire [29:0] _T_1791; // @[Mux.scala 19:72:@2434.4]
  wire [31:0] predict_1_jump_tgt; // @[Cat.scala 30:58:@2437.4]
  wire [1:0] _T_1862; // @[Mux.scala 19:72:@2503.4]
  wire [1:0] _T_1864; // @[Mux.scala 19:72:@2504.4]
  wire [1:0] _T_1866; // @[Mux.scala 19:72:@2505.4]
  wire [1:0] _T_1868; // @[Mux.scala 19:72:@2506.4]
  wire [1:0] _T_1870; // @[Mux.scala 19:72:@2507.4]
  wire [1:0] _T_1872; // @[Mux.scala 19:72:@2508.4]
  wire [1:0] _T_1874; // @[Mux.scala 19:72:@2509.4]
  wire [1:0] _T_1876; // @[Mux.scala 19:72:@2510.4]
  wire [1:0] _T_1878; // @[Mux.scala 19:72:@2511.4]
  wire [1:0] _T_1880; // @[Mux.scala 19:72:@2512.4]
  wire [1:0] _T_1882; // @[Mux.scala 19:72:@2513.4]
  wire [1:0] _T_1884; // @[Mux.scala 19:72:@2514.4]
  wire [1:0] _T_1886; // @[Mux.scala 19:72:@2515.4]
  wire [1:0] _T_1888; // @[Mux.scala 19:72:@2516.4]
  wire [1:0] _T_1890; // @[Mux.scala 19:72:@2517.4]
  wire [1:0] _T_1892; // @[Mux.scala 19:72:@2518.4]
  wire [1:0] _T_1894; // @[Mux.scala 19:72:@2519.4]
  wire [1:0] _T_1896; // @[Mux.scala 19:72:@2520.4]
  wire [1:0] _T_1898; // @[Mux.scala 19:72:@2521.4]
  wire [1:0] _T_1900; // @[Mux.scala 19:72:@2522.4]
  wire [1:0] _T_1902; // @[Mux.scala 19:72:@2523.4]
  wire [1:0] _T_1904; // @[Mux.scala 19:72:@2524.4]
  wire [1:0] _T_1906; // @[Mux.scala 19:72:@2525.4]
  wire [1:0] _T_1908; // @[Mux.scala 19:72:@2526.4]
  wire [1:0] _T_1910; // @[Mux.scala 19:72:@2527.4]
  wire [1:0] _T_1912; // @[Mux.scala 19:72:@2528.4]
  wire [1:0] _T_1914; // @[Mux.scala 19:72:@2529.4]
  wire [1:0] _T_1916; // @[Mux.scala 19:72:@2530.4]
  wire [1:0] _T_1918; // @[Mux.scala 19:72:@2531.4]
  wire [1:0] _T_1920; // @[Mux.scala 19:72:@2532.4]
  wire [1:0] _T_1922; // @[Mux.scala 19:72:@2533.4]
  wire [1:0] _T_1924; // @[Mux.scala 19:72:@2534.4]
  wire [1:0] _T_1926; // @[Mux.scala 19:72:@2535.4]
  wire [1:0] _T_1928; // @[Mux.scala 19:72:@2536.4]
  wire [1:0] _T_1930; // @[Mux.scala 19:72:@2537.4]
  wire [1:0] _T_1932; // @[Mux.scala 19:72:@2538.4]
  wire [1:0] _T_1934; // @[Mux.scala 19:72:@2539.4]
  wire [1:0] _T_1936; // @[Mux.scala 19:72:@2540.4]
  wire [1:0] _T_1938; // @[Mux.scala 19:72:@2541.4]
  wire [1:0] _T_1940; // @[Mux.scala 19:72:@2542.4]
  wire [1:0] _T_1942; // @[Mux.scala 19:72:@2543.4]
  wire [1:0] _T_1944; // @[Mux.scala 19:72:@2544.4]
  wire [1:0] _T_1946; // @[Mux.scala 19:72:@2545.4]
  wire [1:0] _T_1948; // @[Mux.scala 19:72:@2546.4]
  wire [1:0] _T_1950; // @[Mux.scala 19:72:@2547.4]
  wire [1:0] _T_1952; // @[Mux.scala 19:72:@2548.4]
  wire [1:0] _T_1954; // @[Mux.scala 19:72:@2549.4]
  wire [1:0] _T_1956; // @[Mux.scala 19:72:@2550.4]
  wire [1:0] _T_1958; // @[Mux.scala 19:72:@2551.4]
  wire [1:0] _T_1960; // @[Mux.scala 19:72:@2552.4]
  wire [1:0] _T_1962; // @[Mux.scala 19:72:@2553.4]
  wire [1:0] _T_1964; // @[Mux.scala 19:72:@2554.4]
  wire [1:0] _T_1966; // @[Mux.scala 19:72:@2555.4]
  wire [1:0] _T_1968; // @[Mux.scala 19:72:@2556.4]
  wire [1:0] _T_1970; // @[Mux.scala 19:72:@2557.4]
  wire [1:0] _T_1972; // @[Mux.scala 19:72:@2558.4]
  wire [1:0] _T_1974; // @[Mux.scala 19:72:@2559.4]
  wire [1:0] _T_1976; // @[Mux.scala 19:72:@2560.4]
  wire [1:0] _T_1978; // @[Mux.scala 19:72:@2561.4]
  wire [1:0] _T_1980; // @[Mux.scala 19:72:@2562.4]
  wire [1:0] _T_1982; // @[Mux.scala 19:72:@2563.4]
  wire [1:0] _T_1984; // @[Mux.scala 19:72:@2564.4]
  wire [1:0] _T_1986; // @[Mux.scala 19:72:@2565.4]
  wire [1:0] _T_1988; // @[Mux.scala 19:72:@2566.4]
  wire [1:0] _T_1989; // @[Mux.scala 19:72:@2567.4]
  wire [1:0] _T_1990; // @[Mux.scala 19:72:@2568.4]
  wire [1:0] _T_1991; // @[Mux.scala 19:72:@2569.4]
  wire [1:0] _T_1992; // @[Mux.scala 19:72:@2570.4]
  wire [1:0] _T_1993; // @[Mux.scala 19:72:@2571.4]
  wire [1:0] _T_1994; // @[Mux.scala 19:72:@2572.4]
  wire [1:0] _T_1995; // @[Mux.scala 19:72:@2573.4]
  wire [1:0] _T_1996; // @[Mux.scala 19:72:@2574.4]
  wire [1:0] _T_1997; // @[Mux.scala 19:72:@2575.4]
  wire [1:0] _T_1998; // @[Mux.scala 19:72:@2576.4]
  wire [1:0] _T_1999; // @[Mux.scala 19:72:@2577.4]
  wire [1:0] _T_2000; // @[Mux.scala 19:72:@2578.4]
  wire [1:0] _T_2001; // @[Mux.scala 19:72:@2579.4]
  wire [1:0] _T_2002; // @[Mux.scala 19:72:@2580.4]
  wire [1:0] _T_2003; // @[Mux.scala 19:72:@2581.4]
  wire [1:0] _T_2004; // @[Mux.scala 19:72:@2582.4]
  wire [1:0] _T_2005; // @[Mux.scala 19:72:@2583.4]
  wire [1:0] _T_2006; // @[Mux.scala 19:72:@2584.4]
  wire [1:0] _T_2007; // @[Mux.scala 19:72:@2585.4]
  wire [1:0] _T_2008; // @[Mux.scala 19:72:@2586.4]
  wire [1:0] _T_2009; // @[Mux.scala 19:72:@2587.4]
  wire [1:0] _T_2010; // @[Mux.scala 19:72:@2588.4]
  wire [1:0] _T_2011; // @[Mux.scala 19:72:@2589.4]
  wire [1:0] _T_2012; // @[Mux.scala 19:72:@2590.4]
  wire [1:0] _T_2013; // @[Mux.scala 19:72:@2591.4]
  wire [1:0] _T_2014; // @[Mux.scala 19:72:@2592.4]
  wire [1:0] _T_2015; // @[Mux.scala 19:72:@2593.4]
  wire [1:0] _T_2016; // @[Mux.scala 19:72:@2594.4]
  wire [1:0] _T_2017; // @[Mux.scala 19:72:@2595.4]
  wire [1:0] _T_2018; // @[Mux.scala 19:72:@2596.4]
  wire [1:0] _T_2019; // @[Mux.scala 19:72:@2597.4]
  wire [1:0] _T_2020; // @[Mux.scala 19:72:@2598.4]
  wire [1:0] _T_2021; // @[Mux.scala 19:72:@2599.4]
  wire [1:0] _T_2022; // @[Mux.scala 19:72:@2600.4]
  wire [1:0] _T_2023; // @[Mux.scala 19:72:@2601.4]
  wire [1:0] _T_2024; // @[Mux.scala 19:72:@2602.4]
  wire [1:0] _T_2025; // @[Mux.scala 19:72:@2603.4]
  wire [1:0] _T_2026; // @[Mux.scala 19:72:@2604.4]
  wire [1:0] _T_2027; // @[Mux.scala 19:72:@2605.4]
  wire [1:0] _T_2028; // @[Mux.scala 19:72:@2606.4]
  wire [1:0] _T_2029; // @[Mux.scala 19:72:@2607.4]
  wire [1:0] _T_2030; // @[Mux.scala 19:72:@2608.4]
  wire [1:0] _T_2031; // @[Mux.scala 19:72:@2609.4]
  wire [1:0] _T_2032; // @[Mux.scala 19:72:@2610.4]
  wire [1:0] _T_2033; // @[Mux.scala 19:72:@2611.4]
  wire [1:0] _T_2034; // @[Mux.scala 19:72:@2612.4]
  wire [1:0] _T_2035; // @[Mux.scala 19:72:@2613.4]
  wire [1:0] _T_2036; // @[Mux.scala 19:72:@2614.4]
  wire [1:0] _T_2037; // @[Mux.scala 19:72:@2615.4]
  wire [1:0] _T_2038; // @[Mux.scala 19:72:@2616.4]
  wire [1:0] _T_2039; // @[Mux.scala 19:72:@2617.4]
  wire [1:0] _T_2040; // @[Mux.scala 19:72:@2618.4]
  wire [1:0] _T_2041; // @[Mux.scala 19:72:@2619.4]
  wire [1:0] _T_2042; // @[Mux.scala 19:72:@2620.4]
  wire [1:0] _T_2043; // @[Mux.scala 19:72:@2621.4]
  wire [1:0] _T_2044; // @[Mux.scala 19:72:@2622.4]
  wire [1:0] _T_2045; // @[Mux.scala 19:72:@2623.4]
  wire [1:0] _T_2046; // @[Mux.scala 19:72:@2624.4]
  wire [1:0] _T_2047; // @[Mux.scala 19:72:@2625.4]
  wire [1:0] _T_2048; // @[Mux.scala 19:72:@2626.4]
  wire [1:0] _T_2049; // @[Mux.scala 19:72:@2627.4]
  wire [1:0] _T_2050; // @[Mux.scala 19:72:@2628.4]
  wire [1:0] predict_1_bj_type; // @[Mux.scala 19:72:@2629.4]
  wire [1:0] _T_2120; // @[Mux.scala 19:72:@2697.4]
  wire [1:0] _T_2122; // @[Mux.scala 19:72:@2698.4]
  wire [1:0] _T_2124; // @[Mux.scala 19:72:@2699.4]
  wire [1:0] _T_2126; // @[Mux.scala 19:72:@2700.4]
  wire [1:0] _T_2128; // @[Mux.scala 19:72:@2701.4]
  wire [1:0] _T_2130; // @[Mux.scala 19:72:@2702.4]
  wire [1:0] _T_2132; // @[Mux.scala 19:72:@2703.4]
  wire [1:0] _T_2134; // @[Mux.scala 19:72:@2704.4]
  wire [1:0] _T_2136; // @[Mux.scala 19:72:@2705.4]
  wire [1:0] _T_2138; // @[Mux.scala 19:72:@2706.4]
  wire [1:0] _T_2140; // @[Mux.scala 19:72:@2707.4]
  wire [1:0] _T_2142; // @[Mux.scala 19:72:@2708.4]
  wire [1:0] _T_2144; // @[Mux.scala 19:72:@2709.4]
  wire [1:0] _T_2146; // @[Mux.scala 19:72:@2710.4]
  wire [1:0] _T_2148; // @[Mux.scala 19:72:@2711.4]
  wire [1:0] _T_2150; // @[Mux.scala 19:72:@2712.4]
  wire [1:0] _T_2152; // @[Mux.scala 19:72:@2713.4]
  wire [1:0] _T_2154; // @[Mux.scala 19:72:@2714.4]
  wire [1:0] _T_2156; // @[Mux.scala 19:72:@2715.4]
  wire [1:0] _T_2158; // @[Mux.scala 19:72:@2716.4]
  wire [1:0] _T_2160; // @[Mux.scala 19:72:@2717.4]
  wire [1:0] _T_2162; // @[Mux.scala 19:72:@2718.4]
  wire [1:0] _T_2164; // @[Mux.scala 19:72:@2719.4]
  wire [1:0] _T_2166; // @[Mux.scala 19:72:@2720.4]
  wire [1:0] _T_2168; // @[Mux.scala 19:72:@2721.4]
  wire [1:0] _T_2170; // @[Mux.scala 19:72:@2722.4]
  wire [1:0] _T_2172; // @[Mux.scala 19:72:@2723.4]
  wire [1:0] _T_2174; // @[Mux.scala 19:72:@2724.4]
  wire [1:0] _T_2176; // @[Mux.scala 19:72:@2725.4]
  wire [1:0] _T_2178; // @[Mux.scala 19:72:@2726.4]
  wire [1:0] _T_2180; // @[Mux.scala 19:72:@2727.4]
  wire [1:0] _T_2182; // @[Mux.scala 19:72:@2728.4]
  wire [1:0] _T_2184; // @[Mux.scala 19:72:@2729.4]
  wire [1:0] _T_2186; // @[Mux.scala 19:72:@2730.4]
  wire [1:0] _T_2188; // @[Mux.scala 19:72:@2731.4]
  wire [1:0] _T_2190; // @[Mux.scala 19:72:@2732.4]
  wire [1:0] _T_2192; // @[Mux.scala 19:72:@2733.4]
  wire [1:0] _T_2194; // @[Mux.scala 19:72:@2734.4]
  wire [1:0] _T_2196; // @[Mux.scala 19:72:@2735.4]
  wire [1:0] _T_2198; // @[Mux.scala 19:72:@2736.4]
  wire [1:0] _T_2200; // @[Mux.scala 19:72:@2737.4]
  wire [1:0] _T_2202; // @[Mux.scala 19:72:@2738.4]
  wire [1:0] _T_2204; // @[Mux.scala 19:72:@2739.4]
  wire [1:0] _T_2206; // @[Mux.scala 19:72:@2740.4]
  wire [1:0] _T_2208; // @[Mux.scala 19:72:@2741.4]
  wire [1:0] _T_2210; // @[Mux.scala 19:72:@2742.4]
  wire [1:0] _T_2212; // @[Mux.scala 19:72:@2743.4]
  wire [1:0] _T_2214; // @[Mux.scala 19:72:@2744.4]
  wire [1:0] _T_2216; // @[Mux.scala 19:72:@2745.4]
  wire [1:0] _T_2218; // @[Mux.scala 19:72:@2746.4]
  wire [1:0] _T_2220; // @[Mux.scala 19:72:@2747.4]
  wire [1:0] _T_2222; // @[Mux.scala 19:72:@2748.4]
  wire [1:0] _T_2224; // @[Mux.scala 19:72:@2749.4]
  wire [1:0] _T_2226; // @[Mux.scala 19:72:@2750.4]
  wire [1:0] _T_2228; // @[Mux.scala 19:72:@2751.4]
  wire [1:0] _T_2230; // @[Mux.scala 19:72:@2752.4]
  wire [1:0] _T_2232; // @[Mux.scala 19:72:@2753.4]
  wire [1:0] _T_2234; // @[Mux.scala 19:72:@2754.4]
  wire [1:0] _T_2236; // @[Mux.scala 19:72:@2755.4]
  wire [1:0] _T_2238; // @[Mux.scala 19:72:@2756.4]
  wire [1:0] _T_2240; // @[Mux.scala 19:72:@2757.4]
  wire [1:0] _T_2242; // @[Mux.scala 19:72:@2758.4]
  wire [1:0] _T_2244; // @[Mux.scala 19:72:@2759.4]
  wire [1:0] _T_2246; // @[Mux.scala 19:72:@2760.4]
  wire [1:0] _T_2247; // @[Mux.scala 19:72:@2761.4]
  wire [1:0] _T_2248; // @[Mux.scala 19:72:@2762.4]
  wire [1:0] _T_2249; // @[Mux.scala 19:72:@2763.4]
  wire [1:0] _T_2250; // @[Mux.scala 19:72:@2764.4]
  wire [1:0] _T_2251; // @[Mux.scala 19:72:@2765.4]
  wire [1:0] _T_2252; // @[Mux.scala 19:72:@2766.4]
  wire [1:0] _T_2253; // @[Mux.scala 19:72:@2767.4]
  wire [1:0] _T_2254; // @[Mux.scala 19:72:@2768.4]
  wire [1:0] _T_2255; // @[Mux.scala 19:72:@2769.4]
  wire [1:0] _T_2256; // @[Mux.scala 19:72:@2770.4]
  wire [1:0] _T_2257; // @[Mux.scala 19:72:@2771.4]
  wire [1:0] _T_2258; // @[Mux.scala 19:72:@2772.4]
  wire [1:0] _T_2259; // @[Mux.scala 19:72:@2773.4]
  wire [1:0] _T_2260; // @[Mux.scala 19:72:@2774.4]
  wire [1:0] _T_2261; // @[Mux.scala 19:72:@2775.4]
  wire [1:0] _T_2262; // @[Mux.scala 19:72:@2776.4]
  wire [1:0] _T_2263; // @[Mux.scala 19:72:@2777.4]
  wire [1:0] _T_2264; // @[Mux.scala 19:72:@2778.4]
  wire [1:0] _T_2265; // @[Mux.scala 19:72:@2779.4]
  wire [1:0] _T_2266; // @[Mux.scala 19:72:@2780.4]
  wire [1:0] _T_2267; // @[Mux.scala 19:72:@2781.4]
  wire [1:0] _T_2268; // @[Mux.scala 19:72:@2782.4]
  wire [1:0] _T_2269; // @[Mux.scala 19:72:@2783.4]
  wire [1:0] _T_2270; // @[Mux.scala 19:72:@2784.4]
  wire [1:0] _T_2271; // @[Mux.scala 19:72:@2785.4]
  wire [1:0] _T_2272; // @[Mux.scala 19:72:@2786.4]
  wire [1:0] _T_2273; // @[Mux.scala 19:72:@2787.4]
  wire [1:0] _T_2274; // @[Mux.scala 19:72:@2788.4]
  wire [1:0] _T_2275; // @[Mux.scala 19:72:@2789.4]
  wire [1:0] _T_2276; // @[Mux.scala 19:72:@2790.4]
  wire [1:0] _T_2277; // @[Mux.scala 19:72:@2791.4]
  wire [1:0] _T_2278; // @[Mux.scala 19:72:@2792.4]
  wire [1:0] _T_2279; // @[Mux.scala 19:72:@2793.4]
  wire [1:0] _T_2280; // @[Mux.scala 19:72:@2794.4]
  wire [1:0] _T_2281; // @[Mux.scala 19:72:@2795.4]
  wire [1:0] _T_2282; // @[Mux.scala 19:72:@2796.4]
  wire [1:0] _T_2283; // @[Mux.scala 19:72:@2797.4]
  wire [1:0] _T_2284; // @[Mux.scala 19:72:@2798.4]
  wire [1:0] _T_2285; // @[Mux.scala 19:72:@2799.4]
  wire [1:0] _T_2286; // @[Mux.scala 19:72:@2800.4]
  wire [1:0] _T_2287; // @[Mux.scala 19:72:@2801.4]
  wire [1:0] _T_2288; // @[Mux.scala 19:72:@2802.4]
  wire [1:0] _T_2289; // @[Mux.scala 19:72:@2803.4]
  wire [1:0] _T_2290; // @[Mux.scala 19:72:@2804.4]
  wire [1:0] _T_2291; // @[Mux.scala 19:72:@2805.4]
  wire [1:0] _T_2292; // @[Mux.scala 19:72:@2806.4]
  wire [1:0] _T_2293; // @[Mux.scala 19:72:@2807.4]
  wire [1:0] _T_2294; // @[Mux.scala 19:72:@2808.4]
  wire [1:0] _T_2295; // @[Mux.scala 19:72:@2809.4]
  wire [1:0] _T_2296; // @[Mux.scala 19:72:@2810.4]
  wire [1:0] _T_2297; // @[Mux.scala 19:72:@2811.4]
  wire [1:0] _T_2298; // @[Mux.scala 19:72:@2812.4]
  wire [1:0] _T_2299; // @[Mux.scala 19:72:@2813.4]
  wire [1:0] _T_2300; // @[Mux.scala 19:72:@2814.4]
  wire [1:0] _T_2301; // @[Mux.scala 19:72:@2815.4]
  wire [1:0] _T_2302; // @[Mux.scala 19:72:@2816.4]
  wire [1:0] _T_2303; // @[Mux.scala 19:72:@2817.4]
  wire [1:0] _T_2304; // @[Mux.scala 19:72:@2818.4]
  wire [1:0] _T_2305; // @[Mux.scala 19:72:@2819.4]
  wire [1:0] _T_2306; // @[Mux.scala 19:72:@2820.4]
  wire [1:0] _T_2307; // @[Mux.scala 19:72:@2821.4]
  wire [1:0] _T_2308; // @[Mux.scala 19:72:@2822.4]
  wire [1:0] predict_1_h_count; // @[Mux.scala 19:72:@2823.4]
  wire [9:0] _T_2313; // @[BTB.scala 110:54:@2828.4]
  wire [9:0] predict_1_gshxor; // @[BTB.scala 110:44:@2829.4]
  wire [1:0] predict_1_gshare; // @[BTB.scala 98:21:@1087.4 BTB.scala 112:25:@2834.4]
  wire  _T_2318; // @[BTB.scala 47:40:@2836.4]
  wire  _T_2319; // @[BTB.scala 47:52:@2837.4]
  wire  predict_1_select; // @[BTB.scala 98:21:@1087.4 BTB.scala 111:25:@2832.4]
  wire  _T_2320; // @[BTB.scala 47:25:@2838.4]
  wire [9:0] predict_1_history; // @[Cat.scala 30:58:@2839.4]
  wire  _T_2323; // @[BTB.scala 40:28:@2841.4]
  wire  _T_2327; // @[BTB.scala 49:42:@2844.4]
  wire  _T_2331; // @[BTB.scala 49:63:@2848.4]
  wire  _T_2332; // @[BTB.scala 49:30:@2849.4]
  wire  _T_2337; // @[BTB.scala 119:54:@2856.4]
  wire [31:0] _T_2347; // @[BTB.scala 120:34:@2864.4]
  reg  shift_reg; // @[BTB.scala 123:23:@2867.4]
  reg [31:0] _RAND_323;
  wire  shift_wire; // @[BTB.scala 124:30:@2868.4]
  wire  _T_2351; // @[BTB.scala 126:22:@2870.6]
  wire [8:0] _T_2352; // @[BTB.scala 127:44:@2872.8]
  wire [9:0] _T_2353; // @[Cat.scala 30:58:@2873.8]
  wire [9:0] _GEN_0; // @[BTB.scala 126:44:@2871.6]
  wire  _T_2355; // @[BTB.scala 46:30:@2882.8]
  wire  _T_2360; // @[BTB.scala 132:38:@2886.8]
  wire  _T_2362; // @[BTB.scala 132:18:@2887.8]
  wire  _T_2364; // @[BTB.scala 46:30:@2888.8]
  wire  _T_2366; // @[BTB.scala 132:79:@2889.8]
  wire  _T_2367; // @[BTB.scala 132:76:@2890.8]
  wire [9:0] _T_2370; // @[Cat.scala 30:58:@2894.10]
  wire [8:0] _T_2380; // @[BTB.scala 137:45:@2906.14]
  wire [9:0] _T_2384; // @[Cat.scala 30:58:@2910.14]
  wire [9:0] _GEN_1; // @[BTB.scala 136:32:@2905.12]
  wire [9:0] _GEN_2; // @[BTB.scala 141:35:@2919.12]
  wire [9:0] _GEN_3; // @[BTB.scala 135:72:@2903.10]
  wire [9:0] _GEN_4; // @[BTB.scala 133:23:@2892.8]
  wire  _GEN_5; // @[BTB.scala 131:30:@2881.6]
  wire [9:0] _GEN_6; // @[BTB.scala 131:30:@2881.6]
  wire [9:0] _GEN_7; // @[BTB.scala 125:25:@2869.4]
  reg  fb_reg_valid; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_324;
  reg  fb_reg_miss; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_325;
  reg  fb_reg_redirect; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_326;
  reg [1:0] fb_reg_btb_type; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_327;
  reg [29:0] fb_reg_pc; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_328;
  reg [29:0] fb_reg_tgt; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_329;
  reg  fb_reg_diff; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_330;
  reg [9:0] fb_reg_gshxor; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_331;
  reg [5:0] fb_reg_lfsr; // @[BTB.scala 146:23:@2933.4]
  reg [31:0] _RAND_332;
  wire [29:0] _T_2393; // @[BTB.scala 176:35:@2936.4]
  wire [29:0] _T_2394; // @[BTB.scala 177:37:@2938.4]
  wire [9:0] _T_2396; // @[BTB.scala 181:62:@2944.4]
  wire [9:0] _T_2397; // @[BTB.scala 181:47:@2945.4]
  wire  _T_2398; // @[BTB.scala 160:22:@2947.4]
  wire  _T_2399; // @[BTB.scala 160:32:@2948.4]
  wire  _T_2400; // @[BTB.scala 160:26:@2949.4]
  wire [4:0] _T_2401; // @[BTB.scala 160:41:@2950.4]
  wire [5:0] _T_2402; // @[Cat.scala 30:58:@2951.4]
  wire  _T_2404; // @[BTB.scala 192:44:@2954.4]
  wire  _T_2405; // @[BTB.scala 192:44:@2955.4]
  wire  _T_2406; // @[BTB.scala 192:44:@2956.4]
  wire  _T_2407; // @[BTB.scala 192:44:@2957.4]
  wire  _T_2408; // @[BTB.scala 192:44:@2958.4]
  wire  _T_2409; // @[BTB.scala 192:44:@2959.4]
  wire  _T_2410; // @[BTB.scala 192:44:@2960.4]
  wire  _T_2411; // @[BTB.scala 192:44:@2961.4]
  wire  _T_2412; // @[BTB.scala 192:44:@2962.4]
  wire  _T_2413; // @[BTB.scala 192:44:@2963.4]
  wire  _T_2414; // @[BTB.scala 192:44:@2964.4]
  wire  _T_2415; // @[BTB.scala 192:44:@2965.4]
  wire  _T_2416; // @[BTB.scala 192:44:@2966.4]
  wire  _T_2417; // @[BTB.scala 192:44:@2967.4]
  wire  _T_2418; // @[BTB.scala 192:44:@2968.4]
  wire  _T_2419; // @[BTB.scala 192:44:@2969.4]
  wire  _T_2420; // @[BTB.scala 192:44:@2970.4]
  wire  _T_2421; // @[BTB.scala 192:44:@2971.4]
  wire  _T_2422; // @[BTB.scala 192:44:@2972.4]
  wire  _T_2423; // @[BTB.scala 192:44:@2973.4]
  wire  _T_2424; // @[BTB.scala 192:44:@2974.4]
  wire  _T_2425; // @[BTB.scala 192:44:@2975.4]
  wire  _T_2426; // @[BTB.scala 192:44:@2976.4]
  wire  _T_2427; // @[BTB.scala 192:44:@2977.4]
  wire  _T_2428; // @[BTB.scala 192:44:@2978.4]
  wire  _T_2429; // @[BTB.scala 192:44:@2979.4]
  wire  _T_2430; // @[BTB.scala 192:44:@2980.4]
  wire  _T_2431; // @[BTB.scala 192:44:@2981.4]
  wire  _T_2432; // @[BTB.scala 192:44:@2982.4]
  wire  _T_2433; // @[BTB.scala 192:44:@2983.4]
  wire  _T_2434; // @[BTB.scala 192:44:@2984.4]
  wire  _T_2435; // @[BTB.scala 192:44:@2985.4]
  wire  _T_2436; // @[BTB.scala 192:44:@2986.4]
  wire  _T_2437; // @[BTB.scala 192:44:@2987.4]
  wire  _T_2438; // @[BTB.scala 192:44:@2988.4]
  wire  _T_2439; // @[BTB.scala 192:44:@2989.4]
  wire  _T_2440; // @[BTB.scala 192:44:@2990.4]
  wire  _T_2441; // @[BTB.scala 192:44:@2991.4]
  wire  _T_2442; // @[BTB.scala 192:44:@2992.4]
  wire  _T_2443; // @[BTB.scala 192:44:@2993.4]
  wire  _T_2444; // @[BTB.scala 192:44:@2994.4]
  wire  _T_2445; // @[BTB.scala 192:44:@2995.4]
  wire  _T_2446; // @[BTB.scala 192:44:@2996.4]
  wire  _T_2447; // @[BTB.scala 192:44:@2997.4]
  wire  _T_2448; // @[BTB.scala 192:44:@2998.4]
  wire  _T_2449; // @[BTB.scala 192:44:@2999.4]
  wire  _T_2450; // @[BTB.scala 192:44:@3000.4]
  wire  _T_2451; // @[BTB.scala 192:44:@3001.4]
  wire  _T_2452; // @[BTB.scala 192:44:@3002.4]
  wire  _T_2453; // @[BTB.scala 192:44:@3003.4]
  wire  _T_2454; // @[BTB.scala 192:44:@3004.4]
  wire  _T_2455; // @[BTB.scala 192:44:@3005.4]
  wire  _T_2456; // @[BTB.scala 192:44:@3006.4]
  wire  _T_2457; // @[BTB.scala 192:44:@3007.4]
  wire  _T_2458; // @[BTB.scala 192:44:@3008.4]
  wire  _T_2459; // @[BTB.scala 192:44:@3009.4]
  wire  _T_2460; // @[BTB.scala 192:44:@3010.4]
  wire  _T_2461; // @[BTB.scala 192:44:@3011.4]
  wire  _T_2462; // @[BTB.scala 192:44:@3012.4]
  wire  _T_2463; // @[BTB.scala 192:44:@3013.4]
  wire  _T_2464; // @[BTB.scala 192:44:@3014.4]
  wire  _T_2465; // @[BTB.scala 192:44:@3015.4]
  wire  _T_2466; // @[BTB.scala 192:44:@3016.4]
  wire  _T_2467; // @[BTB.scala 192:44:@3017.4]
  wire [7:0] _T_2544; // @[BTB.scala 192:60:@3089.4]
  wire [15:0] _T_2552; // @[BTB.scala 192:60:@3097.4]
  wire [7:0] _T_2559; // @[BTB.scala 192:60:@3104.4]
  wire [31:0] _T_2568; // @[BTB.scala 192:60:@3113.4]
  wire [7:0] _T_2575; // @[BTB.scala 192:60:@3120.4]
  wire [15:0] _T_2583; // @[BTB.scala 192:60:@3128.4]
  wire [7:0] _T_2590; // @[BTB.scala 192:60:@3135.4]
  wire [31:0] _T_2599; // @[BTB.scala 192:60:@3144.4]
  wire [63:0] _T_2600; // @[BTB.scala 192:60:@3145.4]
  wire [63:0] feedback_lookup; // @[BTB.scala 192:67:@3209.4]
  wire  _T_2665; // @[Mux.scala 21:36:@3211.4]
  wire  _T_2666; // @[Mux.scala 21:36:@3212.4]
  wire  _T_2667; // @[Mux.scala 21:36:@3213.4]
  wire  _T_2668; // @[Mux.scala 21:36:@3214.4]
  wire  _T_2669; // @[Mux.scala 21:36:@3215.4]
  wire  _T_2670; // @[Mux.scala 21:36:@3216.4]
  wire  _T_2671; // @[Mux.scala 21:36:@3217.4]
  wire  _T_2672; // @[Mux.scala 21:36:@3218.4]
  wire  _T_2673; // @[Mux.scala 21:36:@3219.4]
  wire  _T_2674; // @[Mux.scala 21:36:@3220.4]
  wire  _T_2675; // @[Mux.scala 21:36:@3221.4]
  wire  _T_2676; // @[Mux.scala 21:36:@3222.4]
  wire  _T_2677; // @[Mux.scala 21:36:@3223.4]
  wire  _T_2678; // @[Mux.scala 21:36:@3224.4]
  wire  _T_2679; // @[Mux.scala 21:36:@3225.4]
  wire  _T_2680; // @[Mux.scala 21:36:@3226.4]
  wire  _T_2681; // @[Mux.scala 21:36:@3227.4]
  wire  _T_2682; // @[Mux.scala 21:36:@3228.4]
  wire  _T_2683; // @[Mux.scala 21:36:@3229.4]
  wire  _T_2684; // @[Mux.scala 21:36:@3230.4]
  wire  _T_2685; // @[Mux.scala 21:36:@3231.4]
  wire  _T_2686; // @[Mux.scala 21:36:@3232.4]
  wire  _T_2687; // @[Mux.scala 21:36:@3233.4]
  wire  _T_2688; // @[Mux.scala 21:36:@3234.4]
  wire  _T_2689; // @[Mux.scala 21:36:@3235.4]
  wire  _T_2690; // @[Mux.scala 21:36:@3236.4]
  wire  _T_2691; // @[Mux.scala 21:36:@3237.4]
  wire  _T_2692; // @[Mux.scala 21:36:@3238.4]
  wire  _T_2693; // @[Mux.scala 21:36:@3239.4]
  wire  _T_2694; // @[Mux.scala 21:36:@3240.4]
  wire  _T_2695; // @[Mux.scala 21:36:@3241.4]
  wire  _T_2696; // @[Mux.scala 21:36:@3242.4]
  wire  _T_2697; // @[Mux.scala 21:36:@3243.4]
  wire  _T_2698; // @[Mux.scala 21:36:@3244.4]
  wire  _T_2699; // @[Mux.scala 21:36:@3245.4]
  wire  _T_2700; // @[Mux.scala 21:36:@3246.4]
  wire  _T_2701; // @[Mux.scala 21:36:@3247.4]
  wire  _T_2702; // @[Mux.scala 21:36:@3248.4]
  wire  _T_2703; // @[Mux.scala 21:36:@3249.4]
  wire  _T_2704; // @[Mux.scala 21:36:@3250.4]
  wire  _T_2705; // @[Mux.scala 21:36:@3251.4]
  wire  _T_2706; // @[Mux.scala 21:36:@3252.4]
  wire  _T_2707; // @[Mux.scala 21:36:@3253.4]
  wire  _T_2708; // @[Mux.scala 21:36:@3254.4]
  wire  _T_2709; // @[Mux.scala 21:36:@3255.4]
  wire  _T_2710; // @[Mux.scala 21:36:@3256.4]
  wire  _T_2711; // @[Mux.scala 21:36:@3257.4]
  wire  _T_2712; // @[Mux.scala 21:36:@3258.4]
  wire  _T_2713; // @[Mux.scala 21:36:@3259.4]
  wire  _T_2714; // @[Mux.scala 21:36:@3260.4]
  wire  _T_2715; // @[Mux.scala 21:36:@3261.4]
  wire  _T_2716; // @[Mux.scala 21:36:@3262.4]
  wire  _T_2717; // @[Mux.scala 21:36:@3263.4]
  wire  _T_2718; // @[Mux.scala 21:36:@3264.4]
  wire  _T_2719; // @[Mux.scala 21:36:@3265.4]
  wire  _T_2720; // @[Mux.scala 21:36:@3266.4]
  wire  _T_2721; // @[Mux.scala 21:36:@3267.4]
  wire  _T_2722; // @[Mux.scala 21:36:@3268.4]
  wire  _T_2723; // @[Mux.scala 21:36:@3269.4]
  wire  _T_2724; // @[Mux.scala 21:36:@3270.4]
  wire  _T_2725; // @[Mux.scala 21:36:@3271.4]
  wire  _T_2726; // @[Mux.scala 21:36:@3272.4]
  wire  _T_2727; // @[Mux.scala 21:36:@3273.4]
  wire  _T_2728; // @[Mux.scala 21:36:@3274.4]
  wire [1:0] _T_2731; // @[Mux.scala 19:72:@3275.4]
  wire [1:0] _T_2733; // @[Mux.scala 19:72:@3276.4]
  wire [1:0] _T_2735; // @[Mux.scala 19:72:@3277.4]
  wire [1:0] _T_2737; // @[Mux.scala 19:72:@3278.4]
  wire [1:0] _T_2739; // @[Mux.scala 19:72:@3279.4]
  wire [1:0] _T_2741; // @[Mux.scala 19:72:@3280.4]
  wire [1:0] _T_2743; // @[Mux.scala 19:72:@3281.4]
  wire [1:0] _T_2745; // @[Mux.scala 19:72:@3282.4]
  wire [1:0] _T_2747; // @[Mux.scala 19:72:@3283.4]
  wire [1:0] _T_2749; // @[Mux.scala 19:72:@3284.4]
  wire [1:0] _T_2751; // @[Mux.scala 19:72:@3285.4]
  wire [1:0] _T_2753; // @[Mux.scala 19:72:@3286.4]
  wire [1:0] _T_2755; // @[Mux.scala 19:72:@3287.4]
  wire [1:0] _T_2757; // @[Mux.scala 19:72:@3288.4]
  wire [1:0] _T_2759; // @[Mux.scala 19:72:@3289.4]
  wire [1:0] _T_2761; // @[Mux.scala 19:72:@3290.4]
  wire [1:0] _T_2763; // @[Mux.scala 19:72:@3291.4]
  wire [1:0] _T_2765; // @[Mux.scala 19:72:@3292.4]
  wire [1:0] _T_2767; // @[Mux.scala 19:72:@3293.4]
  wire [1:0] _T_2769; // @[Mux.scala 19:72:@3294.4]
  wire [1:0] _T_2771; // @[Mux.scala 19:72:@3295.4]
  wire [1:0] _T_2773; // @[Mux.scala 19:72:@3296.4]
  wire [1:0] _T_2775; // @[Mux.scala 19:72:@3297.4]
  wire [1:0] _T_2777; // @[Mux.scala 19:72:@3298.4]
  wire [1:0] _T_2779; // @[Mux.scala 19:72:@3299.4]
  wire [1:0] _T_2781; // @[Mux.scala 19:72:@3300.4]
  wire [1:0] _T_2783; // @[Mux.scala 19:72:@3301.4]
  wire [1:0] _T_2785; // @[Mux.scala 19:72:@3302.4]
  wire [1:0] _T_2787; // @[Mux.scala 19:72:@3303.4]
  wire [1:0] _T_2789; // @[Mux.scala 19:72:@3304.4]
  wire [1:0] _T_2791; // @[Mux.scala 19:72:@3305.4]
  wire [1:0] _T_2793; // @[Mux.scala 19:72:@3306.4]
  wire [1:0] _T_2795; // @[Mux.scala 19:72:@3307.4]
  wire [1:0] _T_2797; // @[Mux.scala 19:72:@3308.4]
  wire [1:0] _T_2799; // @[Mux.scala 19:72:@3309.4]
  wire [1:0] _T_2801; // @[Mux.scala 19:72:@3310.4]
  wire [1:0] _T_2803; // @[Mux.scala 19:72:@3311.4]
  wire [1:0] _T_2805; // @[Mux.scala 19:72:@3312.4]
  wire [1:0] _T_2807; // @[Mux.scala 19:72:@3313.4]
  wire [1:0] _T_2809; // @[Mux.scala 19:72:@3314.4]
  wire [1:0] _T_2811; // @[Mux.scala 19:72:@3315.4]
  wire [1:0] _T_2813; // @[Mux.scala 19:72:@3316.4]
  wire [1:0] _T_2815; // @[Mux.scala 19:72:@3317.4]
  wire [1:0] _T_2817; // @[Mux.scala 19:72:@3318.4]
  wire [1:0] _T_2819; // @[Mux.scala 19:72:@3319.4]
  wire [1:0] _T_2821; // @[Mux.scala 19:72:@3320.4]
  wire [1:0] _T_2823; // @[Mux.scala 19:72:@3321.4]
  wire [1:0] _T_2825; // @[Mux.scala 19:72:@3322.4]
  wire [1:0] _T_2827; // @[Mux.scala 19:72:@3323.4]
  wire [1:0] _T_2829; // @[Mux.scala 19:72:@3324.4]
  wire [1:0] _T_2831; // @[Mux.scala 19:72:@3325.4]
  wire [1:0] _T_2833; // @[Mux.scala 19:72:@3326.4]
  wire [1:0] _T_2835; // @[Mux.scala 19:72:@3327.4]
  wire [1:0] _T_2837; // @[Mux.scala 19:72:@3328.4]
  wire [1:0] _T_2839; // @[Mux.scala 19:72:@3329.4]
  wire [1:0] _T_2841; // @[Mux.scala 19:72:@3330.4]
  wire [1:0] _T_2843; // @[Mux.scala 19:72:@3331.4]
  wire [1:0] _T_2845; // @[Mux.scala 19:72:@3332.4]
  wire [1:0] _T_2847; // @[Mux.scala 19:72:@3333.4]
  wire [1:0] _T_2849; // @[Mux.scala 19:72:@3334.4]
  wire [1:0] _T_2851; // @[Mux.scala 19:72:@3335.4]
  wire [1:0] _T_2853; // @[Mux.scala 19:72:@3336.4]
  wire [1:0] _T_2855; // @[Mux.scala 19:72:@3337.4]
  wire [1:0] _T_2857; // @[Mux.scala 19:72:@3338.4]
  wire [1:0] _T_2858; // @[Mux.scala 19:72:@3339.4]
  wire [1:0] _T_2859; // @[Mux.scala 19:72:@3340.4]
  wire [1:0] _T_2860; // @[Mux.scala 19:72:@3341.4]
  wire [1:0] _T_2861; // @[Mux.scala 19:72:@3342.4]
  wire [1:0] _T_2862; // @[Mux.scala 19:72:@3343.4]
  wire [1:0] _T_2863; // @[Mux.scala 19:72:@3344.4]
  wire [1:0] _T_2864; // @[Mux.scala 19:72:@3345.4]
  wire [1:0] _T_2865; // @[Mux.scala 19:72:@3346.4]
  wire [1:0] _T_2866; // @[Mux.scala 19:72:@3347.4]
  wire [1:0] _T_2867; // @[Mux.scala 19:72:@3348.4]
  wire [1:0] _T_2868; // @[Mux.scala 19:72:@3349.4]
  wire [1:0] _T_2869; // @[Mux.scala 19:72:@3350.4]
  wire [1:0] _T_2870; // @[Mux.scala 19:72:@3351.4]
  wire [1:0] _T_2871; // @[Mux.scala 19:72:@3352.4]
  wire [1:0] _T_2872; // @[Mux.scala 19:72:@3353.4]
  wire [1:0] _T_2873; // @[Mux.scala 19:72:@3354.4]
  wire [1:0] _T_2874; // @[Mux.scala 19:72:@3355.4]
  wire [1:0] _T_2875; // @[Mux.scala 19:72:@3356.4]
  wire [1:0] _T_2876; // @[Mux.scala 19:72:@3357.4]
  wire [1:0] _T_2877; // @[Mux.scala 19:72:@3358.4]
  wire [1:0] _T_2878; // @[Mux.scala 19:72:@3359.4]
  wire [1:0] _T_2879; // @[Mux.scala 19:72:@3360.4]
  wire [1:0] _T_2880; // @[Mux.scala 19:72:@3361.4]
  wire [1:0] _T_2881; // @[Mux.scala 19:72:@3362.4]
  wire [1:0] _T_2882; // @[Mux.scala 19:72:@3363.4]
  wire [1:0] _T_2883; // @[Mux.scala 19:72:@3364.4]
  wire [1:0] _T_2884; // @[Mux.scala 19:72:@3365.4]
  wire [1:0] _T_2885; // @[Mux.scala 19:72:@3366.4]
  wire [1:0] _T_2886; // @[Mux.scala 19:72:@3367.4]
  wire [1:0] _T_2887; // @[Mux.scala 19:72:@3368.4]
  wire [1:0] _T_2888; // @[Mux.scala 19:72:@3369.4]
  wire [1:0] _T_2889; // @[Mux.scala 19:72:@3370.4]
  wire [1:0] _T_2890; // @[Mux.scala 19:72:@3371.4]
  wire [1:0] _T_2891; // @[Mux.scala 19:72:@3372.4]
  wire [1:0] _T_2892; // @[Mux.scala 19:72:@3373.4]
  wire [1:0] _T_2893; // @[Mux.scala 19:72:@3374.4]
  wire [1:0] _T_2894; // @[Mux.scala 19:72:@3375.4]
  wire [1:0] _T_2895; // @[Mux.scala 19:72:@3376.4]
  wire [1:0] _T_2896; // @[Mux.scala 19:72:@3377.4]
  wire [1:0] _T_2897; // @[Mux.scala 19:72:@3378.4]
  wire [1:0] _T_2898; // @[Mux.scala 19:72:@3379.4]
  wire [1:0] _T_2899; // @[Mux.scala 19:72:@3380.4]
  wire [1:0] _T_2900; // @[Mux.scala 19:72:@3381.4]
  wire [1:0] _T_2901; // @[Mux.scala 19:72:@3382.4]
  wire [1:0] _T_2902; // @[Mux.scala 19:72:@3383.4]
  wire [1:0] _T_2903; // @[Mux.scala 19:72:@3384.4]
  wire [1:0] _T_2904; // @[Mux.scala 19:72:@3385.4]
  wire [1:0] _T_2905; // @[Mux.scala 19:72:@3386.4]
  wire [1:0] _T_2906; // @[Mux.scala 19:72:@3387.4]
  wire [1:0] _T_2907; // @[Mux.scala 19:72:@3388.4]
  wire [1:0] _T_2908; // @[Mux.scala 19:72:@3389.4]
  wire [1:0] _T_2909; // @[Mux.scala 19:72:@3390.4]
  wire [1:0] _T_2910; // @[Mux.scala 19:72:@3391.4]
  wire [1:0] _T_2911; // @[Mux.scala 19:72:@3392.4]
  wire [1:0] _T_2912; // @[Mux.scala 19:72:@3393.4]
  wire [1:0] _T_2913; // @[Mux.scala 19:72:@3394.4]
  wire [1:0] _T_2914; // @[Mux.scala 19:72:@3395.4]
  wire [1:0] _T_2915; // @[Mux.scala 19:72:@3396.4]
  wire [1:0] _T_2916; // @[Mux.scala 19:72:@3397.4]
  wire [1:0] _T_2917; // @[Mux.scala 19:72:@3398.4]
  wire [1:0] _T_2918; // @[Mux.scala 19:72:@3399.4]
  wire [1:0] _T_2919; // @[Mux.scala 19:72:@3400.4]
  wire [1:0] feedback_h_count; // @[Mux.scala 19:72:@3401.4]
  wire  _T_2925; // @[BTB.scala 186:30:@3407.4]
  wire [31:0] _T_2926; // @[OneHot.scala 26:18:@3408.4]
  wire [31:0] _T_2927; // @[OneHot.scala 27:18:@3409.4]
  wire  _T_2929; // @[OneHot.scala 28:14:@3410.4]
  wire [31:0] _T_2930; // @[OneHot.scala 28:28:@3411.4]
  wire [15:0] _T_2931; // @[OneHot.scala 26:18:@3412.4]
  wire [15:0] _T_2932; // @[OneHot.scala 27:18:@3413.4]
  wire  _T_2934; // @[OneHot.scala 28:14:@3414.4]
  wire [15:0] _T_2935; // @[OneHot.scala 28:28:@3415.4]
  wire [7:0] _T_2936; // @[OneHot.scala 26:18:@3416.4]
  wire [7:0] _T_2937; // @[OneHot.scala 27:18:@3417.4]
  wire  _T_2939; // @[OneHot.scala 28:14:@3418.4]
  wire [7:0] _T_2940; // @[OneHot.scala 28:28:@3419.4]
  wire [3:0] _T_2941; // @[OneHot.scala 26:18:@3420.4]
  wire [3:0] _T_2942; // @[OneHot.scala 27:18:@3421.4]
  wire  _T_2944; // @[OneHot.scala 28:14:@3422.4]
  wire [3:0] _T_2945; // @[OneHot.scala 28:28:@3423.4]
  wire [1:0] _T_2946; // @[OneHot.scala 26:18:@3424.4]
  wire [1:0] _T_2947; // @[OneHot.scala 27:18:@3425.4]
  wire  _T_2949; // @[OneHot.scala 28:14:@3426.4]
  wire [1:0] _T_2950; // @[OneHot.scala 28:28:@3427.4]
  wire  _T_2951; // @[CircuitMath.scala 30:8:@3428.4]
  wire [5:0] _T_2956; // @[Cat.scala 30:58:@3433.4]
  wire [63:0] _T_3020; // @[BTB.scala 196:26:@3497.4]
  wire  _T_3022; // @[BTB.scala 196:26:@3498.4]
  wire  _T_3087; // @[OneHot.scala 39:40:@3563.4]
  wire  _T_3088; // @[OneHot.scala 39:40:@3564.4]
  wire  _T_3089; // @[OneHot.scala 39:40:@3565.4]
  wire  _T_3090; // @[OneHot.scala 39:40:@3566.4]
  wire  _T_3091; // @[OneHot.scala 39:40:@3567.4]
  wire  _T_3092; // @[OneHot.scala 39:40:@3568.4]
  wire  _T_3093; // @[OneHot.scala 39:40:@3569.4]
  wire  _T_3094; // @[OneHot.scala 39:40:@3570.4]
  wire  _T_3095; // @[OneHot.scala 39:40:@3571.4]
  wire  _T_3096; // @[OneHot.scala 39:40:@3572.4]
  wire  _T_3097; // @[OneHot.scala 39:40:@3573.4]
  wire  _T_3098; // @[OneHot.scala 39:40:@3574.4]
  wire  _T_3099; // @[OneHot.scala 39:40:@3575.4]
  wire  _T_3100; // @[OneHot.scala 39:40:@3576.4]
  wire  _T_3101; // @[OneHot.scala 39:40:@3577.4]
  wire  _T_3102; // @[OneHot.scala 39:40:@3578.4]
  wire  _T_3103; // @[OneHot.scala 39:40:@3579.4]
  wire  _T_3104; // @[OneHot.scala 39:40:@3580.4]
  wire  _T_3105; // @[OneHot.scala 39:40:@3581.4]
  wire  _T_3106; // @[OneHot.scala 39:40:@3582.4]
  wire  _T_3107; // @[OneHot.scala 39:40:@3583.4]
  wire  _T_3108; // @[OneHot.scala 39:40:@3584.4]
  wire  _T_3109; // @[OneHot.scala 39:40:@3585.4]
  wire  _T_3110; // @[OneHot.scala 39:40:@3586.4]
  wire  _T_3111; // @[OneHot.scala 39:40:@3587.4]
  wire  _T_3112; // @[OneHot.scala 39:40:@3588.4]
  wire  _T_3113; // @[OneHot.scala 39:40:@3589.4]
  wire  _T_3114; // @[OneHot.scala 39:40:@3590.4]
  wire  _T_3115; // @[OneHot.scala 39:40:@3591.4]
  wire  _T_3116; // @[OneHot.scala 39:40:@3592.4]
  wire  _T_3117; // @[OneHot.scala 39:40:@3593.4]
  wire  _T_3118; // @[OneHot.scala 39:40:@3594.4]
  wire  _T_3119; // @[OneHot.scala 39:40:@3595.4]
  wire  _T_3120; // @[OneHot.scala 39:40:@3596.4]
  wire  _T_3121; // @[OneHot.scala 39:40:@3597.4]
  wire  _T_3122; // @[OneHot.scala 39:40:@3598.4]
  wire  _T_3123; // @[OneHot.scala 39:40:@3599.4]
  wire  _T_3124; // @[OneHot.scala 39:40:@3600.4]
  wire  _T_3125; // @[OneHot.scala 39:40:@3601.4]
  wire  _T_3126; // @[OneHot.scala 39:40:@3602.4]
  wire  _T_3127; // @[OneHot.scala 39:40:@3603.4]
  wire  _T_3128; // @[OneHot.scala 39:40:@3604.4]
  wire  _T_3129; // @[OneHot.scala 39:40:@3605.4]
  wire  _T_3130; // @[OneHot.scala 39:40:@3606.4]
  wire  _T_3131; // @[OneHot.scala 39:40:@3607.4]
  wire  _T_3132; // @[OneHot.scala 39:40:@3608.4]
  wire  _T_3133; // @[OneHot.scala 39:40:@3609.4]
  wire  _T_3134; // @[OneHot.scala 39:40:@3610.4]
  wire  _T_3135; // @[OneHot.scala 39:40:@3611.4]
  wire  _T_3136; // @[OneHot.scala 39:40:@3612.4]
  wire  _T_3137; // @[OneHot.scala 39:40:@3613.4]
  wire  _T_3138; // @[OneHot.scala 39:40:@3614.4]
  wire  _T_3139; // @[OneHot.scala 39:40:@3615.4]
  wire  _T_3140; // @[OneHot.scala 39:40:@3616.4]
  wire  _T_3141; // @[OneHot.scala 39:40:@3617.4]
  wire  _T_3142; // @[OneHot.scala 39:40:@3618.4]
  wire  _T_3143; // @[OneHot.scala 39:40:@3619.4]
  wire  _T_3144; // @[OneHot.scala 39:40:@3620.4]
  wire  _T_3145; // @[OneHot.scala 39:40:@3621.4]
  wire  _T_3146; // @[OneHot.scala 39:40:@3622.4]
  wire  _T_3147; // @[OneHot.scala 39:40:@3623.4]
  wire  _T_3148; // @[OneHot.scala 39:40:@3624.4]
  wire  _T_3149; // @[OneHot.scala 39:40:@3625.4]
  wire [5:0] _T_3215; // @[Mux.scala 31:69:@3627.4]
  wire [5:0] _T_3216; // @[Mux.scala 31:69:@3628.4]
  wire [5:0] _T_3217; // @[Mux.scala 31:69:@3629.4]
  wire [5:0] _T_3218; // @[Mux.scala 31:69:@3630.4]
  wire [5:0] _T_3219; // @[Mux.scala 31:69:@3631.4]
  wire [5:0] _T_3220; // @[Mux.scala 31:69:@3632.4]
  wire [5:0] _T_3221; // @[Mux.scala 31:69:@3633.4]
  wire [5:0] _T_3222; // @[Mux.scala 31:69:@3634.4]
  wire [5:0] _T_3223; // @[Mux.scala 31:69:@3635.4]
  wire [5:0] _T_3224; // @[Mux.scala 31:69:@3636.4]
  wire [5:0] _T_3225; // @[Mux.scala 31:69:@3637.4]
  wire [5:0] _T_3226; // @[Mux.scala 31:69:@3638.4]
  wire [5:0] _T_3227; // @[Mux.scala 31:69:@3639.4]
  wire [5:0] _T_3228; // @[Mux.scala 31:69:@3640.4]
  wire [5:0] _T_3229; // @[Mux.scala 31:69:@3641.4]
  wire [5:0] _T_3230; // @[Mux.scala 31:69:@3642.4]
  wire [5:0] _T_3231; // @[Mux.scala 31:69:@3643.4]
  wire [5:0] _T_3232; // @[Mux.scala 31:69:@3644.4]
  wire [5:0] _T_3233; // @[Mux.scala 31:69:@3645.4]
  wire [5:0] _T_3234; // @[Mux.scala 31:69:@3646.4]
  wire [5:0] _T_3235; // @[Mux.scala 31:69:@3647.4]
  wire [5:0] _T_3236; // @[Mux.scala 31:69:@3648.4]
  wire [5:0] _T_3237; // @[Mux.scala 31:69:@3649.4]
  wire [5:0] _T_3238; // @[Mux.scala 31:69:@3650.4]
  wire [5:0] _T_3239; // @[Mux.scala 31:69:@3651.4]
  wire [5:0] _T_3240; // @[Mux.scala 31:69:@3652.4]
  wire [5:0] _T_3241; // @[Mux.scala 31:69:@3653.4]
  wire [5:0] _T_3242; // @[Mux.scala 31:69:@3654.4]
  wire [5:0] _T_3243; // @[Mux.scala 31:69:@3655.4]
  wire [5:0] _T_3244; // @[Mux.scala 31:69:@3656.4]
  wire [5:0] _T_3245; // @[Mux.scala 31:69:@3657.4]
  wire [5:0] _T_3246; // @[Mux.scala 31:69:@3658.4]
  wire [5:0] _T_3247; // @[Mux.scala 31:69:@3659.4]
  wire [5:0] _T_3248; // @[Mux.scala 31:69:@3660.4]
  wire [5:0] _T_3249; // @[Mux.scala 31:69:@3661.4]
  wire [5:0] _T_3250; // @[Mux.scala 31:69:@3662.4]
  wire [5:0] _T_3251; // @[Mux.scala 31:69:@3663.4]
  wire [5:0] _T_3252; // @[Mux.scala 31:69:@3664.4]
  wire [5:0] _T_3253; // @[Mux.scala 31:69:@3665.4]
  wire [5:0] _T_3254; // @[Mux.scala 31:69:@3666.4]
  wire [5:0] _T_3255; // @[Mux.scala 31:69:@3667.4]
  wire [5:0] _T_3256; // @[Mux.scala 31:69:@3668.4]
  wire [5:0] _T_3257; // @[Mux.scala 31:69:@3669.4]
  wire [5:0] _T_3258; // @[Mux.scala 31:69:@3670.4]
  wire [5:0] _T_3259; // @[Mux.scala 31:69:@3671.4]
  wire [5:0] _T_3260; // @[Mux.scala 31:69:@3672.4]
  wire [5:0] _T_3261; // @[Mux.scala 31:69:@3673.4]
  wire [5:0] _T_3262; // @[Mux.scala 31:69:@3674.4]
  wire [5:0] _T_3263; // @[Mux.scala 31:69:@3675.4]
  wire [5:0] _T_3264; // @[Mux.scala 31:69:@3676.4]
  wire [5:0] _T_3265; // @[Mux.scala 31:69:@3677.4]
  wire [5:0] _T_3266; // @[Mux.scala 31:69:@3678.4]
  wire [5:0] _T_3267; // @[Mux.scala 31:69:@3679.4]
  wire [5:0] _T_3268; // @[Mux.scala 31:69:@3680.4]
  wire [5:0] _T_3269; // @[Mux.scala 31:69:@3681.4]
  wire [5:0] _T_3270; // @[Mux.scala 31:69:@3682.4]
  wire [5:0] _T_3271; // @[Mux.scala 31:69:@3683.4]
  wire [5:0] _T_3272; // @[Mux.scala 31:69:@3684.4]
  wire [5:0] _T_3273; // @[Mux.scala 31:69:@3685.4]
  wire [5:0] _T_3274; // @[Mux.scala 31:69:@3686.4]
  wire [5:0] _T_3275; // @[Mux.scala 31:69:@3687.4]
  wire [5:0] _T_3276; // @[Mux.scala 31:69:@3688.4]
  wire [5:0] _T_3277; // @[Mux.scala 31:69:@3689.4]
  wire [5:0] _T_3278; // @[BTB.scala 196:8:@3690.4]
  wire [5:0] feedback_idx; // @[BTB.scala 195:26:@3691.4]
  wire  _GEN_9; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_10; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_11; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_12; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_13; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_14; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_15; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_16; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_17; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_18; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_19; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_20; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_21; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_22; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_23; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_24; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_25; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_26; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_27; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_28; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_29; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_30; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_31; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_32; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_33; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_34; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_35; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_36; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_37; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_38; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_39; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_40; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_41; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_42; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_43; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_44; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_45; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_46; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_47; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_48; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_49; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_50; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_51; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_52; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_53; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_54; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_55; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_56; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_57; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_58; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_59; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_60; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_61; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_62; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_63; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_64; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_65; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_66; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_67; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_68; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_69; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_70; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_71; // @[BTB.scala 201:32:@3697.8]
  wire  _GEN_72; // @[BTB.scala 201:32:@3697.8]
  wire  _T_3285; // @[BTB.scala 203:51:@3702.10]
  wire  _GEN_73; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_74; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_75; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_76; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_77; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_78; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_79; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_80; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_81; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_82; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_83; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_84; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_85; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_86; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_87; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_88; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_89; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_90; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_91; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_92; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_93; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_94; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_95; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_96; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_97; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_98; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_99; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_100; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_101; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_102; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_103; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_104; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_105; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_106; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_107; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_108; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_109; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_110; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_111; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_112; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_113; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_114; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_115; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_116; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_117; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_118; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_119; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_120; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_121; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_122; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_123; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_124; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_125; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_126; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_127; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_128; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_129; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_130; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_131; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_132; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_133; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_134; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_135; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_136; // @[BTB.scala 203:32:@3703.10]
  wire  _GEN_137; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_138; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_139; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_140; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_141; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_142; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_143; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_144; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_145; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_146; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_147; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_148; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_149; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_150; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_151; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_152; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_153; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_154; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_155; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_156; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_157; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_158; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_159; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_160; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_161; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_162; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_163; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_164; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_165; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_166; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_167; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_168; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_169; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_170; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_171; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_172; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_173; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_174; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_175; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_176; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_177; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_178; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_179; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_180; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_181; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_182; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_183; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_184; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_185; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_186; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_187; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_188; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_189; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_190; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_191; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_192; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_193; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_194; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_195; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_196; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_197; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_198; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_199; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_200; // @[BTB.scala 202:32:@3701.8]
  wire  _GEN_201; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_202; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_203; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_204; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_205; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_206; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_207; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_208; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_209; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_210; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_211; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_212; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_213; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_214; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_215; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_216; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_217; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_218; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_219; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_220; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_221; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_222; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_223; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_224; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_225; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_226; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_227; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_228; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_229; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_230; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_231; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_232; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_233; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_234; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_235; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_236; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_237; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_238; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_239; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_240; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_241; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_242; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_243; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_244; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_245; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_246; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_247; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_248; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_249; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_250; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_251; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_252; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_253; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_254; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_255; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_256; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_257; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_258; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_259; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_260; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_261; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_262; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_263; // @[BTB.scala 200:28:@3696.6]
  wire  _GEN_264; // @[BTB.scala 200:28:@3696.6]
  wire [29:0] _GEN_265; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_266; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_267; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_268; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_269; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_270; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_271; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_272; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_273; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_274; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_275; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_276; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_277; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_278; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_279; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_280; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_281; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_282; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_283; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_284; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_285; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_286; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_287; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_288; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_289; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_290; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_291; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_292; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_293; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_294; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_295; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_296; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_297; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_298; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_299; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_300; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_301; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_302; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_303; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_304; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_305; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_306; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_307; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_308; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_309; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_310; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_311; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_312; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_313; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_314; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_315; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_316; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_317; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_318; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_319; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_320; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_321; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_322; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_323; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_324; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_325; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_326; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_327; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_328; // @[BTB.scala 206:33:@3706.8]
  wire [29:0] _GEN_329; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_330; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_331; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_332; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_333; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_334; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_335; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_336; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_337; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_338; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_339; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_340; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_341; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_342; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_343; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_344; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_345; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_346; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_347; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_348; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_349; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_350; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_351; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_352; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_353; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_354; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_355; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_356; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_357; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_358; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_359; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_360; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_361; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_362; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_363; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_364; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_365; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_366; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_367; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_368; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_369; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_370; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_371; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_372; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_373; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_374; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_375; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_376; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_377; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_378; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_379; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_380; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_381; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_382; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_383; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_384; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_385; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_386; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_387; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_388; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_389; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_390; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_391; // @[BTB.scala 207:33:@3707.8]
  wire [29:0] _GEN_392; // @[BTB.scala 207:33:@3707.8]
  wire [1:0] _GEN_393; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_394; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_395; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_396; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_397; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_398; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_399; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_400; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_401; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_402; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_403; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_404; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_405; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_406; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_407; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_408; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_409; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_410; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_411; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_412; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_413; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_414; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_415; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_416; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_417; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_418; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_419; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_420; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_421; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_422; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_423; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_424; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_425; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_426; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_427; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_428; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_429; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_430; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_431; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_432; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_433; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_434; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_435; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_436; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_437; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_438; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_439; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_440; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_441; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_442; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_443; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_444; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_445; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_446; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_447; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_448; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_449; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_450; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_451; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_452; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_453; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_454; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_455; // @[BTB.scala 208:33:@3708.8]
  wire [1:0] _GEN_456; // @[BTB.scala 208:33:@3708.8]
  wire [29:0] _GEN_457; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_458; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_459; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_460; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_461; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_462; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_463; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_464; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_465; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_466; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_467; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_468; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_469; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_470; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_471; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_472; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_473; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_474; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_475; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_476; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_477; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_478; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_479; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_480; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_481; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_482; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_483; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_484; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_485; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_486; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_487; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_488; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_489; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_490; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_491; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_492; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_493; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_494; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_495; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_496; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_497; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_498; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_499; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_500; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_501; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_502; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_503; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_504; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_505; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_506; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_507; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_508; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_509; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_510; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_511; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_512; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_513; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_514; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_515; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_516; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_517; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_518; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_519; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_520; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_521; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_522; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_523; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_524; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_525; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_526; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_527; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_528; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_529; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_530; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_531; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_532; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_533; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_534; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_535; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_536; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_537; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_538; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_539; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_540; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_541; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_542; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_543; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_544; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_545; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_546; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_547; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_548; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_549; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_550; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_551; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_552; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_553; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_554; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_555; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_556; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_557; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_558; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_559; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_560; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_561; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_562; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_563; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_564; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_565; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_566; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_567; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_568; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_569; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_570; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_571; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_572; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_573; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_574; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_575; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_576; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_577; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_578; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_579; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_580; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_581; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_582; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_583; // @[BTB.scala 205:28:@3705.6]
  wire [29:0] _GEN_584; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_585; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_586; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_587; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_588; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_589; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_590; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_591; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_592; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_593; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_594; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_595; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_596; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_597; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_598; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_599; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_600; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_601; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_602; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_603; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_604; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_605; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_606; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_607; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_608; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_609; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_610; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_611; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_612; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_613; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_614; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_615; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_616; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_617; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_618; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_619; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_620; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_621; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_622; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_623; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_624; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_625; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_626; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_627; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_628; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_629; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_630; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_631; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_632; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_633; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_634; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_635; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_636; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_637; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_638; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_639; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_640; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_641; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_642; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_643; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_644; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_645; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_646; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_647; // @[BTB.scala 205:28:@3705.6]
  wire [1:0] _GEN_648; // @[BTB.scala 205:28:@3705.6]
  wire  _T_3291; // @[BTB.scala 72:38:@3715.12]
  wire  _T_3292; // @[BTB.scala 72:45:@3716.12]
  wire  _T_3293; // @[BTB.scala 72:54:@3717.12]
  wire  _T_3295; // @[BTB.scala 72:52:@3718.12]
  wire  _T_3296; // @[BTB.scala 72:49:@3719.12]
  wire [1:0] _T_3297; // @[Cat.scala 30:58:@3720.12]
  wire [1:0] _GEN_649; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_650; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_651; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_652; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_653; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_654; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_655; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_656; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_657; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_658; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_659; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_660; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_661; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_662; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_663; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_664; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_665; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_666; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_667; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_668; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_669; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_670; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_671; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_672; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_673; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_674; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_675; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_676; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_677; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_678; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_679; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_680; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_681; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_682; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_683; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_684; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_685; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_686; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_687; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_688; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_689; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_690; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_691; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_692; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_693; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_694; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_695; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_696; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_697; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_698; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_699; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_700; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_701; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_702; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_703; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_704; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_705; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_706; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_707; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_708; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_709; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_710; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_711; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] _GEN_712; // @[BTB.scala 214:37:@3721.12]
  wire [1:0] feedback_gshare; // @[BTB.scala 184:22:@2953.4 BTB.scala 194:20:@3406.4]
  wire  _T_3300; // @[BTB.scala 72:38:@3723.12]
  wire  _T_3301; // @[BTB.scala 72:45:@3724.12]
  wire  _T_3302; // @[BTB.scala 72:54:@3725.12]
  wire  _T_3304; // @[BTB.scala 72:52:@3726.12]
  wire  _T_3305; // @[BTB.scala 72:49:@3727.12]
  wire [1:0] _T_3307; // @[BTB.scala 74:38:@3732.12]
  wire  _T_3309; // @[BTB.scala 74:38:@3733.12]
  wire  _T_3314; // @[BTB.scala 74:49:@3737.12]
  wire [1:0] _T_3315; // @[Cat.scala 30:58:@3738.12]
  wire [1:0] _GEN_713; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_714; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_715; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_716; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_717; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_718; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_719; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_720; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_721; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_722; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_723; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_724; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_725; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_726; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_727; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_728; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_729; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_730; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_731; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_732; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_733; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_734; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_735; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_736; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_737; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_738; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_739; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_740; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_741; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_742; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_743; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_744; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_745; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_746; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_747; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_748; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_749; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_750; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_751; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_752; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_753; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_754; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_755; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_756; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_757; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_758; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_759; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_760; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_761; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_762; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_763; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_764; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_765; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_766; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_767; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_768; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_769; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_770; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_771; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_772; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_773; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_774; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_775; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _GEN_776; // @[BTB.scala 217:37:@3739.12]
  wire [1:0] _T_3317; // @[BTB.scala 74:38:@3741.12]
  wire  _T_3319; // @[BTB.scala 74:38:@3742.12]
  wire  _T_3324; // @[BTB.scala 74:49:@3746.12]
  wire [1:0] _GEN_777; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_778; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_779; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_780; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_781; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_782; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_783; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_784; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_785; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_786; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_787; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_788; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_789; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_790; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_791; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_792; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_793; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_794; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_795; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_796; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_797; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_798; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_799; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_800; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_801; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_802; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_803; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_804; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_805; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_806; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_807; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_808; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_809; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_810; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_811; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_812; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_813; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_814; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_815; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_816; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_817; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_818; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_819; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_820; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_821; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_822; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_823; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_824; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_825; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_826; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_827; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_828; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_829; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_830; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_831; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_832; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_833; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_834; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_835; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_836; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_837; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_838; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_839; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_840; // @[BTB.scala 213:32:@3714.10]
  wire  _GEN_848; // @[BTB.scala 213:32:@3714.10]
  wire [1:0] _GEN_851; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_852; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_853; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_854; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_855; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_856; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_857; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_858; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_859; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_860; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_861; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_862; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_863; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_864; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_865; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_866; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_867; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_868; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_869; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_870; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_871; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_872; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_873; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_874; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_875; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_876; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_877; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_878; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_879; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_880; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_881; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_882; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_883; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_884; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_885; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_886; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_887; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_888; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_889; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_890; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_891; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_892; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_893; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_894; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_895; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_896; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_897; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_898; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_899; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_900; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_901; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_902; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_903; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_904; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_905; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_906; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_907; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_908; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_909; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_910; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_911; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_912; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_913; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_914; // @[BTB.scala 221:35:@3753.12]
  wire [1:0] _GEN_915; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_916; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_917; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_918; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_919; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_920; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_921; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_922; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_923; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_924; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_925; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_926; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_927; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_928; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_929; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_930; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_931; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_932; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_933; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_934; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_935; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_936; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_937; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_938; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_939; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_940; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_941; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_942; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_943; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_944; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_945; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_946; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_947; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_948; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_949; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_950; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_951; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_952; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_953; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_954; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_955; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_956; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_957; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_958; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_959; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_960; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_961; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_962; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_963; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_964; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_965; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_966; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_967; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_968; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_969; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_970; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_971; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_972; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_973; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_974; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_975; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_976; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_977; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_978; // @[BTB.scala 220:35:@3752.10]
  wire [1:0] _GEN_980; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_981; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_982; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_983; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_984; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_985; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_986; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_987; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_988; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_989; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_990; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_991; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_992; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_993; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_994; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_995; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_996; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_997; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_998; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_999; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1000; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1001; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1002; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1003; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1004; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1005; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1006; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1007; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1008; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1009; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1010; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1011; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1012; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1013; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1014; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1015; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1016; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1017; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1018; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1019; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1020; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1021; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1022; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1023; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1024; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1025; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1026; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1027; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1028; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1029; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1030; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1031; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1032; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1033; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1034; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1035; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1036; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1037; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1038; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1039; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1040; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1041; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1042; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1043; // @[BTB.scala 212:29:@3713.8]
  wire  _GEN_1046; // @[BTB.scala 212:29:@3713.8]
  wire  _GEN_1051; // @[BTB.scala 212:29:@3713.8]
  wire  _GEN_1056; // @[BTB.scala 212:29:@3713.8]
  wire [1:0] _GEN_1059; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1060; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1061; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1062; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1063; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1064; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1065; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1066; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1067; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1068; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1069; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1070; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1071; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1072; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1073; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1074; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1075; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1076; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1077; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1078; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1079; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1080; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1081; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1082; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1083; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1084; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1085; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1086; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1087; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1088; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1089; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1090; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1091; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1092; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1093; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1094; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1095; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1096; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1097; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1098; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1099; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1100; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1101; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1102; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1103; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1104; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1105; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1106; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1107; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1108; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1109; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1110; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1111; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1112; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1113; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1114; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1115; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1116; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1117; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1118; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1119; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1120; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1121; // @[BTB.scala 211:49:@3711.6]
  wire [1:0] _GEN_1122; // @[BTB.scala 211:49:@3711.6]
  wire  _GEN_1125; // @[BTB.scala 211:49:@3711.6]
  wire  _GEN_1130; // @[BTB.scala 211:49:@3711.6]
  wire  _GEN_1135; // @[BTB.scala 211:49:@3711.6]
  wire  _GEN_1138; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1139; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1140; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1141; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1142; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1143; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1144; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1145; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1146; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1147; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1148; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1149; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1150; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1151; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1152; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1153; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1154; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1155; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1156; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1157; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1158; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1159; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1160; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1161; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1162; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1163; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1164; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1165; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1166; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1167; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1168; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1169; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1170; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1171; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1172; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1173; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1174; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1175; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1176; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1177; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1178; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1179; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1180; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1181; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1182; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1183; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1184; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1185; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1186; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1187; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1188; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1189; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1190; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1191; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1192; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1193; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1194; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1195; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1196; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1197; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1198; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1199; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1200; // @[BTB.scala 199:23:@3695.4]
  wire  _GEN_1201; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1202; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1203; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1204; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1205; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1206; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1207; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1208; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1209; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1210; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1211; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1212; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1213; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1214; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1215; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1216; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1217; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1218; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1219; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1220; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1221; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1222; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1223; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1224; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1225; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1226; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1227; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1228; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1229; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1230; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1231; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1232; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1233; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1234; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1235; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1236; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1237; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1238; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1239; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1240; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1241; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1242; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1243; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1244; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1245; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1246; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1247; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1248; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1249; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1250; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1251; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1252; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1253; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1254; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1255; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1256; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1257; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1258; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1259; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1260; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1261; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1262; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1263; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1264; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1265; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1266; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1267; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1268; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1269; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1270; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1271; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1272; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1273; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1274; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1275; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1276; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1277; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1278; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1279; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1280; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1281; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1282; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1283; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1284; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1285; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1286; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1287; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1288; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1289; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1290; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1291; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1292; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1293; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1294; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1295; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1296; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1297; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1298; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1299; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1300; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1301; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1302; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1303; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1304; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1305; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1306; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1307; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1308; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1309; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1310; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1311; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1312; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1313; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1314; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1315; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1316; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1317; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1318; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1319; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1320; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1321; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1322; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1323; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1324; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1325; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1326; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1327; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1328; // @[BTB.scala 199:23:@3695.4]
  wire [29:0] _GEN_1329; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1330; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1331; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1332; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1333; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1334; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1335; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1336; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1337; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1338; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1339; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1340; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1341; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1342; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1343; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1344; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1345; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1346; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1347; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1348; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1349; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1350; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1351; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1352; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1353; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1354; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1355; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1356; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1357; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1358; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1359; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1360; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1361; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1362; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1363; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1364; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1365; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1366; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1367; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1368; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1369; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1370; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1371; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1372; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1373; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1374; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1375; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1376; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1377; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1378; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1379; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1380; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1381; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1382; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1383; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1384; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1385; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1386; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1387; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1388; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1389; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1390; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1391; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1392; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1393; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1394; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1395; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1396; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1397; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1398; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1399; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1400; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1401; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1402; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1403; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1404; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1405; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1406; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1407; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1408; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1409; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1410; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1411; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1412; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1413; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1414; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1415; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1416; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1417; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1418; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1419; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1420; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1421; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1422; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1423; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1424; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1425; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1426; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1427; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1428; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1429; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1430; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1431; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1432; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1433; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1434; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1435; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1436; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1437; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1438; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1439; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1440; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1441; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1442; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1443; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1444; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1445; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1446; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1447; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1448; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1449; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1450; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1451; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1452; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1453; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1454; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1455; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1456; // @[BTB.scala 199:23:@3695.4]
  wire [1:0] _GEN_1457; // @[BTB.scala 199:23:@3695.4]
  wire  _T_3331; // @[BTB.scala 227:21:@3760.4]
  wire  feedback_select; // @[BTB.scala 184:22:@2953.4 BTB.scala 197:20:@3694.4]
  wire  _T_3333; // @[BTB.scala 228:26:@3762.6]
  wire  _T_3334; // @[BTB.scala 228:23:@3763.6]
  wire  _GEN_1479; // @[BTB.scala 228:44:@3764.6]
  wire [31:0] _T_3342; // @[Cat.scala 30:58:@3775.6]
  wire [31:0] _T_3352; // @[OneHot.scala 26:18:@3783.6]
  wire [31:0] _T_3353; // @[OneHot.scala 27:18:@3784.6]
  wire  _T_3355; // @[OneHot.scala 28:14:@3785.6]
  wire [31:0] _T_3356; // @[OneHot.scala 28:28:@3786.6]
  wire [15:0] _T_3357; // @[OneHot.scala 26:18:@3787.6]
  wire [15:0] _T_3358; // @[OneHot.scala 27:18:@3788.6]
  wire  _T_3360; // @[OneHot.scala 28:14:@3789.6]
  wire [15:0] _T_3361; // @[OneHot.scala 28:28:@3790.6]
  wire [7:0] _T_3362; // @[OneHot.scala 26:18:@3791.6]
  wire [7:0] _T_3363; // @[OneHot.scala 27:18:@3792.6]
  wire  _T_3365; // @[OneHot.scala 28:14:@3793.6]
  wire [7:0] _T_3366; // @[OneHot.scala 28:28:@3794.6]
  wire [3:0] _T_3367; // @[OneHot.scala 26:18:@3795.6]
  wire [3:0] _T_3368; // @[OneHot.scala 27:18:@3796.6]
  wire  _T_3370; // @[OneHot.scala 28:14:@3797.6]
  wire [3:0] _T_3371; // @[OneHot.scala 28:28:@3798.6]
  wire [1:0] _T_3372; // @[OneHot.scala 26:18:@3799.6]
  wire [1:0] _T_3373; // @[OneHot.scala 27:18:@3800.6]
  wire  _T_3375; // @[OneHot.scala 28:14:@3801.6]
  wire [1:0] _T_3376; // @[OneHot.scala 28:28:@3802.6]
  wire  _T_3377; // @[CircuitMath.scala 30:8:@3803.6]
  wire [5:0] _T_3382; // @[Cat.scala 30:58:@3808.6]
  wire  _T_3385; // @[BTB.scala 237:13:@3810.6]
  wire  _T_3386; // @[BTB.scala 248:50:@3814.6]
  wire  _T_3390; // @[BTB.scala 248:50:@3820.6]
  wire  _T_3394; // @[BTB.scala 248:50:@3826.6]
  wire  _T_3398; // @[BTB.scala 248:50:@3832.6]
  wire  _T_3402; // @[BTB.scala 248:50:@3838.6]
  wire  _T_3406; // @[BTB.scala 248:50:@3844.6]
  wire  _T_3410; // @[BTB.scala 248:50:@3850.6]
  wire  _T_3414; // @[BTB.scala 248:50:@3856.6]
  wire  _T_3418; // @[BTB.scala 248:50:@3862.6]
  wire  _T_3422; // @[BTB.scala 249:28:@3868.6]
  wire [31:0] _T_3439; // @[OneHot.scala 26:18:@3885.6]
  wire [31:0] _T_3440; // @[OneHot.scala 27:18:@3886.6]
  wire  _T_3442; // @[OneHot.scala 28:14:@3887.6]
  wire [31:0] _T_3443; // @[OneHot.scala 28:28:@3888.6]
  wire [15:0] _T_3444; // @[OneHot.scala 26:18:@3889.6]
  wire [15:0] _T_3445; // @[OneHot.scala 27:18:@3890.6]
  wire  _T_3447; // @[OneHot.scala 28:14:@3891.6]
  wire [15:0] _T_3448; // @[OneHot.scala 28:28:@3892.6]
  wire [7:0] _T_3449; // @[OneHot.scala 26:18:@3893.6]
  wire [7:0] _T_3450; // @[OneHot.scala 27:18:@3894.6]
  wire  _T_3452; // @[OneHot.scala 28:14:@3895.6]
  wire [7:0] _T_3453; // @[OneHot.scala 28:28:@3896.6]
  wire [3:0] _T_3454; // @[OneHot.scala 26:18:@3897.6]
  wire [3:0] _T_3455; // @[OneHot.scala 27:18:@3898.6]
  wire  _T_3457; // @[OneHot.scala 28:14:@3899.6]
  wire [3:0] _T_3458; // @[OneHot.scala 28:28:@3900.6]
  wire [1:0] _T_3459; // @[OneHot.scala 26:18:@3901.6]
  wire [1:0] _T_3460; // @[OneHot.scala 27:18:@3902.6]
  wire  _T_3462; // @[OneHot.scala 28:14:@3903.6]
  wire [1:0] _T_3463; // @[OneHot.scala 28:28:@3904.6]
  wire  _T_3464; // @[CircuitMath.scala 30:8:@3905.6]
  wire [5:0] _T_3469; // @[Cat.scala 30:58:@3910.6]
  RAS RAS ( // @[BTB.scala 79:19:@759.4]
    .clock(RAS_clock),
    .reset(RAS_reset),
    .io_push_valid(RAS_io_push_valid),
    .io_push_bits(RAS_io_push_bits),
    .io_pop(RAS_io_pop),
    .io_peek(RAS_io_peek)
  );
  assign bht__T_1239_addr = gb_history ^ _T_1236;
  assign bht__T_1239_data = bht[bht__T_1239_addr]; // @[BTB.scala 77:16:@757.4]
  assign bht__T_2316_addr = gb_history ^ _T_2313;
  assign bht__T_2316_data = bht[bht__T_2316_addr]; // @[BTB.scala 77:16:@757.4]
  assign bht__T_2923_addr = fb_reg_gshxor;
  assign bht__T_2923_data = bht[bht__T_2923_addr]; // @[BTB.scala 77:16:@757.4]
  assign bht__T_3298_data = {_T_3300,_T_3305};
  assign bht__T_3298_addr = fb_reg_gshxor;
  assign bht__T_3298_mask = 1'h1;
  assign bht__T_3298_en = fb_reg_valid ? _GEN_1125 : 1'h0;
  assign bht__T_3316_data = {_T_3319,_T_3324};
  assign bht__T_3316_addr = fb_reg_gshxor;
  assign bht__T_3316_mask = 1'h1;
  assign bht__T_3316_en = fb_reg_valid ? _GEN_1130 : 1'h0;
  assign bht__T_3327_data = 2'h2;
  assign bht__T_3327_addr = fb_reg_gshxor;
  assign bht__T_3327_mask = 1'h1;
  assign bht__T_3327_en = fb_reg_valid ? _GEN_1135 : 1'h0;
  assign arb__T_1238_addr = gb_history ^ _T_1236;
  assign arb__T_1238_data = arb[arb__T_1238_addr]; // @[BTB.scala 78:16:@758.4]
  assign arb__T_2315_addr = gb_history ^ _T_2313;
  assign arb__T_2315_data = arb[arb__T_2315_addr]; // @[BTB.scala 78:16:@758.4]
  assign arb__T_3280_addr = fb_reg_gshxor;
  assign arb__T_3280_data = arb[arb__T_3280_addr]; // @[BTB.scala 78:16:@758.4]
  assign arb__T_3335_data = 1'h1;
  assign arb__T_3335_addr = fb_reg_gshxor;
  assign arb__T_3335_mask = 1'h1;
  assign arb__T_3335_en = _T_3331 ? _T_3334 : 1'h0;
  assign arb__T_3337_data = 1'h0;
  assign arb__T_3337_addr = fb_reg_gshxor;
  assign arb__T_3337_mask = 1'h1;
  assign arb__T_3337_en = _T_3331 ? _GEN_1479 : 1'h0;
  assign _T_175 = io_if_pc_bits[31:3]; // @[BTB.scala 99:43:@1088.4]
  assign _T_178 = {_T_175,1'h1}; // @[Cat.scala 30:58:@1089.4]
  assign predict_0_cont_tgt = {_T_175,1'h1,2'h0}; // @[Cat.scala 30:58:@1090.4]
  assign _T_181 = predict_0_cont_tgt + 32'h4; // @[BTB.scala 100:46:@1092.4]
  assign predict_1_cont_tgt = predict_0_cont_tgt + 32'h4; // @[BTB.scala 100:46:@1093.4]
  assign _T_183 = io_if_pc_bits[2]; // @[BTB.scala 101:55:@1095.4]
  assign _T_186 = _T_183 == 1'h0; // @[BTB.scala 101:41:@1097.4]
  assign if_pc_0 = {_T_175,1'h0}; // @[Cat.scala 30:58:@1102.4]
  assign _T_198 = btb_pc_0 == if_pc_0; // @[BTB.scala 105:47:@1104.4]
  assign _T_199 = btb_pc_1 == if_pc_0; // @[BTB.scala 105:47:@1105.4]
  assign _T_200 = btb_pc_2 == if_pc_0; // @[BTB.scala 105:47:@1106.4]
  assign _T_201 = btb_pc_3 == if_pc_0; // @[BTB.scala 105:47:@1107.4]
  assign _T_202 = btb_pc_4 == if_pc_0; // @[BTB.scala 105:47:@1108.4]
  assign _T_203 = btb_pc_5 == if_pc_0; // @[BTB.scala 105:47:@1109.4]
  assign _T_204 = btb_pc_6 == if_pc_0; // @[BTB.scala 105:47:@1110.4]
  assign _T_205 = btb_pc_7 == if_pc_0; // @[BTB.scala 105:47:@1111.4]
  assign _T_206 = btb_pc_8 == if_pc_0; // @[BTB.scala 105:47:@1112.4]
  assign _T_207 = btb_pc_9 == if_pc_0; // @[BTB.scala 105:47:@1113.4]
  assign _T_208 = btb_pc_10 == if_pc_0; // @[BTB.scala 105:47:@1114.4]
  assign _T_209 = btb_pc_11 == if_pc_0; // @[BTB.scala 105:47:@1115.4]
  assign _T_210 = btb_pc_12 == if_pc_0; // @[BTB.scala 105:47:@1116.4]
  assign _T_211 = btb_pc_13 == if_pc_0; // @[BTB.scala 105:47:@1117.4]
  assign _T_212 = btb_pc_14 == if_pc_0; // @[BTB.scala 105:47:@1118.4]
  assign _T_213 = btb_pc_15 == if_pc_0; // @[BTB.scala 105:47:@1119.4]
  assign _T_214 = btb_pc_16 == if_pc_0; // @[BTB.scala 105:47:@1120.4]
  assign _T_215 = btb_pc_17 == if_pc_0; // @[BTB.scala 105:47:@1121.4]
  assign _T_216 = btb_pc_18 == if_pc_0; // @[BTB.scala 105:47:@1122.4]
  assign _T_217 = btb_pc_19 == if_pc_0; // @[BTB.scala 105:47:@1123.4]
  assign _T_218 = btb_pc_20 == if_pc_0; // @[BTB.scala 105:47:@1124.4]
  assign _T_219 = btb_pc_21 == if_pc_0; // @[BTB.scala 105:47:@1125.4]
  assign _T_220 = btb_pc_22 == if_pc_0; // @[BTB.scala 105:47:@1126.4]
  assign _T_221 = btb_pc_23 == if_pc_0; // @[BTB.scala 105:47:@1127.4]
  assign _T_222 = btb_pc_24 == if_pc_0; // @[BTB.scala 105:47:@1128.4]
  assign _T_223 = btb_pc_25 == if_pc_0; // @[BTB.scala 105:47:@1129.4]
  assign _T_224 = btb_pc_26 == if_pc_0; // @[BTB.scala 105:47:@1130.4]
  assign _T_225 = btb_pc_27 == if_pc_0; // @[BTB.scala 105:47:@1131.4]
  assign _T_226 = btb_pc_28 == if_pc_0; // @[BTB.scala 105:47:@1132.4]
  assign _T_227 = btb_pc_29 == if_pc_0; // @[BTB.scala 105:47:@1133.4]
  assign _T_228 = btb_pc_30 == if_pc_0; // @[BTB.scala 105:47:@1134.4]
  assign _T_229 = btb_pc_31 == if_pc_0; // @[BTB.scala 105:47:@1135.4]
  assign _T_230 = btb_pc_32 == if_pc_0; // @[BTB.scala 105:47:@1136.4]
  assign _T_231 = btb_pc_33 == if_pc_0; // @[BTB.scala 105:47:@1137.4]
  assign _T_232 = btb_pc_34 == if_pc_0; // @[BTB.scala 105:47:@1138.4]
  assign _T_233 = btb_pc_35 == if_pc_0; // @[BTB.scala 105:47:@1139.4]
  assign _T_234 = btb_pc_36 == if_pc_0; // @[BTB.scala 105:47:@1140.4]
  assign _T_235 = btb_pc_37 == if_pc_0; // @[BTB.scala 105:47:@1141.4]
  assign _T_236 = btb_pc_38 == if_pc_0; // @[BTB.scala 105:47:@1142.4]
  assign _T_237 = btb_pc_39 == if_pc_0; // @[BTB.scala 105:47:@1143.4]
  assign _T_238 = btb_pc_40 == if_pc_0; // @[BTB.scala 105:47:@1144.4]
  assign _T_239 = btb_pc_41 == if_pc_0; // @[BTB.scala 105:47:@1145.4]
  assign _T_240 = btb_pc_42 == if_pc_0; // @[BTB.scala 105:47:@1146.4]
  assign _T_241 = btb_pc_43 == if_pc_0; // @[BTB.scala 105:47:@1147.4]
  assign _T_242 = btb_pc_44 == if_pc_0; // @[BTB.scala 105:47:@1148.4]
  assign _T_243 = btb_pc_45 == if_pc_0; // @[BTB.scala 105:47:@1149.4]
  assign _T_244 = btb_pc_46 == if_pc_0; // @[BTB.scala 105:47:@1150.4]
  assign _T_245 = btb_pc_47 == if_pc_0; // @[BTB.scala 105:47:@1151.4]
  assign _T_246 = btb_pc_48 == if_pc_0; // @[BTB.scala 105:47:@1152.4]
  assign _T_247 = btb_pc_49 == if_pc_0; // @[BTB.scala 105:47:@1153.4]
  assign _T_248 = btb_pc_50 == if_pc_0; // @[BTB.scala 105:47:@1154.4]
  assign _T_249 = btb_pc_51 == if_pc_0; // @[BTB.scala 105:47:@1155.4]
  assign _T_250 = btb_pc_52 == if_pc_0; // @[BTB.scala 105:47:@1156.4]
  assign _T_251 = btb_pc_53 == if_pc_0; // @[BTB.scala 105:47:@1157.4]
  assign _T_252 = btb_pc_54 == if_pc_0; // @[BTB.scala 105:47:@1158.4]
  assign _T_253 = btb_pc_55 == if_pc_0; // @[BTB.scala 105:47:@1159.4]
  assign _T_254 = btb_pc_56 == if_pc_0; // @[BTB.scala 105:47:@1160.4]
  assign _T_255 = btb_pc_57 == if_pc_0; // @[BTB.scala 105:47:@1161.4]
  assign _T_256 = btb_pc_58 == if_pc_0; // @[BTB.scala 105:47:@1162.4]
  assign _T_257 = btb_pc_59 == if_pc_0; // @[BTB.scala 105:47:@1163.4]
  assign _T_258 = btb_pc_60 == if_pc_0; // @[BTB.scala 105:47:@1164.4]
  assign _T_259 = btb_pc_61 == if_pc_0; // @[BTB.scala 105:47:@1165.4]
  assign _T_260 = btb_pc_62 == if_pc_0; // @[BTB.scala 105:47:@1166.4]
  assign _T_261 = btb_pc_63 == if_pc_0; // @[BTB.scala 105:47:@1167.4]
  assign _T_338 = {_T_205,_T_204,_T_203,_T_202,_T_201,_T_200,_T_199,_T_198}; // @[BTB.scala 105:62:@1239.4]
  assign _T_346 = {_T_213,_T_212,_T_211,_T_210,_T_209,_T_208,_T_207,_T_206,_T_338}; // @[BTB.scala 105:62:@1247.4]
  assign _T_353 = {_T_221,_T_220,_T_219,_T_218,_T_217,_T_216,_T_215,_T_214}; // @[BTB.scala 105:62:@1254.4]
  assign _T_362 = {_T_229,_T_228,_T_227,_T_226,_T_225,_T_224,_T_223,_T_222,_T_353,_T_346}; // @[BTB.scala 105:62:@1263.4]
  assign _T_369 = {_T_237,_T_236,_T_235,_T_234,_T_233,_T_232,_T_231,_T_230}; // @[BTB.scala 105:62:@1270.4]
  assign _T_377 = {_T_245,_T_244,_T_243,_T_242,_T_241,_T_240,_T_239,_T_238,_T_369}; // @[BTB.scala 105:62:@1278.4]
  assign _T_384 = {_T_253,_T_252,_T_251,_T_250,_T_249,_T_248,_T_247,_T_246}; // @[BTB.scala 105:62:@1285.4]
  assign _T_393 = {_T_261,_T_260,_T_259,_T_258,_T_257,_T_256,_T_255,_T_254,_T_384,_T_377}; // @[BTB.scala 105:62:@1294.4]
  assign _T_394 = {_T_393,_T_362}; // @[BTB.scala 105:62:@1295.4]
  assign _T_401 = {btb_valid_7,btb_valid_6,btb_valid_5,btb_valid_4,btb_valid_3,btb_valid_2,btb_valid_1,btb_valid_0}; // @[BTB.scala 105:81:@1302.4]
  assign _T_409 = {btb_valid_15,btb_valid_14,btb_valid_13,btb_valid_12,btb_valid_11,btb_valid_10,btb_valid_9,btb_valid_8,_T_401}; // @[BTB.scala 105:81:@1310.4]
  assign _T_416 = {btb_valid_23,btb_valid_22,btb_valid_21,btb_valid_20,btb_valid_19,btb_valid_18,btb_valid_17,btb_valid_16}; // @[BTB.scala 105:81:@1317.4]
  assign _T_425 = {btb_valid_31,btb_valid_30,btb_valid_29,btb_valid_28,btb_valid_27,btb_valid_26,btb_valid_25,btb_valid_24,_T_416,_T_409}; // @[BTB.scala 105:81:@1326.4]
  assign _T_432 = {btb_valid_39,btb_valid_38,btb_valid_37,btb_valid_36,btb_valid_35,btb_valid_34,btb_valid_33,btb_valid_32}; // @[BTB.scala 105:81:@1333.4]
  assign _T_440 = {btb_valid_47,btb_valid_46,btb_valid_45,btb_valid_44,btb_valid_43,btb_valid_42,btb_valid_41,btb_valid_40,_T_432}; // @[BTB.scala 105:81:@1341.4]
  assign _T_447 = {btb_valid_55,btb_valid_54,btb_valid_53,btb_valid_52,btb_valid_51,btb_valid_50,btb_valid_49,btb_valid_48}; // @[BTB.scala 105:81:@1348.4]
  assign _T_456 = {btb_valid_63,btb_valid_62,btb_valid_61,btb_valid_60,btb_valid_59,btb_valid_58,btb_valid_57,btb_valid_56,_T_447,_T_440}; // @[BTB.scala 105:81:@1357.4]
  assign _T_457 = {_T_456,_T_425}; // @[BTB.scala 105:81:@1358.4]
  assign predict_0_lookup = _T_394 & _T_457; // @[BTB.scala 105:69:@1359.4]
  assign _T_459 = predict_0_lookup[0]; // @[Mux.scala 21:36:@1361.4]
  assign _T_460 = predict_0_lookup[1]; // @[Mux.scala 21:36:@1362.4]
  assign _T_461 = predict_0_lookup[2]; // @[Mux.scala 21:36:@1363.4]
  assign _T_462 = predict_0_lookup[3]; // @[Mux.scala 21:36:@1364.4]
  assign _T_463 = predict_0_lookup[4]; // @[Mux.scala 21:36:@1365.4]
  assign _T_464 = predict_0_lookup[5]; // @[Mux.scala 21:36:@1366.4]
  assign _T_465 = predict_0_lookup[6]; // @[Mux.scala 21:36:@1367.4]
  assign _T_466 = predict_0_lookup[7]; // @[Mux.scala 21:36:@1368.4]
  assign _T_467 = predict_0_lookup[8]; // @[Mux.scala 21:36:@1369.4]
  assign _T_468 = predict_0_lookup[9]; // @[Mux.scala 21:36:@1370.4]
  assign _T_469 = predict_0_lookup[10]; // @[Mux.scala 21:36:@1371.4]
  assign _T_470 = predict_0_lookup[11]; // @[Mux.scala 21:36:@1372.4]
  assign _T_471 = predict_0_lookup[12]; // @[Mux.scala 21:36:@1373.4]
  assign _T_472 = predict_0_lookup[13]; // @[Mux.scala 21:36:@1374.4]
  assign _T_473 = predict_0_lookup[14]; // @[Mux.scala 21:36:@1375.4]
  assign _T_474 = predict_0_lookup[15]; // @[Mux.scala 21:36:@1376.4]
  assign _T_475 = predict_0_lookup[16]; // @[Mux.scala 21:36:@1377.4]
  assign _T_476 = predict_0_lookup[17]; // @[Mux.scala 21:36:@1378.4]
  assign _T_477 = predict_0_lookup[18]; // @[Mux.scala 21:36:@1379.4]
  assign _T_478 = predict_0_lookup[19]; // @[Mux.scala 21:36:@1380.4]
  assign _T_479 = predict_0_lookup[20]; // @[Mux.scala 21:36:@1381.4]
  assign _T_480 = predict_0_lookup[21]; // @[Mux.scala 21:36:@1382.4]
  assign _T_481 = predict_0_lookup[22]; // @[Mux.scala 21:36:@1383.4]
  assign _T_482 = predict_0_lookup[23]; // @[Mux.scala 21:36:@1384.4]
  assign _T_483 = predict_0_lookup[24]; // @[Mux.scala 21:36:@1385.4]
  assign _T_484 = predict_0_lookup[25]; // @[Mux.scala 21:36:@1386.4]
  assign _T_485 = predict_0_lookup[26]; // @[Mux.scala 21:36:@1387.4]
  assign _T_486 = predict_0_lookup[27]; // @[Mux.scala 21:36:@1388.4]
  assign _T_487 = predict_0_lookup[28]; // @[Mux.scala 21:36:@1389.4]
  assign _T_488 = predict_0_lookup[29]; // @[Mux.scala 21:36:@1390.4]
  assign _T_489 = predict_0_lookup[30]; // @[Mux.scala 21:36:@1391.4]
  assign _T_490 = predict_0_lookup[31]; // @[Mux.scala 21:36:@1392.4]
  assign _T_491 = predict_0_lookup[32]; // @[Mux.scala 21:36:@1393.4]
  assign _T_492 = predict_0_lookup[33]; // @[Mux.scala 21:36:@1394.4]
  assign _T_493 = predict_0_lookup[34]; // @[Mux.scala 21:36:@1395.4]
  assign _T_494 = predict_0_lookup[35]; // @[Mux.scala 21:36:@1396.4]
  assign _T_495 = predict_0_lookup[36]; // @[Mux.scala 21:36:@1397.4]
  assign _T_496 = predict_0_lookup[37]; // @[Mux.scala 21:36:@1398.4]
  assign _T_497 = predict_0_lookup[38]; // @[Mux.scala 21:36:@1399.4]
  assign _T_498 = predict_0_lookup[39]; // @[Mux.scala 21:36:@1400.4]
  assign _T_499 = predict_0_lookup[40]; // @[Mux.scala 21:36:@1401.4]
  assign _T_500 = predict_0_lookup[41]; // @[Mux.scala 21:36:@1402.4]
  assign _T_501 = predict_0_lookup[42]; // @[Mux.scala 21:36:@1403.4]
  assign _T_502 = predict_0_lookup[43]; // @[Mux.scala 21:36:@1404.4]
  assign _T_503 = predict_0_lookup[44]; // @[Mux.scala 21:36:@1405.4]
  assign _T_504 = predict_0_lookup[45]; // @[Mux.scala 21:36:@1406.4]
  assign _T_505 = predict_0_lookup[46]; // @[Mux.scala 21:36:@1407.4]
  assign _T_506 = predict_0_lookup[47]; // @[Mux.scala 21:36:@1408.4]
  assign _T_507 = predict_0_lookup[48]; // @[Mux.scala 21:36:@1409.4]
  assign _T_508 = predict_0_lookup[49]; // @[Mux.scala 21:36:@1410.4]
  assign _T_509 = predict_0_lookup[50]; // @[Mux.scala 21:36:@1411.4]
  assign _T_510 = predict_0_lookup[51]; // @[Mux.scala 21:36:@1412.4]
  assign _T_511 = predict_0_lookup[52]; // @[Mux.scala 21:36:@1413.4]
  assign _T_512 = predict_0_lookup[53]; // @[Mux.scala 21:36:@1414.4]
  assign _T_513 = predict_0_lookup[54]; // @[Mux.scala 21:36:@1415.4]
  assign _T_514 = predict_0_lookup[55]; // @[Mux.scala 21:36:@1416.4]
  assign _T_515 = predict_0_lookup[56]; // @[Mux.scala 21:36:@1417.4]
  assign _T_516 = predict_0_lookup[57]; // @[Mux.scala 21:36:@1418.4]
  assign _T_517 = predict_0_lookup[58]; // @[Mux.scala 21:36:@1419.4]
  assign _T_518 = predict_0_lookup[59]; // @[Mux.scala 21:36:@1420.4]
  assign _T_519 = predict_0_lookup[60]; // @[Mux.scala 21:36:@1421.4]
  assign _T_520 = predict_0_lookup[61]; // @[Mux.scala 21:36:@1422.4]
  assign _T_521 = predict_0_lookup[62]; // @[Mux.scala 21:36:@1423.4]
  assign _T_522 = predict_0_lookup[63]; // @[Mux.scala 21:36:@1424.4]
  assign _T_525 = _T_459 ? btb_tgt_0 : 30'h0; // @[Mux.scala 19:72:@1425.4]
  assign _T_527 = _T_460 ? btb_tgt_1 : 30'h0; // @[Mux.scala 19:72:@1426.4]
  assign _T_529 = _T_461 ? btb_tgt_2 : 30'h0; // @[Mux.scala 19:72:@1427.4]
  assign _T_531 = _T_462 ? btb_tgt_3 : 30'h0; // @[Mux.scala 19:72:@1428.4]
  assign _T_533 = _T_463 ? btb_tgt_4 : 30'h0; // @[Mux.scala 19:72:@1429.4]
  assign _T_535 = _T_464 ? btb_tgt_5 : 30'h0; // @[Mux.scala 19:72:@1430.4]
  assign _T_537 = _T_465 ? btb_tgt_6 : 30'h0; // @[Mux.scala 19:72:@1431.4]
  assign _T_539 = _T_466 ? btb_tgt_7 : 30'h0; // @[Mux.scala 19:72:@1432.4]
  assign _T_541 = _T_467 ? btb_tgt_8 : 30'h0; // @[Mux.scala 19:72:@1433.4]
  assign _T_543 = _T_468 ? btb_tgt_9 : 30'h0; // @[Mux.scala 19:72:@1434.4]
  assign _T_545 = _T_469 ? btb_tgt_10 : 30'h0; // @[Mux.scala 19:72:@1435.4]
  assign _T_547 = _T_470 ? btb_tgt_11 : 30'h0; // @[Mux.scala 19:72:@1436.4]
  assign _T_549 = _T_471 ? btb_tgt_12 : 30'h0; // @[Mux.scala 19:72:@1437.4]
  assign _T_551 = _T_472 ? btb_tgt_13 : 30'h0; // @[Mux.scala 19:72:@1438.4]
  assign _T_553 = _T_473 ? btb_tgt_14 : 30'h0; // @[Mux.scala 19:72:@1439.4]
  assign _T_555 = _T_474 ? btb_tgt_15 : 30'h0; // @[Mux.scala 19:72:@1440.4]
  assign _T_557 = _T_475 ? btb_tgt_16 : 30'h0; // @[Mux.scala 19:72:@1441.4]
  assign _T_559 = _T_476 ? btb_tgt_17 : 30'h0; // @[Mux.scala 19:72:@1442.4]
  assign _T_561 = _T_477 ? btb_tgt_18 : 30'h0; // @[Mux.scala 19:72:@1443.4]
  assign _T_563 = _T_478 ? btb_tgt_19 : 30'h0; // @[Mux.scala 19:72:@1444.4]
  assign _T_565 = _T_479 ? btb_tgt_20 : 30'h0; // @[Mux.scala 19:72:@1445.4]
  assign _T_567 = _T_480 ? btb_tgt_21 : 30'h0; // @[Mux.scala 19:72:@1446.4]
  assign _T_569 = _T_481 ? btb_tgt_22 : 30'h0; // @[Mux.scala 19:72:@1447.4]
  assign _T_571 = _T_482 ? btb_tgt_23 : 30'h0; // @[Mux.scala 19:72:@1448.4]
  assign _T_573 = _T_483 ? btb_tgt_24 : 30'h0; // @[Mux.scala 19:72:@1449.4]
  assign _T_575 = _T_484 ? btb_tgt_25 : 30'h0; // @[Mux.scala 19:72:@1450.4]
  assign _T_577 = _T_485 ? btb_tgt_26 : 30'h0; // @[Mux.scala 19:72:@1451.4]
  assign _T_579 = _T_486 ? btb_tgt_27 : 30'h0; // @[Mux.scala 19:72:@1452.4]
  assign _T_581 = _T_487 ? btb_tgt_28 : 30'h0; // @[Mux.scala 19:72:@1453.4]
  assign _T_583 = _T_488 ? btb_tgt_29 : 30'h0; // @[Mux.scala 19:72:@1454.4]
  assign _T_585 = _T_489 ? btb_tgt_30 : 30'h0; // @[Mux.scala 19:72:@1455.4]
  assign _T_587 = _T_490 ? btb_tgt_31 : 30'h0; // @[Mux.scala 19:72:@1456.4]
  assign _T_589 = _T_491 ? btb_tgt_32 : 30'h0; // @[Mux.scala 19:72:@1457.4]
  assign _T_591 = _T_492 ? btb_tgt_33 : 30'h0; // @[Mux.scala 19:72:@1458.4]
  assign _T_593 = _T_493 ? btb_tgt_34 : 30'h0; // @[Mux.scala 19:72:@1459.4]
  assign _T_595 = _T_494 ? btb_tgt_35 : 30'h0; // @[Mux.scala 19:72:@1460.4]
  assign _T_597 = _T_495 ? btb_tgt_36 : 30'h0; // @[Mux.scala 19:72:@1461.4]
  assign _T_599 = _T_496 ? btb_tgt_37 : 30'h0; // @[Mux.scala 19:72:@1462.4]
  assign _T_601 = _T_497 ? btb_tgt_38 : 30'h0; // @[Mux.scala 19:72:@1463.4]
  assign _T_603 = _T_498 ? btb_tgt_39 : 30'h0; // @[Mux.scala 19:72:@1464.4]
  assign _T_605 = _T_499 ? btb_tgt_40 : 30'h0; // @[Mux.scala 19:72:@1465.4]
  assign _T_607 = _T_500 ? btb_tgt_41 : 30'h0; // @[Mux.scala 19:72:@1466.4]
  assign _T_609 = _T_501 ? btb_tgt_42 : 30'h0; // @[Mux.scala 19:72:@1467.4]
  assign _T_611 = _T_502 ? btb_tgt_43 : 30'h0; // @[Mux.scala 19:72:@1468.4]
  assign _T_613 = _T_503 ? btb_tgt_44 : 30'h0; // @[Mux.scala 19:72:@1469.4]
  assign _T_615 = _T_504 ? btb_tgt_45 : 30'h0; // @[Mux.scala 19:72:@1470.4]
  assign _T_617 = _T_505 ? btb_tgt_46 : 30'h0; // @[Mux.scala 19:72:@1471.4]
  assign _T_619 = _T_506 ? btb_tgt_47 : 30'h0; // @[Mux.scala 19:72:@1472.4]
  assign _T_621 = _T_507 ? btb_tgt_48 : 30'h0; // @[Mux.scala 19:72:@1473.4]
  assign _T_623 = _T_508 ? btb_tgt_49 : 30'h0; // @[Mux.scala 19:72:@1474.4]
  assign _T_625 = _T_509 ? btb_tgt_50 : 30'h0; // @[Mux.scala 19:72:@1475.4]
  assign _T_627 = _T_510 ? btb_tgt_51 : 30'h0; // @[Mux.scala 19:72:@1476.4]
  assign _T_629 = _T_511 ? btb_tgt_52 : 30'h0; // @[Mux.scala 19:72:@1477.4]
  assign _T_631 = _T_512 ? btb_tgt_53 : 30'h0; // @[Mux.scala 19:72:@1478.4]
  assign _T_633 = _T_513 ? btb_tgt_54 : 30'h0; // @[Mux.scala 19:72:@1479.4]
  assign _T_635 = _T_514 ? btb_tgt_55 : 30'h0; // @[Mux.scala 19:72:@1480.4]
  assign _T_637 = _T_515 ? btb_tgt_56 : 30'h0; // @[Mux.scala 19:72:@1481.4]
  assign _T_639 = _T_516 ? btb_tgt_57 : 30'h0; // @[Mux.scala 19:72:@1482.4]
  assign _T_641 = _T_517 ? btb_tgt_58 : 30'h0; // @[Mux.scala 19:72:@1483.4]
  assign _T_643 = _T_518 ? btb_tgt_59 : 30'h0; // @[Mux.scala 19:72:@1484.4]
  assign _T_645 = _T_519 ? btb_tgt_60 : 30'h0; // @[Mux.scala 19:72:@1485.4]
  assign _T_647 = _T_520 ? btb_tgt_61 : 30'h0; // @[Mux.scala 19:72:@1486.4]
  assign _T_649 = _T_521 ? btb_tgt_62 : 30'h0; // @[Mux.scala 19:72:@1487.4]
  assign _T_651 = _T_522 ? btb_tgt_63 : 30'h0; // @[Mux.scala 19:72:@1488.4]
  assign _T_652 = _T_525 | _T_527; // @[Mux.scala 19:72:@1489.4]
  assign _T_653 = _T_652 | _T_529; // @[Mux.scala 19:72:@1490.4]
  assign _T_654 = _T_653 | _T_531; // @[Mux.scala 19:72:@1491.4]
  assign _T_655 = _T_654 | _T_533; // @[Mux.scala 19:72:@1492.4]
  assign _T_656 = _T_655 | _T_535; // @[Mux.scala 19:72:@1493.4]
  assign _T_657 = _T_656 | _T_537; // @[Mux.scala 19:72:@1494.4]
  assign _T_658 = _T_657 | _T_539; // @[Mux.scala 19:72:@1495.4]
  assign _T_659 = _T_658 | _T_541; // @[Mux.scala 19:72:@1496.4]
  assign _T_660 = _T_659 | _T_543; // @[Mux.scala 19:72:@1497.4]
  assign _T_661 = _T_660 | _T_545; // @[Mux.scala 19:72:@1498.4]
  assign _T_662 = _T_661 | _T_547; // @[Mux.scala 19:72:@1499.4]
  assign _T_663 = _T_662 | _T_549; // @[Mux.scala 19:72:@1500.4]
  assign _T_664 = _T_663 | _T_551; // @[Mux.scala 19:72:@1501.4]
  assign _T_665 = _T_664 | _T_553; // @[Mux.scala 19:72:@1502.4]
  assign _T_666 = _T_665 | _T_555; // @[Mux.scala 19:72:@1503.4]
  assign _T_667 = _T_666 | _T_557; // @[Mux.scala 19:72:@1504.4]
  assign _T_668 = _T_667 | _T_559; // @[Mux.scala 19:72:@1505.4]
  assign _T_669 = _T_668 | _T_561; // @[Mux.scala 19:72:@1506.4]
  assign _T_670 = _T_669 | _T_563; // @[Mux.scala 19:72:@1507.4]
  assign _T_671 = _T_670 | _T_565; // @[Mux.scala 19:72:@1508.4]
  assign _T_672 = _T_671 | _T_567; // @[Mux.scala 19:72:@1509.4]
  assign _T_673 = _T_672 | _T_569; // @[Mux.scala 19:72:@1510.4]
  assign _T_674 = _T_673 | _T_571; // @[Mux.scala 19:72:@1511.4]
  assign _T_675 = _T_674 | _T_573; // @[Mux.scala 19:72:@1512.4]
  assign _T_676 = _T_675 | _T_575; // @[Mux.scala 19:72:@1513.4]
  assign _T_677 = _T_676 | _T_577; // @[Mux.scala 19:72:@1514.4]
  assign _T_678 = _T_677 | _T_579; // @[Mux.scala 19:72:@1515.4]
  assign _T_679 = _T_678 | _T_581; // @[Mux.scala 19:72:@1516.4]
  assign _T_680 = _T_679 | _T_583; // @[Mux.scala 19:72:@1517.4]
  assign _T_681 = _T_680 | _T_585; // @[Mux.scala 19:72:@1518.4]
  assign _T_682 = _T_681 | _T_587; // @[Mux.scala 19:72:@1519.4]
  assign _T_683 = _T_682 | _T_589; // @[Mux.scala 19:72:@1520.4]
  assign _T_684 = _T_683 | _T_591; // @[Mux.scala 19:72:@1521.4]
  assign _T_685 = _T_684 | _T_593; // @[Mux.scala 19:72:@1522.4]
  assign _T_686 = _T_685 | _T_595; // @[Mux.scala 19:72:@1523.4]
  assign _T_687 = _T_686 | _T_597; // @[Mux.scala 19:72:@1524.4]
  assign _T_688 = _T_687 | _T_599; // @[Mux.scala 19:72:@1525.4]
  assign _T_689 = _T_688 | _T_601; // @[Mux.scala 19:72:@1526.4]
  assign _T_690 = _T_689 | _T_603; // @[Mux.scala 19:72:@1527.4]
  assign _T_691 = _T_690 | _T_605; // @[Mux.scala 19:72:@1528.4]
  assign _T_692 = _T_691 | _T_607; // @[Mux.scala 19:72:@1529.4]
  assign _T_693 = _T_692 | _T_609; // @[Mux.scala 19:72:@1530.4]
  assign _T_694 = _T_693 | _T_611; // @[Mux.scala 19:72:@1531.4]
  assign _T_695 = _T_694 | _T_613; // @[Mux.scala 19:72:@1532.4]
  assign _T_696 = _T_695 | _T_615; // @[Mux.scala 19:72:@1533.4]
  assign _T_697 = _T_696 | _T_617; // @[Mux.scala 19:72:@1534.4]
  assign _T_698 = _T_697 | _T_619; // @[Mux.scala 19:72:@1535.4]
  assign _T_699 = _T_698 | _T_621; // @[Mux.scala 19:72:@1536.4]
  assign _T_700 = _T_699 | _T_623; // @[Mux.scala 19:72:@1537.4]
  assign _T_701 = _T_700 | _T_625; // @[Mux.scala 19:72:@1538.4]
  assign _T_702 = _T_701 | _T_627; // @[Mux.scala 19:72:@1539.4]
  assign _T_703 = _T_702 | _T_629; // @[Mux.scala 19:72:@1540.4]
  assign _T_704 = _T_703 | _T_631; // @[Mux.scala 19:72:@1541.4]
  assign _T_705 = _T_704 | _T_633; // @[Mux.scala 19:72:@1542.4]
  assign _T_706 = _T_705 | _T_635; // @[Mux.scala 19:72:@1543.4]
  assign _T_707 = _T_706 | _T_637; // @[Mux.scala 19:72:@1544.4]
  assign _T_708 = _T_707 | _T_639; // @[Mux.scala 19:72:@1545.4]
  assign _T_709 = _T_708 | _T_641; // @[Mux.scala 19:72:@1546.4]
  assign _T_710 = _T_709 | _T_643; // @[Mux.scala 19:72:@1547.4]
  assign _T_711 = _T_710 | _T_645; // @[Mux.scala 19:72:@1548.4]
  assign _T_712 = _T_711 | _T_647; // @[Mux.scala 19:72:@1549.4]
  assign _T_713 = _T_712 | _T_649; // @[Mux.scala 19:72:@1550.4]
  assign _T_714 = _T_713 | _T_651; // @[Mux.scala 19:72:@1551.4]
  assign predict_0_jump_tgt = {_T_714,2'h0}; // @[Cat.scala 30:58:@1554.4]
  assign _T_785 = _T_459 ? btb_bj_type_0 : 2'h0; // @[Mux.scala 19:72:@1620.4]
  assign _T_787 = _T_460 ? btb_bj_type_1 : 2'h0; // @[Mux.scala 19:72:@1621.4]
  assign _T_789 = _T_461 ? btb_bj_type_2 : 2'h0; // @[Mux.scala 19:72:@1622.4]
  assign _T_791 = _T_462 ? btb_bj_type_3 : 2'h0; // @[Mux.scala 19:72:@1623.4]
  assign _T_793 = _T_463 ? btb_bj_type_4 : 2'h0; // @[Mux.scala 19:72:@1624.4]
  assign _T_795 = _T_464 ? btb_bj_type_5 : 2'h0; // @[Mux.scala 19:72:@1625.4]
  assign _T_797 = _T_465 ? btb_bj_type_6 : 2'h0; // @[Mux.scala 19:72:@1626.4]
  assign _T_799 = _T_466 ? btb_bj_type_7 : 2'h0; // @[Mux.scala 19:72:@1627.4]
  assign _T_801 = _T_467 ? btb_bj_type_8 : 2'h0; // @[Mux.scala 19:72:@1628.4]
  assign _T_803 = _T_468 ? btb_bj_type_9 : 2'h0; // @[Mux.scala 19:72:@1629.4]
  assign _T_805 = _T_469 ? btb_bj_type_10 : 2'h0; // @[Mux.scala 19:72:@1630.4]
  assign _T_807 = _T_470 ? btb_bj_type_11 : 2'h0; // @[Mux.scala 19:72:@1631.4]
  assign _T_809 = _T_471 ? btb_bj_type_12 : 2'h0; // @[Mux.scala 19:72:@1632.4]
  assign _T_811 = _T_472 ? btb_bj_type_13 : 2'h0; // @[Mux.scala 19:72:@1633.4]
  assign _T_813 = _T_473 ? btb_bj_type_14 : 2'h0; // @[Mux.scala 19:72:@1634.4]
  assign _T_815 = _T_474 ? btb_bj_type_15 : 2'h0; // @[Mux.scala 19:72:@1635.4]
  assign _T_817 = _T_475 ? btb_bj_type_16 : 2'h0; // @[Mux.scala 19:72:@1636.4]
  assign _T_819 = _T_476 ? btb_bj_type_17 : 2'h0; // @[Mux.scala 19:72:@1637.4]
  assign _T_821 = _T_477 ? btb_bj_type_18 : 2'h0; // @[Mux.scala 19:72:@1638.4]
  assign _T_823 = _T_478 ? btb_bj_type_19 : 2'h0; // @[Mux.scala 19:72:@1639.4]
  assign _T_825 = _T_479 ? btb_bj_type_20 : 2'h0; // @[Mux.scala 19:72:@1640.4]
  assign _T_827 = _T_480 ? btb_bj_type_21 : 2'h0; // @[Mux.scala 19:72:@1641.4]
  assign _T_829 = _T_481 ? btb_bj_type_22 : 2'h0; // @[Mux.scala 19:72:@1642.4]
  assign _T_831 = _T_482 ? btb_bj_type_23 : 2'h0; // @[Mux.scala 19:72:@1643.4]
  assign _T_833 = _T_483 ? btb_bj_type_24 : 2'h0; // @[Mux.scala 19:72:@1644.4]
  assign _T_835 = _T_484 ? btb_bj_type_25 : 2'h0; // @[Mux.scala 19:72:@1645.4]
  assign _T_837 = _T_485 ? btb_bj_type_26 : 2'h0; // @[Mux.scala 19:72:@1646.4]
  assign _T_839 = _T_486 ? btb_bj_type_27 : 2'h0; // @[Mux.scala 19:72:@1647.4]
  assign _T_841 = _T_487 ? btb_bj_type_28 : 2'h0; // @[Mux.scala 19:72:@1648.4]
  assign _T_843 = _T_488 ? btb_bj_type_29 : 2'h0; // @[Mux.scala 19:72:@1649.4]
  assign _T_845 = _T_489 ? btb_bj_type_30 : 2'h0; // @[Mux.scala 19:72:@1650.4]
  assign _T_847 = _T_490 ? btb_bj_type_31 : 2'h0; // @[Mux.scala 19:72:@1651.4]
  assign _T_849 = _T_491 ? btb_bj_type_32 : 2'h0; // @[Mux.scala 19:72:@1652.4]
  assign _T_851 = _T_492 ? btb_bj_type_33 : 2'h0; // @[Mux.scala 19:72:@1653.4]
  assign _T_853 = _T_493 ? btb_bj_type_34 : 2'h0; // @[Mux.scala 19:72:@1654.4]
  assign _T_855 = _T_494 ? btb_bj_type_35 : 2'h0; // @[Mux.scala 19:72:@1655.4]
  assign _T_857 = _T_495 ? btb_bj_type_36 : 2'h0; // @[Mux.scala 19:72:@1656.4]
  assign _T_859 = _T_496 ? btb_bj_type_37 : 2'h0; // @[Mux.scala 19:72:@1657.4]
  assign _T_861 = _T_497 ? btb_bj_type_38 : 2'h0; // @[Mux.scala 19:72:@1658.4]
  assign _T_863 = _T_498 ? btb_bj_type_39 : 2'h0; // @[Mux.scala 19:72:@1659.4]
  assign _T_865 = _T_499 ? btb_bj_type_40 : 2'h0; // @[Mux.scala 19:72:@1660.4]
  assign _T_867 = _T_500 ? btb_bj_type_41 : 2'h0; // @[Mux.scala 19:72:@1661.4]
  assign _T_869 = _T_501 ? btb_bj_type_42 : 2'h0; // @[Mux.scala 19:72:@1662.4]
  assign _T_871 = _T_502 ? btb_bj_type_43 : 2'h0; // @[Mux.scala 19:72:@1663.4]
  assign _T_873 = _T_503 ? btb_bj_type_44 : 2'h0; // @[Mux.scala 19:72:@1664.4]
  assign _T_875 = _T_504 ? btb_bj_type_45 : 2'h0; // @[Mux.scala 19:72:@1665.4]
  assign _T_877 = _T_505 ? btb_bj_type_46 : 2'h0; // @[Mux.scala 19:72:@1666.4]
  assign _T_879 = _T_506 ? btb_bj_type_47 : 2'h0; // @[Mux.scala 19:72:@1667.4]
  assign _T_881 = _T_507 ? btb_bj_type_48 : 2'h0; // @[Mux.scala 19:72:@1668.4]
  assign _T_883 = _T_508 ? btb_bj_type_49 : 2'h0; // @[Mux.scala 19:72:@1669.4]
  assign _T_885 = _T_509 ? btb_bj_type_50 : 2'h0; // @[Mux.scala 19:72:@1670.4]
  assign _T_887 = _T_510 ? btb_bj_type_51 : 2'h0; // @[Mux.scala 19:72:@1671.4]
  assign _T_889 = _T_511 ? btb_bj_type_52 : 2'h0; // @[Mux.scala 19:72:@1672.4]
  assign _T_891 = _T_512 ? btb_bj_type_53 : 2'h0; // @[Mux.scala 19:72:@1673.4]
  assign _T_893 = _T_513 ? btb_bj_type_54 : 2'h0; // @[Mux.scala 19:72:@1674.4]
  assign _T_895 = _T_514 ? btb_bj_type_55 : 2'h0; // @[Mux.scala 19:72:@1675.4]
  assign _T_897 = _T_515 ? btb_bj_type_56 : 2'h0; // @[Mux.scala 19:72:@1676.4]
  assign _T_899 = _T_516 ? btb_bj_type_57 : 2'h0; // @[Mux.scala 19:72:@1677.4]
  assign _T_901 = _T_517 ? btb_bj_type_58 : 2'h0; // @[Mux.scala 19:72:@1678.4]
  assign _T_903 = _T_518 ? btb_bj_type_59 : 2'h0; // @[Mux.scala 19:72:@1679.4]
  assign _T_905 = _T_519 ? btb_bj_type_60 : 2'h0; // @[Mux.scala 19:72:@1680.4]
  assign _T_907 = _T_520 ? btb_bj_type_61 : 2'h0; // @[Mux.scala 19:72:@1681.4]
  assign _T_909 = _T_521 ? btb_bj_type_62 : 2'h0; // @[Mux.scala 19:72:@1682.4]
  assign _T_911 = _T_522 ? btb_bj_type_63 : 2'h0; // @[Mux.scala 19:72:@1683.4]
  assign _T_912 = _T_785 | _T_787; // @[Mux.scala 19:72:@1684.4]
  assign _T_913 = _T_912 | _T_789; // @[Mux.scala 19:72:@1685.4]
  assign _T_914 = _T_913 | _T_791; // @[Mux.scala 19:72:@1686.4]
  assign _T_915 = _T_914 | _T_793; // @[Mux.scala 19:72:@1687.4]
  assign _T_916 = _T_915 | _T_795; // @[Mux.scala 19:72:@1688.4]
  assign _T_917 = _T_916 | _T_797; // @[Mux.scala 19:72:@1689.4]
  assign _T_918 = _T_917 | _T_799; // @[Mux.scala 19:72:@1690.4]
  assign _T_919 = _T_918 | _T_801; // @[Mux.scala 19:72:@1691.4]
  assign _T_920 = _T_919 | _T_803; // @[Mux.scala 19:72:@1692.4]
  assign _T_921 = _T_920 | _T_805; // @[Mux.scala 19:72:@1693.4]
  assign _T_922 = _T_921 | _T_807; // @[Mux.scala 19:72:@1694.4]
  assign _T_923 = _T_922 | _T_809; // @[Mux.scala 19:72:@1695.4]
  assign _T_924 = _T_923 | _T_811; // @[Mux.scala 19:72:@1696.4]
  assign _T_925 = _T_924 | _T_813; // @[Mux.scala 19:72:@1697.4]
  assign _T_926 = _T_925 | _T_815; // @[Mux.scala 19:72:@1698.4]
  assign _T_927 = _T_926 | _T_817; // @[Mux.scala 19:72:@1699.4]
  assign _T_928 = _T_927 | _T_819; // @[Mux.scala 19:72:@1700.4]
  assign _T_929 = _T_928 | _T_821; // @[Mux.scala 19:72:@1701.4]
  assign _T_930 = _T_929 | _T_823; // @[Mux.scala 19:72:@1702.4]
  assign _T_931 = _T_930 | _T_825; // @[Mux.scala 19:72:@1703.4]
  assign _T_932 = _T_931 | _T_827; // @[Mux.scala 19:72:@1704.4]
  assign _T_933 = _T_932 | _T_829; // @[Mux.scala 19:72:@1705.4]
  assign _T_934 = _T_933 | _T_831; // @[Mux.scala 19:72:@1706.4]
  assign _T_935 = _T_934 | _T_833; // @[Mux.scala 19:72:@1707.4]
  assign _T_936 = _T_935 | _T_835; // @[Mux.scala 19:72:@1708.4]
  assign _T_937 = _T_936 | _T_837; // @[Mux.scala 19:72:@1709.4]
  assign _T_938 = _T_937 | _T_839; // @[Mux.scala 19:72:@1710.4]
  assign _T_939 = _T_938 | _T_841; // @[Mux.scala 19:72:@1711.4]
  assign _T_940 = _T_939 | _T_843; // @[Mux.scala 19:72:@1712.4]
  assign _T_941 = _T_940 | _T_845; // @[Mux.scala 19:72:@1713.4]
  assign _T_942 = _T_941 | _T_847; // @[Mux.scala 19:72:@1714.4]
  assign _T_943 = _T_942 | _T_849; // @[Mux.scala 19:72:@1715.4]
  assign _T_944 = _T_943 | _T_851; // @[Mux.scala 19:72:@1716.4]
  assign _T_945 = _T_944 | _T_853; // @[Mux.scala 19:72:@1717.4]
  assign _T_946 = _T_945 | _T_855; // @[Mux.scala 19:72:@1718.4]
  assign _T_947 = _T_946 | _T_857; // @[Mux.scala 19:72:@1719.4]
  assign _T_948 = _T_947 | _T_859; // @[Mux.scala 19:72:@1720.4]
  assign _T_949 = _T_948 | _T_861; // @[Mux.scala 19:72:@1721.4]
  assign _T_950 = _T_949 | _T_863; // @[Mux.scala 19:72:@1722.4]
  assign _T_951 = _T_950 | _T_865; // @[Mux.scala 19:72:@1723.4]
  assign _T_952 = _T_951 | _T_867; // @[Mux.scala 19:72:@1724.4]
  assign _T_953 = _T_952 | _T_869; // @[Mux.scala 19:72:@1725.4]
  assign _T_954 = _T_953 | _T_871; // @[Mux.scala 19:72:@1726.4]
  assign _T_955 = _T_954 | _T_873; // @[Mux.scala 19:72:@1727.4]
  assign _T_956 = _T_955 | _T_875; // @[Mux.scala 19:72:@1728.4]
  assign _T_957 = _T_956 | _T_877; // @[Mux.scala 19:72:@1729.4]
  assign _T_958 = _T_957 | _T_879; // @[Mux.scala 19:72:@1730.4]
  assign _T_959 = _T_958 | _T_881; // @[Mux.scala 19:72:@1731.4]
  assign _T_960 = _T_959 | _T_883; // @[Mux.scala 19:72:@1732.4]
  assign _T_961 = _T_960 | _T_885; // @[Mux.scala 19:72:@1733.4]
  assign _T_962 = _T_961 | _T_887; // @[Mux.scala 19:72:@1734.4]
  assign _T_963 = _T_962 | _T_889; // @[Mux.scala 19:72:@1735.4]
  assign _T_964 = _T_963 | _T_891; // @[Mux.scala 19:72:@1736.4]
  assign _T_965 = _T_964 | _T_893; // @[Mux.scala 19:72:@1737.4]
  assign _T_966 = _T_965 | _T_895; // @[Mux.scala 19:72:@1738.4]
  assign _T_967 = _T_966 | _T_897; // @[Mux.scala 19:72:@1739.4]
  assign _T_968 = _T_967 | _T_899; // @[Mux.scala 19:72:@1740.4]
  assign _T_969 = _T_968 | _T_901; // @[Mux.scala 19:72:@1741.4]
  assign _T_970 = _T_969 | _T_903; // @[Mux.scala 19:72:@1742.4]
  assign _T_971 = _T_970 | _T_905; // @[Mux.scala 19:72:@1743.4]
  assign _T_972 = _T_971 | _T_907; // @[Mux.scala 19:72:@1744.4]
  assign _T_973 = _T_972 | _T_909; // @[Mux.scala 19:72:@1745.4]
  assign predict_0_bj_type = _T_973 | _T_911; // @[Mux.scala 19:72:@1746.4]
  assign _T_1043 = _T_459 ? btb_h_count_0 : 2'h0; // @[Mux.scala 19:72:@1814.4]
  assign _T_1045 = _T_460 ? btb_h_count_1 : 2'h0; // @[Mux.scala 19:72:@1815.4]
  assign _T_1047 = _T_461 ? btb_h_count_2 : 2'h0; // @[Mux.scala 19:72:@1816.4]
  assign _T_1049 = _T_462 ? btb_h_count_3 : 2'h0; // @[Mux.scala 19:72:@1817.4]
  assign _T_1051 = _T_463 ? btb_h_count_4 : 2'h0; // @[Mux.scala 19:72:@1818.4]
  assign _T_1053 = _T_464 ? btb_h_count_5 : 2'h0; // @[Mux.scala 19:72:@1819.4]
  assign _T_1055 = _T_465 ? btb_h_count_6 : 2'h0; // @[Mux.scala 19:72:@1820.4]
  assign _T_1057 = _T_466 ? btb_h_count_7 : 2'h0; // @[Mux.scala 19:72:@1821.4]
  assign _T_1059 = _T_467 ? btb_h_count_8 : 2'h0; // @[Mux.scala 19:72:@1822.4]
  assign _T_1061 = _T_468 ? btb_h_count_9 : 2'h0; // @[Mux.scala 19:72:@1823.4]
  assign _T_1063 = _T_469 ? btb_h_count_10 : 2'h0; // @[Mux.scala 19:72:@1824.4]
  assign _T_1065 = _T_470 ? btb_h_count_11 : 2'h0; // @[Mux.scala 19:72:@1825.4]
  assign _T_1067 = _T_471 ? btb_h_count_12 : 2'h0; // @[Mux.scala 19:72:@1826.4]
  assign _T_1069 = _T_472 ? btb_h_count_13 : 2'h0; // @[Mux.scala 19:72:@1827.4]
  assign _T_1071 = _T_473 ? btb_h_count_14 : 2'h0; // @[Mux.scala 19:72:@1828.4]
  assign _T_1073 = _T_474 ? btb_h_count_15 : 2'h0; // @[Mux.scala 19:72:@1829.4]
  assign _T_1075 = _T_475 ? btb_h_count_16 : 2'h0; // @[Mux.scala 19:72:@1830.4]
  assign _T_1077 = _T_476 ? btb_h_count_17 : 2'h0; // @[Mux.scala 19:72:@1831.4]
  assign _T_1079 = _T_477 ? btb_h_count_18 : 2'h0; // @[Mux.scala 19:72:@1832.4]
  assign _T_1081 = _T_478 ? btb_h_count_19 : 2'h0; // @[Mux.scala 19:72:@1833.4]
  assign _T_1083 = _T_479 ? btb_h_count_20 : 2'h0; // @[Mux.scala 19:72:@1834.4]
  assign _T_1085 = _T_480 ? btb_h_count_21 : 2'h0; // @[Mux.scala 19:72:@1835.4]
  assign _T_1087 = _T_481 ? btb_h_count_22 : 2'h0; // @[Mux.scala 19:72:@1836.4]
  assign _T_1089 = _T_482 ? btb_h_count_23 : 2'h0; // @[Mux.scala 19:72:@1837.4]
  assign _T_1091 = _T_483 ? btb_h_count_24 : 2'h0; // @[Mux.scala 19:72:@1838.4]
  assign _T_1093 = _T_484 ? btb_h_count_25 : 2'h0; // @[Mux.scala 19:72:@1839.4]
  assign _T_1095 = _T_485 ? btb_h_count_26 : 2'h0; // @[Mux.scala 19:72:@1840.4]
  assign _T_1097 = _T_486 ? btb_h_count_27 : 2'h0; // @[Mux.scala 19:72:@1841.4]
  assign _T_1099 = _T_487 ? btb_h_count_28 : 2'h0; // @[Mux.scala 19:72:@1842.4]
  assign _T_1101 = _T_488 ? btb_h_count_29 : 2'h0; // @[Mux.scala 19:72:@1843.4]
  assign _T_1103 = _T_489 ? btb_h_count_30 : 2'h0; // @[Mux.scala 19:72:@1844.4]
  assign _T_1105 = _T_490 ? btb_h_count_31 : 2'h0; // @[Mux.scala 19:72:@1845.4]
  assign _T_1107 = _T_491 ? btb_h_count_32 : 2'h0; // @[Mux.scala 19:72:@1846.4]
  assign _T_1109 = _T_492 ? btb_h_count_33 : 2'h0; // @[Mux.scala 19:72:@1847.4]
  assign _T_1111 = _T_493 ? btb_h_count_34 : 2'h0; // @[Mux.scala 19:72:@1848.4]
  assign _T_1113 = _T_494 ? btb_h_count_35 : 2'h0; // @[Mux.scala 19:72:@1849.4]
  assign _T_1115 = _T_495 ? btb_h_count_36 : 2'h0; // @[Mux.scala 19:72:@1850.4]
  assign _T_1117 = _T_496 ? btb_h_count_37 : 2'h0; // @[Mux.scala 19:72:@1851.4]
  assign _T_1119 = _T_497 ? btb_h_count_38 : 2'h0; // @[Mux.scala 19:72:@1852.4]
  assign _T_1121 = _T_498 ? btb_h_count_39 : 2'h0; // @[Mux.scala 19:72:@1853.4]
  assign _T_1123 = _T_499 ? btb_h_count_40 : 2'h0; // @[Mux.scala 19:72:@1854.4]
  assign _T_1125 = _T_500 ? btb_h_count_41 : 2'h0; // @[Mux.scala 19:72:@1855.4]
  assign _T_1127 = _T_501 ? btb_h_count_42 : 2'h0; // @[Mux.scala 19:72:@1856.4]
  assign _T_1129 = _T_502 ? btb_h_count_43 : 2'h0; // @[Mux.scala 19:72:@1857.4]
  assign _T_1131 = _T_503 ? btb_h_count_44 : 2'h0; // @[Mux.scala 19:72:@1858.4]
  assign _T_1133 = _T_504 ? btb_h_count_45 : 2'h0; // @[Mux.scala 19:72:@1859.4]
  assign _T_1135 = _T_505 ? btb_h_count_46 : 2'h0; // @[Mux.scala 19:72:@1860.4]
  assign _T_1137 = _T_506 ? btb_h_count_47 : 2'h0; // @[Mux.scala 19:72:@1861.4]
  assign _T_1139 = _T_507 ? btb_h_count_48 : 2'h0; // @[Mux.scala 19:72:@1862.4]
  assign _T_1141 = _T_508 ? btb_h_count_49 : 2'h0; // @[Mux.scala 19:72:@1863.4]
  assign _T_1143 = _T_509 ? btb_h_count_50 : 2'h0; // @[Mux.scala 19:72:@1864.4]
  assign _T_1145 = _T_510 ? btb_h_count_51 : 2'h0; // @[Mux.scala 19:72:@1865.4]
  assign _T_1147 = _T_511 ? btb_h_count_52 : 2'h0; // @[Mux.scala 19:72:@1866.4]
  assign _T_1149 = _T_512 ? btb_h_count_53 : 2'h0; // @[Mux.scala 19:72:@1867.4]
  assign _T_1151 = _T_513 ? btb_h_count_54 : 2'h0; // @[Mux.scala 19:72:@1868.4]
  assign _T_1153 = _T_514 ? btb_h_count_55 : 2'h0; // @[Mux.scala 19:72:@1869.4]
  assign _T_1155 = _T_515 ? btb_h_count_56 : 2'h0; // @[Mux.scala 19:72:@1870.4]
  assign _T_1157 = _T_516 ? btb_h_count_57 : 2'h0; // @[Mux.scala 19:72:@1871.4]
  assign _T_1159 = _T_517 ? btb_h_count_58 : 2'h0; // @[Mux.scala 19:72:@1872.4]
  assign _T_1161 = _T_518 ? btb_h_count_59 : 2'h0; // @[Mux.scala 19:72:@1873.4]
  assign _T_1163 = _T_519 ? btb_h_count_60 : 2'h0; // @[Mux.scala 19:72:@1874.4]
  assign _T_1165 = _T_520 ? btb_h_count_61 : 2'h0; // @[Mux.scala 19:72:@1875.4]
  assign _T_1167 = _T_521 ? btb_h_count_62 : 2'h0; // @[Mux.scala 19:72:@1876.4]
  assign _T_1169 = _T_522 ? btb_h_count_63 : 2'h0; // @[Mux.scala 19:72:@1877.4]
  assign _T_1170 = _T_1043 | _T_1045; // @[Mux.scala 19:72:@1878.4]
  assign _T_1171 = _T_1170 | _T_1047; // @[Mux.scala 19:72:@1879.4]
  assign _T_1172 = _T_1171 | _T_1049; // @[Mux.scala 19:72:@1880.4]
  assign _T_1173 = _T_1172 | _T_1051; // @[Mux.scala 19:72:@1881.4]
  assign _T_1174 = _T_1173 | _T_1053; // @[Mux.scala 19:72:@1882.4]
  assign _T_1175 = _T_1174 | _T_1055; // @[Mux.scala 19:72:@1883.4]
  assign _T_1176 = _T_1175 | _T_1057; // @[Mux.scala 19:72:@1884.4]
  assign _T_1177 = _T_1176 | _T_1059; // @[Mux.scala 19:72:@1885.4]
  assign _T_1178 = _T_1177 | _T_1061; // @[Mux.scala 19:72:@1886.4]
  assign _T_1179 = _T_1178 | _T_1063; // @[Mux.scala 19:72:@1887.4]
  assign _T_1180 = _T_1179 | _T_1065; // @[Mux.scala 19:72:@1888.4]
  assign _T_1181 = _T_1180 | _T_1067; // @[Mux.scala 19:72:@1889.4]
  assign _T_1182 = _T_1181 | _T_1069; // @[Mux.scala 19:72:@1890.4]
  assign _T_1183 = _T_1182 | _T_1071; // @[Mux.scala 19:72:@1891.4]
  assign _T_1184 = _T_1183 | _T_1073; // @[Mux.scala 19:72:@1892.4]
  assign _T_1185 = _T_1184 | _T_1075; // @[Mux.scala 19:72:@1893.4]
  assign _T_1186 = _T_1185 | _T_1077; // @[Mux.scala 19:72:@1894.4]
  assign _T_1187 = _T_1186 | _T_1079; // @[Mux.scala 19:72:@1895.4]
  assign _T_1188 = _T_1187 | _T_1081; // @[Mux.scala 19:72:@1896.4]
  assign _T_1189 = _T_1188 | _T_1083; // @[Mux.scala 19:72:@1897.4]
  assign _T_1190 = _T_1189 | _T_1085; // @[Mux.scala 19:72:@1898.4]
  assign _T_1191 = _T_1190 | _T_1087; // @[Mux.scala 19:72:@1899.4]
  assign _T_1192 = _T_1191 | _T_1089; // @[Mux.scala 19:72:@1900.4]
  assign _T_1193 = _T_1192 | _T_1091; // @[Mux.scala 19:72:@1901.4]
  assign _T_1194 = _T_1193 | _T_1093; // @[Mux.scala 19:72:@1902.4]
  assign _T_1195 = _T_1194 | _T_1095; // @[Mux.scala 19:72:@1903.4]
  assign _T_1196 = _T_1195 | _T_1097; // @[Mux.scala 19:72:@1904.4]
  assign _T_1197 = _T_1196 | _T_1099; // @[Mux.scala 19:72:@1905.4]
  assign _T_1198 = _T_1197 | _T_1101; // @[Mux.scala 19:72:@1906.4]
  assign _T_1199 = _T_1198 | _T_1103; // @[Mux.scala 19:72:@1907.4]
  assign _T_1200 = _T_1199 | _T_1105; // @[Mux.scala 19:72:@1908.4]
  assign _T_1201 = _T_1200 | _T_1107; // @[Mux.scala 19:72:@1909.4]
  assign _T_1202 = _T_1201 | _T_1109; // @[Mux.scala 19:72:@1910.4]
  assign _T_1203 = _T_1202 | _T_1111; // @[Mux.scala 19:72:@1911.4]
  assign _T_1204 = _T_1203 | _T_1113; // @[Mux.scala 19:72:@1912.4]
  assign _T_1205 = _T_1204 | _T_1115; // @[Mux.scala 19:72:@1913.4]
  assign _T_1206 = _T_1205 | _T_1117; // @[Mux.scala 19:72:@1914.4]
  assign _T_1207 = _T_1206 | _T_1119; // @[Mux.scala 19:72:@1915.4]
  assign _T_1208 = _T_1207 | _T_1121; // @[Mux.scala 19:72:@1916.4]
  assign _T_1209 = _T_1208 | _T_1123; // @[Mux.scala 19:72:@1917.4]
  assign _T_1210 = _T_1209 | _T_1125; // @[Mux.scala 19:72:@1918.4]
  assign _T_1211 = _T_1210 | _T_1127; // @[Mux.scala 19:72:@1919.4]
  assign _T_1212 = _T_1211 | _T_1129; // @[Mux.scala 19:72:@1920.4]
  assign _T_1213 = _T_1212 | _T_1131; // @[Mux.scala 19:72:@1921.4]
  assign _T_1214 = _T_1213 | _T_1133; // @[Mux.scala 19:72:@1922.4]
  assign _T_1215 = _T_1214 | _T_1135; // @[Mux.scala 19:72:@1923.4]
  assign _T_1216 = _T_1215 | _T_1137; // @[Mux.scala 19:72:@1924.4]
  assign _T_1217 = _T_1216 | _T_1139; // @[Mux.scala 19:72:@1925.4]
  assign _T_1218 = _T_1217 | _T_1141; // @[Mux.scala 19:72:@1926.4]
  assign _T_1219 = _T_1218 | _T_1143; // @[Mux.scala 19:72:@1927.4]
  assign _T_1220 = _T_1219 | _T_1145; // @[Mux.scala 19:72:@1928.4]
  assign _T_1221 = _T_1220 | _T_1147; // @[Mux.scala 19:72:@1929.4]
  assign _T_1222 = _T_1221 | _T_1149; // @[Mux.scala 19:72:@1930.4]
  assign _T_1223 = _T_1222 | _T_1151; // @[Mux.scala 19:72:@1931.4]
  assign _T_1224 = _T_1223 | _T_1153; // @[Mux.scala 19:72:@1932.4]
  assign _T_1225 = _T_1224 | _T_1155; // @[Mux.scala 19:72:@1933.4]
  assign _T_1226 = _T_1225 | _T_1157; // @[Mux.scala 19:72:@1934.4]
  assign _T_1227 = _T_1226 | _T_1159; // @[Mux.scala 19:72:@1935.4]
  assign _T_1228 = _T_1227 | _T_1161; // @[Mux.scala 19:72:@1936.4]
  assign _T_1229 = _T_1228 | _T_1163; // @[Mux.scala 19:72:@1937.4]
  assign _T_1230 = _T_1229 | _T_1165; // @[Mux.scala 19:72:@1938.4]
  assign _T_1231 = _T_1230 | _T_1167; // @[Mux.scala 19:72:@1939.4]
  assign predict_0_h_count = _T_1231 | _T_1169; // @[Mux.scala 19:72:@1940.4]
  assign _T_1236 = if_pc_0[9:0]; // @[BTB.scala 110:54:@1945.4]
  assign predict_0_gshxor = gb_history ^ _T_1236; // @[BTB.scala 110:44:@1946.4]
  assign _T_1240 = gb_history[8:0]; // @[BTB.scala 113:42:@1952.4]
  assign predict_0_gshare = bht__T_1239_data; // @[BTB.scala 98:21:@1087.4 BTB.scala 112:25:@1951.4]
  assign _T_1241 = predict_0_gshare[1]; // @[BTB.scala 47:40:@1953.4]
  assign _T_1242 = predict_0_h_count[1]; // @[BTB.scala 47:52:@1954.4]
  assign predict_0_select = arb__T_1238_data; // @[BTB.scala 98:21:@1087.4 BTB.scala 111:25:@1949.4]
  assign _T_1243 = predict_0_select ? _T_1241 : _T_1242; // @[BTB.scala 47:25:@1955.4]
  assign predict_0_history = {_T_1240,_T_1243}; // @[Cat.scala 30:58:@1956.4]
  assign _T_1246 = predict_0_lookup != 64'h0; // @[BTB.scala 40:28:@1958.4]
  assign _T_1250 = predict_0_bj_type != 2'h2; // @[BTB.scala 49:42:@1961.4]
  assign _T_1254 = _T_1250 | _T_1243; // @[BTB.scala 49:63:@1965.4]
  assign _T_1255 = _T_1246 & _T_1254; // @[BTB.scala 49:30:@1966.4]
  assign _T_1260 = predict_0_bj_type == 2'h1; // @[BTB.scala 119:54:@1973.4]
  assign _T_1270 = _T_1255 ? predict_0_jump_tgt : predict_0_cont_tgt; // @[BTB.scala 120:34:@1981.4]
  assign _T_1275 = btb_pc_0 == _T_178; // @[BTB.scala 105:47:@1987.4]
  assign _T_1276 = btb_pc_1 == _T_178; // @[BTB.scala 105:47:@1988.4]
  assign _T_1277 = btb_pc_2 == _T_178; // @[BTB.scala 105:47:@1989.4]
  assign _T_1278 = btb_pc_3 == _T_178; // @[BTB.scala 105:47:@1990.4]
  assign _T_1279 = btb_pc_4 == _T_178; // @[BTB.scala 105:47:@1991.4]
  assign _T_1280 = btb_pc_5 == _T_178; // @[BTB.scala 105:47:@1992.4]
  assign _T_1281 = btb_pc_6 == _T_178; // @[BTB.scala 105:47:@1993.4]
  assign _T_1282 = btb_pc_7 == _T_178; // @[BTB.scala 105:47:@1994.4]
  assign _T_1283 = btb_pc_8 == _T_178; // @[BTB.scala 105:47:@1995.4]
  assign _T_1284 = btb_pc_9 == _T_178; // @[BTB.scala 105:47:@1996.4]
  assign _T_1285 = btb_pc_10 == _T_178; // @[BTB.scala 105:47:@1997.4]
  assign _T_1286 = btb_pc_11 == _T_178; // @[BTB.scala 105:47:@1998.4]
  assign _T_1287 = btb_pc_12 == _T_178; // @[BTB.scala 105:47:@1999.4]
  assign _T_1288 = btb_pc_13 == _T_178; // @[BTB.scala 105:47:@2000.4]
  assign _T_1289 = btb_pc_14 == _T_178; // @[BTB.scala 105:47:@2001.4]
  assign _T_1290 = btb_pc_15 == _T_178; // @[BTB.scala 105:47:@2002.4]
  assign _T_1291 = btb_pc_16 == _T_178; // @[BTB.scala 105:47:@2003.4]
  assign _T_1292 = btb_pc_17 == _T_178; // @[BTB.scala 105:47:@2004.4]
  assign _T_1293 = btb_pc_18 == _T_178; // @[BTB.scala 105:47:@2005.4]
  assign _T_1294 = btb_pc_19 == _T_178; // @[BTB.scala 105:47:@2006.4]
  assign _T_1295 = btb_pc_20 == _T_178; // @[BTB.scala 105:47:@2007.4]
  assign _T_1296 = btb_pc_21 == _T_178; // @[BTB.scala 105:47:@2008.4]
  assign _T_1297 = btb_pc_22 == _T_178; // @[BTB.scala 105:47:@2009.4]
  assign _T_1298 = btb_pc_23 == _T_178; // @[BTB.scala 105:47:@2010.4]
  assign _T_1299 = btb_pc_24 == _T_178; // @[BTB.scala 105:47:@2011.4]
  assign _T_1300 = btb_pc_25 == _T_178; // @[BTB.scala 105:47:@2012.4]
  assign _T_1301 = btb_pc_26 == _T_178; // @[BTB.scala 105:47:@2013.4]
  assign _T_1302 = btb_pc_27 == _T_178; // @[BTB.scala 105:47:@2014.4]
  assign _T_1303 = btb_pc_28 == _T_178; // @[BTB.scala 105:47:@2015.4]
  assign _T_1304 = btb_pc_29 == _T_178; // @[BTB.scala 105:47:@2016.4]
  assign _T_1305 = btb_pc_30 == _T_178; // @[BTB.scala 105:47:@2017.4]
  assign _T_1306 = btb_pc_31 == _T_178; // @[BTB.scala 105:47:@2018.4]
  assign _T_1307 = btb_pc_32 == _T_178; // @[BTB.scala 105:47:@2019.4]
  assign _T_1308 = btb_pc_33 == _T_178; // @[BTB.scala 105:47:@2020.4]
  assign _T_1309 = btb_pc_34 == _T_178; // @[BTB.scala 105:47:@2021.4]
  assign _T_1310 = btb_pc_35 == _T_178; // @[BTB.scala 105:47:@2022.4]
  assign _T_1311 = btb_pc_36 == _T_178; // @[BTB.scala 105:47:@2023.4]
  assign _T_1312 = btb_pc_37 == _T_178; // @[BTB.scala 105:47:@2024.4]
  assign _T_1313 = btb_pc_38 == _T_178; // @[BTB.scala 105:47:@2025.4]
  assign _T_1314 = btb_pc_39 == _T_178; // @[BTB.scala 105:47:@2026.4]
  assign _T_1315 = btb_pc_40 == _T_178; // @[BTB.scala 105:47:@2027.4]
  assign _T_1316 = btb_pc_41 == _T_178; // @[BTB.scala 105:47:@2028.4]
  assign _T_1317 = btb_pc_42 == _T_178; // @[BTB.scala 105:47:@2029.4]
  assign _T_1318 = btb_pc_43 == _T_178; // @[BTB.scala 105:47:@2030.4]
  assign _T_1319 = btb_pc_44 == _T_178; // @[BTB.scala 105:47:@2031.4]
  assign _T_1320 = btb_pc_45 == _T_178; // @[BTB.scala 105:47:@2032.4]
  assign _T_1321 = btb_pc_46 == _T_178; // @[BTB.scala 105:47:@2033.4]
  assign _T_1322 = btb_pc_47 == _T_178; // @[BTB.scala 105:47:@2034.4]
  assign _T_1323 = btb_pc_48 == _T_178; // @[BTB.scala 105:47:@2035.4]
  assign _T_1324 = btb_pc_49 == _T_178; // @[BTB.scala 105:47:@2036.4]
  assign _T_1325 = btb_pc_50 == _T_178; // @[BTB.scala 105:47:@2037.4]
  assign _T_1326 = btb_pc_51 == _T_178; // @[BTB.scala 105:47:@2038.4]
  assign _T_1327 = btb_pc_52 == _T_178; // @[BTB.scala 105:47:@2039.4]
  assign _T_1328 = btb_pc_53 == _T_178; // @[BTB.scala 105:47:@2040.4]
  assign _T_1329 = btb_pc_54 == _T_178; // @[BTB.scala 105:47:@2041.4]
  assign _T_1330 = btb_pc_55 == _T_178; // @[BTB.scala 105:47:@2042.4]
  assign _T_1331 = btb_pc_56 == _T_178; // @[BTB.scala 105:47:@2043.4]
  assign _T_1332 = btb_pc_57 == _T_178; // @[BTB.scala 105:47:@2044.4]
  assign _T_1333 = btb_pc_58 == _T_178; // @[BTB.scala 105:47:@2045.4]
  assign _T_1334 = btb_pc_59 == _T_178; // @[BTB.scala 105:47:@2046.4]
  assign _T_1335 = btb_pc_60 == _T_178; // @[BTB.scala 105:47:@2047.4]
  assign _T_1336 = btb_pc_61 == _T_178; // @[BTB.scala 105:47:@2048.4]
  assign _T_1337 = btb_pc_62 == _T_178; // @[BTB.scala 105:47:@2049.4]
  assign _T_1338 = btb_pc_63 == _T_178; // @[BTB.scala 105:47:@2050.4]
  assign _T_1415 = {_T_1282,_T_1281,_T_1280,_T_1279,_T_1278,_T_1277,_T_1276,_T_1275}; // @[BTB.scala 105:62:@2122.4]
  assign _T_1423 = {_T_1290,_T_1289,_T_1288,_T_1287,_T_1286,_T_1285,_T_1284,_T_1283,_T_1415}; // @[BTB.scala 105:62:@2130.4]
  assign _T_1430 = {_T_1298,_T_1297,_T_1296,_T_1295,_T_1294,_T_1293,_T_1292,_T_1291}; // @[BTB.scala 105:62:@2137.4]
  assign _T_1439 = {_T_1306,_T_1305,_T_1304,_T_1303,_T_1302,_T_1301,_T_1300,_T_1299,_T_1430,_T_1423}; // @[BTB.scala 105:62:@2146.4]
  assign _T_1446 = {_T_1314,_T_1313,_T_1312,_T_1311,_T_1310,_T_1309,_T_1308,_T_1307}; // @[BTB.scala 105:62:@2153.4]
  assign _T_1454 = {_T_1322,_T_1321,_T_1320,_T_1319,_T_1318,_T_1317,_T_1316,_T_1315,_T_1446}; // @[BTB.scala 105:62:@2161.4]
  assign _T_1461 = {_T_1330,_T_1329,_T_1328,_T_1327,_T_1326,_T_1325,_T_1324,_T_1323}; // @[BTB.scala 105:62:@2168.4]
  assign _T_1470 = {_T_1338,_T_1337,_T_1336,_T_1335,_T_1334,_T_1333,_T_1332,_T_1331,_T_1461,_T_1454}; // @[BTB.scala 105:62:@2177.4]
  assign _T_1471 = {_T_1470,_T_1439}; // @[BTB.scala 105:62:@2178.4]
  assign predict_1_lookup = _T_1471 & _T_457; // @[BTB.scala 105:69:@2242.4]
  assign _T_1536 = predict_1_lookup[0]; // @[Mux.scala 21:36:@2244.4]
  assign _T_1537 = predict_1_lookup[1]; // @[Mux.scala 21:36:@2245.4]
  assign _T_1538 = predict_1_lookup[2]; // @[Mux.scala 21:36:@2246.4]
  assign _T_1539 = predict_1_lookup[3]; // @[Mux.scala 21:36:@2247.4]
  assign _T_1540 = predict_1_lookup[4]; // @[Mux.scala 21:36:@2248.4]
  assign _T_1541 = predict_1_lookup[5]; // @[Mux.scala 21:36:@2249.4]
  assign _T_1542 = predict_1_lookup[6]; // @[Mux.scala 21:36:@2250.4]
  assign _T_1543 = predict_1_lookup[7]; // @[Mux.scala 21:36:@2251.4]
  assign _T_1544 = predict_1_lookup[8]; // @[Mux.scala 21:36:@2252.4]
  assign _T_1545 = predict_1_lookup[9]; // @[Mux.scala 21:36:@2253.4]
  assign _T_1546 = predict_1_lookup[10]; // @[Mux.scala 21:36:@2254.4]
  assign _T_1547 = predict_1_lookup[11]; // @[Mux.scala 21:36:@2255.4]
  assign _T_1548 = predict_1_lookup[12]; // @[Mux.scala 21:36:@2256.4]
  assign _T_1549 = predict_1_lookup[13]; // @[Mux.scala 21:36:@2257.4]
  assign _T_1550 = predict_1_lookup[14]; // @[Mux.scala 21:36:@2258.4]
  assign _T_1551 = predict_1_lookup[15]; // @[Mux.scala 21:36:@2259.4]
  assign _T_1552 = predict_1_lookup[16]; // @[Mux.scala 21:36:@2260.4]
  assign _T_1553 = predict_1_lookup[17]; // @[Mux.scala 21:36:@2261.4]
  assign _T_1554 = predict_1_lookup[18]; // @[Mux.scala 21:36:@2262.4]
  assign _T_1555 = predict_1_lookup[19]; // @[Mux.scala 21:36:@2263.4]
  assign _T_1556 = predict_1_lookup[20]; // @[Mux.scala 21:36:@2264.4]
  assign _T_1557 = predict_1_lookup[21]; // @[Mux.scala 21:36:@2265.4]
  assign _T_1558 = predict_1_lookup[22]; // @[Mux.scala 21:36:@2266.4]
  assign _T_1559 = predict_1_lookup[23]; // @[Mux.scala 21:36:@2267.4]
  assign _T_1560 = predict_1_lookup[24]; // @[Mux.scala 21:36:@2268.4]
  assign _T_1561 = predict_1_lookup[25]; // @[Mux.scala 21:36:@2269.4]
  assign _T_1562 = predict_1_lookup[26]; // @[Mux.scala 21:36:@2270.4]
  assign _T_1563 = predict_1_lookup[27]; // @[Mux.scala 21:36:@2271.4]
  assign _T_1564 = predict_1_lookup[28]; // @[Mux.scala 21:36:@2272.4]
  assign _T_1565 = predict_1_lookup[29]; // @[Mux.scala 21:36:@2273.4]
  assign _T_1566 = predict_1_lookup[30]; // @[Mux.scala 21:36:@2274.4]
  assign _T_1567 = predict_1_lookup[31]; // @[Mux.scala 21:36:@2275.4]
  assign _T_1568 = predict_1_lookup[32]; // @[Mux.scala 21:36:@2276.4]
  assign _T_1569 = predict_1_lookup[33]; // @[Mux.scala 21:36:@2277.4]
  assign _T_1570 = predict_1_lookup[34]; // @[Mux.scala 21:36:@2278.4]
  assign _T_1571 = predict_1_lookup[35]; // @[Mux.scala 21:36:@2279.4]
  assign _T_1572 = predict_1_lookup[36]; // @[Mux.scala 21:36:@2280.4]
  assign _T_1573 = predict_1_lookup[37]; // @[Mux.scala 21:36:@2281.4]
  assign _T_1574 = predict_1_lookup[38]; // @[Mux.scala 21:36:@2282.4]
  assign _T_1575 = predict_1_lookup[39]; // @[Mux.scala 21:36:@2283.4]
  assign _T_1576 = predict_1_lookup[40]; // @[Mux.scala 21:36:@2284.4]
  assign _T_1577 = predict_1_lookup[41]; // @[Mux.scala 21:36:@2285.4]
  assign _T_1578 = predict_1_lookup[42]; // @[Mux.scala 21:36:@2286.4]
  assign _T_1579 = predict_1_lookup[43]; // @[Mux.scala 21:36:@2287.4]
  assign _T_1580 = predict_1_lookup[44]; // @[Mux.scala 21:36:@2288.4]
  assign _T_1581 = predict_1_lookup[45]; // @[Mux.scala 21:36:@2289.4]
  assign _T_1582 = predict_1_lookup[46]; // @[Mux.scala 21:36:@2290.4]
  assign _T_1583 = predict_1_lookup[47]; // @[Mux.scala 21:36:@2291.4]
  assign _T_1584 = predict_1_lookup[48]; // @[Mux.scala 21:36:@2292.4]
  assign _T_1585 = predict_1_lookup[49]; // @[Mux.scala 21:36:@2293.4]
  assign _T_1586 = predict_1_lookup[50]; // @[Mux.scala 21:36:@2294.4]
  assign _T_1587 = predict_1_lookup[51]; // @[Mux.scala 21:36:@2295.4]
  assign _T_1588 = predict_1_lookup[52]; // @[Mux.scala 21:36:@2296.4]
  assign _T_1589 = predict_1_lookup[53]; // @[Mux.scala 21:36:@2297.4]
  assign _T_1590 = predict_1_lookup[54]; // @[Mux.scala 21:36:@2298.4]
  assign _T_1591 = predict_1_lookup[55]; // @[Mux.scala 21:36:@2299.4]
  assign _T_1592 = predict_1_lookup[56]; // @[Mux.scala 21:36:@2300.4]
  assign _T_1593 = predict_1_lookup[57]; // @[Mux.scala 21:36:@2301.4]
  assign _T_1594 = predict_1_lookup[58]; // @[Mux.scala 21:36:@2302.4]
  assign _T_1595 = predict_1_lookup[59]; // @[Mux.scala 21:36:@2303.4]
  assign _T_1596 = predict_1_lookup[60]; // @[Mux.scala 21:36:@2304.4]
  assign _T_1597 = predict_1_lookup[61]; // @[Mux.scala 21:36:@2305.4]
  assign _T_1598 = predict_1_lookup[62]; // @[Mux.scala 21:36:@2306.4]
  assign _T_1599 = predict_1_lookup[63]; // @[Mux.scala 21:36:@2307.4]
  assign _T_1602 = _T_1536 ? btb_tgt_0 : 30'h0; // @[Mux.scala 19:72:@2308.4]
  assign _T_1604 = _T_1537 ? btb_tgt_1 : 30'h0; // @[Mux.scala 19:72:@2309.4]
  assign _T_1606 = _T_1538 ? btb_tgt_2 : 30'h0; // @[Mux.scala 19:72:@2310.4]
  assign _T_1608 = _T_1539 ? btb_tgt_3 : 30'h0; // @[Mux.scala 19:72:@2311.4]
  assign _T_1610 = _T_1540 ? btb_tgt_4 : 30'h0; // @[Mux.scala 19:72:@2312.4]
  assign _T_1612 = _T_1541 ? btb_tgt_5 : 30'h0; // @[Mux.scala 19:72:@2313.4]
  assign _T_1614 = _T_1542 ? btb_tgt_6 : 30'h0; // @[Mux.scala 19:72:@2314.4]
  assign _T_1616 = _T_1543 ? btb_tgt_7 : 30'h0; // @[Mux.scala 19:72:@2315.4]
  assign _T_1618 = _T_1544 ? btb_tgt_8 : 30'h0; // @[Mux.scala 19:72:@2316.4]
  assign _T_1620 = _T_1545 ? btb_tgt_9 : 30'h0; // @[Mux.scala 19:72:@2317.4]
  assign _T_1622 = _T_1546 ? btb_tgt_10 : 30'h0; // @[Mux.scala 19:72:@2318.4]
  assign _T_1624 = _T_1547 ? btb_tgt_11 : 30'h0; // @[Mux.scala 19:72:@2319.4]
  assign _T_1626 = _T_1548 ? btb_tgt_12 : 30'h0; // @[Mux.scala 19:72:@2320.4]
  assign _T_1628 = _T_1549 ? btb_tgt_13 : 30'h0; // @[Mux.scala 19:72:@2321.4]
  assign _T_1630 = _T_1550 ? btb_tgt_14 : 30'h0; // @[Mux.scala 19:72:@2322.4]
  assign _T_1632 = _T_1551 ? btb_tgt_15 : 30'h0; // @[Mux.scala 19:72:@2323.4]
  assign _T_1634 = _T_1552 ? btb_tgt_16 : 30'h0; // @[Mux.scala 19:72:@2324.4]
  assign _T_1636 = _T_1553 ? btb_tgt_17 : 30'h0; // @[Mux.scala 19:72:@2325.4]
  assign _T_1638 = _T_1554 ? btb_tgt_18 : 30'h0; // @[Mux.scala 19:72:@2326.4]
  assign _T_1640 = _T_1555 ? btb_tgt_19 : 30'h0; // @[Mux.scala 19:72:@2327.4]
  assign _T_1642 = _T_1556 ? btb_tgt_20 : 30'h0; // @[Mux.scala 19:72:@2328.4]
  assign _T_1644 = _T_1557 ? btb_tgt_21 : 30'h0; // @[Mux.scala 19:72:@2329.4]
  assign _T_1646 = _T_1558 ? btb_tgt_22 : 30'h0; // @[Mux.scala 19:72:@2330.4]
  assign _T_1648 = _T_1559 ? btb_tgt_23 : 30'h0; // @[Mux.scala 19:72:@2331.4]
  assign _T_1650 = _T_1560 ? btb_tgt_24 : 30'h0; // @[Mux.scala 19:72:@2332.4]
  assign _T_1652 = _T_1561 ? btb_tgt_25 : 30'h0; // @[Mux.scala 19:72:@2333.4]
  assign _T_1654 = _T_1562 ? btb_tgt_26 : 30'h0; // @[Mux.scala 19:72:@2334.4]
  assign _T_1656 = _T_1563 ? btb_tgt_27 : 30'h0; // @[Mux.scala 19:72:@2335.4]
  assign _T_1658 = _T_1564 ? btb_tgt_28 : 30'h0; // @[Mux.scala 19:72:@2336.4]
  assign _T_1660 = _T_1565 ? btb_tgt_29 : 30'h0; // @[Mux.scala 19:72:@2337.4]
  assign _T_1662 = _T_1566 ? btb_tgt_30 : 30'h0; // @[Mux.scala 19:72:@2338.4]
  assign _T_1664 = _T_1567 ? btb_tgt_31 : 30'h0; // @[Mux.scala 19:72:@2339.4]
  assign _T_1666 = _T_1568 ? btb_tgt_32 : 30'h0; // @[Mux.scala 19:72:@2340.4]
  assign _T_1668 = _T_1569 ? btb_tgt_33 : 30'h0; // @[Mux.scala 19:72:@2341.4]
  assign _T_1670 = _T_1570 ? btb_tgt_34 : 30'h0; // @[Mux.scala 19:72:@2342.4]
  assign _T_1672 = _T_1571 ? btb_tgt_35 : 30'h0; // @[Mux.scala 19:72:@2343.4]
  assign _T_1674 = _T_1572 ? btb_tgt_36 : 30'h0; // @[Mux.scala 19:72:@2344.4]
  assign _T_1676 = _T_1573 ? btb_tgt_37 : 30'h0; // @[Mux.scala 19:72:@2345.4]
  assign _T_1678 = _T_1574 ? btb_tgt_38 : 30'h0; // @[Mux.scala 19:72:@2346.4]
  assign _T_1680 = _T_1575 ? btb_tgt_39 : 30'h0; // @[Mux.scala 19:72:@2347.4]
  assign _T_1682 = _T_1576 ? btb_tgt_40 : 30'h0; // @[Mux.scala 19:72:@2348.4]
  assign _T_1684 = _T_1577 ? btb_tgt_41 : 30'h0; // @[Mux.scala 19:72:@2349.4]
  assign _T_1686 = _T_1578 ? btb_tgt_42 : 30'h0; // @[Mux.scala 19:72:@2350.4]
  assign _T_1688 = _T_1579 ? btb_tgt_43 : 30'h0; // @[Mux.scala 19:72:@2351.4]
  assign _T_1690 = _T_1580 ? btb_tgt_44 : 30'h0; // @[Mux.scala 19:72:@2352.4]
  assign _T_1692 = _T_1581 ? btb_tgt_45 : 30'h0; // @[Mux.scala 19:72:@2353.4]
  assign _T_1694 = _T_1582 ? btb_tgt_46 : 30'h0; // @[Mux.scala 19:72:@2354.4]
  assign _T_1696 = _T_1583 ? btb_tgt_47 : 30'h0; // @[Mux.scala 19:72:@2355.4]
  assign _T_1698 = _T_1584 ? btb_tgt_48 : 30'h0; // @[Mux.scala 19:72:@2356.4]
  assign _T_1700 = _T_1585 ? btb_tgt_49 : 30'h0; // @[Mux.scala 19:72:@2357.4]
  assign _T_1702 = _T_1586 ? btb_tgt_50 : 30'h0; // @[Mux.scala 19:72:@2358.4]
  assign _T_1704 = _T_1587 ? btb_tgt_51 : 30'h0; // @[Mux.scala 19:72:@2359.4]
  assign _T_1706 = _T_1588 ? btb_tgt_52 : 30'h0; // @[Mux.scala 19:72:@2360.4]
  assign _T_1708 = _T_1589 ? btb_tgt_53 : 30'h0; // @[Mux.scala 19:72:@2361.4]
  assign _T_1710 = _T_1590 ? btb_tgt_54 : 30'h0; // @[Mux.scala 19:72:@2362.4]
  assign _T_1712 = _T_1591 ? btb_tgt_55 : 30'h0; // @[Mux.scala 19:72:@2363.4]
  assign _T_1714 = _T_1592 ? btb_tgt_56 : 30'h0; // @[Mux.scala 19:72:@2364.4]
  assign _T_1716 = _T_1593 ? btb_tgt_57 : 30'h0; // @[Mux.scala 19:72:@2365.4]
  assign _T_1718 = _T_1594 ? btb_tgt_58 : 30'h0; // @[Mux.scala 19:72:@2366.4]
  assign _T_1720 = _T_1595 ? btb_tgt_59 : 30'h0; // @[Mux.scala 19:72:@2367.4]
  assign _T_1722 = _T_1596 ? btb_tgt_60 : 30'h0; // @[Mux.scala 19:72:@2368.4]
  assign _T_1724 = _T_1597 ? btb_tgt_61 : 30'h0; // @[Mux.scala 19:72:@2369.4]
  assign _T_1726 = _T_1598 ? btb_tgt_62 : 30'h0; // @[Mux.scala 19:72:@2370.4]
  assign _T_1728 = _T_1599 ? btb_tgt_63 : 30'h0; // @[Mux.scala 19:72:@2371.4]
  assign _T_1729 = _T_1602 | _T_1604; // @[Mux.scala 19:72:@2372.4]
  assign _T_1730 = _T_1729 | _T_1606; // @[Mux.scala 19:72:@2373.4]
  assign _T_1731 = _T_1730 | _T_1608; // @[Mux.scala 19:72:@2374.4]
  assign _T_1732 = _T_1731 | _T_1610; // @[Mux.scala 19:72:@2375.4]
  assign _T_1733 = _T_1732 | _T_1612; // @[Mux.scala 19:72:@2376.4]
  assign _T_1734 = _T_1733 | _T_1614; // @[Mux.scala 19:72:@2377.4]
  assign _T_1735 = _T_1734 | _T_1616; // @[Mux.scala 19:72:@2378.4]
  assign _T_1736 = _T_1735 | _T_1618; // @[Mux.scala 19:72:@2379.4]
  assign _T_1737 = _T_1736 | _T_1620; // @[Mux.scala 19:72:@2380.4]
  assign _T_1738 = _T_1737 | _T_1622; // @[Mux.scala 19:72:@2381.4]
  assign _T_1739 = _T_1738 | _T_1624; // @[Mux.scala 19:72:@2382.4]
  assign _T_1740 = _T_1739 | _T_1626; // @[Mux.scala 19:72:@2383.4]
  assign _T_1741 = _T_1740 | _T_1628; // @[Mux.scala 19:72:@2384.4]
  assign _T_1742 = _T_1741 | _T_1630; // @[Mux.scala 19:72:@2385.4]
  assign _T_1743 = _T_1742 | _T_1632; // @[Mux.scala 19:72:@2386.4]
  assign _T_1744 = _T_1743 | _T_1634; // @[Mux.scala 19:72:@2387.4]
  assign _T_1745 = _T_1744 | _T_1636; // @[Mux.scala 19:72:@2388.4]
  assign _T_1746 = _T_1745 | _T_1638; // @[Mux.scala 19:72:@2389.4]
  assign _T_1747 = _T_1746 | _T_1640; // @[Mux.scala 19:72:@2390.4]
  assign _T_1748 = _T_1747 | _T_1642; // @[Mux.scala 19:72:@2391.4]
  assign _T_1749 = _T_1748 | _T_1644; // @[Mux.scala 19:72:@2392.4]
  assign _T_1750 = _T_1749 | _T_1646; // @[Mux.scala 19:72:@2393.4]
  assign _T_1751 = _T_1750 | _T_1648; // @[Mux.scala 19:72:@2394.4]
  assign _T_1752 = _T_1751 | _T_1650; // @[Mux.scala 19:72:@2395.4]
  assign _T_1753 = _T_1752 | _T_1652; // @[Mux.scala 19:72:@2396.4]
  assign _T_1754 = _T_1753 | _T_1654; // @[Mux.scala 19:72:@2397.4]
  assign _T_1755 = _T_1754 | _T_1656; // @[Mux.scala 19:72:@2398.4]
  assign _T_1756 = _T_1755 | _T_1658; // @[Mux.scala 19:72:@2399.4]
  assign _T_1757 = _T_1756 | _T_1660; // @[Mux.scala 19:72:@2400.4]
  assign _T_1758 = _T_1757 | _T_1662; // @[Mux.scala 19:72:@2401.4]
  assign _T_1759 = _T_1758 | _T_1664; // @[Mux.scala 19:72:@2402.4]
  assign _T_1760 = _T_1759 | _T_1666; // @[Mux.scala 19:72:@2403.4]
  assign _T_1761 = _T_1760 | _T_1668; // @[Mux.scala 19:72:@2404.4]
  assign _T_1762 = _T_1761 | _T_1670; // @[Mux.scala 19:72:@2405.4]
  assign _T_1763 = _T_1762 | _T_1672; // @[Mux.scala 19:72:@2406.4]
  assign _T_1764 = _T_1763 | _T_1674; // @[Mux.scala 19:72:@2407.4]
  assign _T_1765 = _T_1764 | _T_1676; // @[Mux.scala 19:72:@2408.4]
  assign _T_1766 = _T_1765 | _T_1678; // @[Mux.scala 19:72:@2409.4]
  assign _T_1767 = _T_1766 | _T_1680; // @[Mux.scala 19:72:@2410.4]
  assign _T_1768 = _T_1767 | _T_1682; // @[Mux.scala 19:72:@2411.4]
  assign _T_1769 = _T_1768 | _T_1684; // @[Mux.scala 19:72:@2412.4]
  assign _T_1770 = _T_1769 | _T_1686; // @[Mux.scala 19:72:@2413.4]
  assign _T_1771 = _T_1770 | _T_1688; // @[Mux.scala 19:72:@2414.4]
  assign _T_1772 = _T_1771 | _T_1690; // @[Mux.scala 19:72:@2415.4]
  assign _T_1773 = _T_1772 | _T_1692; // @[Mux.scala 19:72:@2416.4]
  assign _T_1774 = _T_1773 | _T_1694; // @[Mux.scala 19:72:@2417.4]
  assign _T_1775 = _T_1774 | _T_1696; // @[Mux.scala 19:72:@2418.4]
  assign _T_1776 = _T_1775 | _T_1698; // @[Mux.scala 19:72:@2419.4]
  assign _T_1777 = _T_1776 | _T_1700; // @[Mux.scala 19:72:@2420.4]
  assign _T_1778 = _T_1777 | _T_1702; // @[Mux.scala 19:72:@2421.4]
  assign _T_1779 = _T_1778 | _T_1704; // @[Mux.scala 19:72:@2422.4]
  assign _T_1780 = _T_1779 | _T_1706; // @[Mux.scala 19:72:@2423.4]
  assign _T_1781 = _T_1780 | _T_1708; // @[Mux.scala 19:72:@2424.4]
  assign _T_1782 = _T_1781 | _T_1710; // @[Mux.scala 19:72:@2425.4]
  assign _T_1783 = _T_1782 | _T_1712; // @[Mux.scala 19:72:@2426.4]
  assign _T_1784 = _T_1783 | _T_1714; // @[Mux.scala 19:72:@2427.4]
  assign _T_1785 = _T_1784 | _T_1716; // @[Mux.scala 19:72:@2428.4]
  assign _T_1786 = _T_1785 | _T_1718; // @[Mux.scala 19:72:@2429.4]
  assign _T_1787 = _T_1786 | _T_1720; // @[Mux.scala 19:72:@2430.4]
  assign _T_1788 = _T_1787 | _T_1722; // @[Mux.scala 19:72:@2431.4]
  assign _T_1789 = _T_1788 | _T_1724; // @[Mux.scala 19:72:@2432.4]
  assign _T_1790 = _T_1789 | _T_1726; // @[Mux.scala 19:72:@2433.4]
  assign _T_1791 = _T_1790 | _T_1728; // @[Mux.scala 19:72:@2434.4]
  assign predict_1_jump_tgt = {_T_1791,2'h0}; // @[Cat.scala 30:58:@2437.4]
  assign _T_1862 = _T_1536 ? btb_bj_type_0 : 2'h0; // @[Mux.scala 19:72:@2503.4]
  assign _T_1864 = _T_1537 ? btb_bj_type_1 : 2'h0; // @[Mux.scala 19:72:@2504.4]
  assign _T_1866 = _T_1538 ? btb_bj_type_2 : 2'h0; // @[Mux.scala 19:72:@2505.4]
  assign _T_1868 = _T_1539 ? btb_bj_type_3 : 2'h0; // @[Mux.scala 19:72:@2506.4]
  assign _T_1870 = _T_1540 ? btb_bj_type_4 : 2'h0; // @[Mux.scala 19:72:@2507.4]
  assign _T_1872 = _T_1541 ? btb_bj_type_5 : 2'h0; // @[Mux.scala 19:72:@2508.4]
  assign _T_1874 = _T_1542 ? btb_bj_type_6 : 2'h0; // @[Mux.scala 19:72:@2509.4]
  assign _T_1876 = _T_1543 ? btb_bj_type_7 : 2'h0; // @[Mux.scala 19:72:@2510.4]
  assign _T_1878 = _T_1544 ? btb_bj_type_8 : 2'h0; // @[Mux.scala 19:72:@2511.4]
  assign _T_1880 = _T_1545 ? btb_bj_type_9 : 2'h0; // @[Mux.scala 19:72:@2512.4]
  assign _T_1882 = _T_1546 ? btb_bj_type_10 : 2'h0; // @[Mux.scala 19:72:@2513.4]
  assign _T_1884 = _T_1547 ? btb_bj_type_11 : 2'h0; // @[Mux.scala 19:72:@2514.4]
  assign _T_1886 = _T_1548 ? btb_bj_type_12 : 2'h0; // @[Mux.scala 19:72:@2515.4]
  assign _T_1888 = _T_1549 ? btb_bj_type_13 : 2'h0; // @[Mux.scala 19:72:@2516.4]
  assign _T_1890 = _T_1550 ? btb_bj_type_14 : 2'h0; // @[Mux.scala 19:72:@2517.4]
  assign _T_1892 = _T_1551 ? btb_bj_type_15 : 2'h0; // @[Mux.scala 19:72:@2518.4]
  assign _T_1894 = _T_1552 ? btb_bj_type_16 : 2'h0; // @[Mux.scala 19:72:@2519.4]
  assign _T_1896 = _T_1553 ? btb_bj_type_17 : 2'h0; // @[Mux.scala 19:72:@2520.4]
  assign _T_1898 = _T_1554 ? btb_bj_type_18 : 2'h0; // @[Mux.scala 19:72:@2521.4]
  assign _T_1900 = _T_1555 ? btb_bj_type_19 : 2'h0; // @[Mux.scala 19:72:@2522.4]
  assign _T_1902 = _T_1556 ? btb_bj_type_20 : 2'h0; // @[Mux.scala 19:72:@2523.4]
  assign _T_1904 = _T_1557 ? btb_bj_type_21 : 2'h0; // @[Mux.scala 19:72:@2524.4]
  assign _T_1906 = _T_1558 ? btb_bj_type_22 : 2'h0; // @[Mux.scala 19:72:@2525.4]
  assign _T_1908 = _T_1559 ? btb_bj_type_23 : 2'h0; // @[Mux.scala 19:72:@2526.4]
  assign _T_1910 = _T_1560 ? btb_bj_type_24 : 2'h0; // @[Mux.scala 19:72:@2527.4]
  assign _T_1912 = _T_1561 ? btb_bj_type_25 : 2'h0; // @[Mux.scala 19:72:@2528.4]
  assign _T_1914 = _T_1562 ? btb_bj_type_26 : 2'h0; // @[Mux.scala 19:72:@2529.4]
  assign _T_1916 = _T_1563 ? btb_bj_type_27 : 2'h0; // @[Mux.scala 19:72:@2530.4]
  assign _T_1918 = _T_1564 ? btb_bj_type_28 : 2'h0; // @[Mux.scala 19:72:@2531.4]
  assign _T_1920 = _T_1565 ? btb_bj_type_29 : 2'h0; // @[Mux.scala 19:72:@2532.4]
  assign _T_1922 = _T_1566 ? btb_bj_type_30 : 2'h0; // @[Mux.scala 19:72:@2533.4]
  assign _T_1924 = _T_1567 ? btb_bj_type_31 : 2'h0; // @[Mux.scala 19:72:@2534.4]
  assign _T_1926 = _T_1568 ? btb_bj_type_32 : 2'h0; // @[Mux.scala 19:72:@2535.4]
  assign _T_1928 = _T_1569 ? btb_bj_type_33 : 2'h0; // @[Mux.scala 19:72:@2536.4]
  assign _T_1930 = _T_1570 ? btb_bj_type_34 : 2'h0; // @[Mux.scala 19:72:@2537.4]
  assign _T_1932 = _T_1571 ? btb_bj_type_35 : 2'h0; // @[Mux.scala 19:72:@2538.4]
  assign _T_1934 = _T_1572 ? btb_bj_type_36 : 2'h0; // @[Mux.scala 19:72:@2539.4]
  assign _T_1936 = _T_1573 ? btb_bj_type_37 : 2'h0; // @[Mux.scala 19:72:@2540.4]
  assign _T_1938 = _T_1574 ? btb_bj_type_38 : 2'h0; // @[Mux.scala 19:72:@2541.4]
  assign _T_1940 = _T_1575 ? btb_bj_type_39 : 2'h0; // @[Mux.scala 19:72:@2542.4]
  assign _T_1942 = _T_1576 ? btb_bj_type_40 : 2'h0; // @[Mux.scala 19:72:@2543.4]
  assign _T_1944 = _T_1577 ? btb_bj_type_41 : 2'h0; // @[Mux.scala 19:72:@2544.4]
  assign _T_1946 = _T_1578 ? btb_bj_type_42 : 2'h0; // @[Mux.scala 19:72:@2545.4]
  assign _T_1948 = _T_1579 ? btb_bj_type_43 : 2'h0; // @[Mux.scala 19:72:@2546.4]
  assign _T_1950 = _T_1580 ? btb_bj_type_44 : 2'h0; // @[Mux.scala 19:72:@2547.4]
  assign _T_1952 = _T_1581 ? btb_bj_type_45 : 2'h0; // @[Mux.scala 19:72:@2548.4]
  assign _T_1954 = _T_1582 ? btb_bj_type_46 : 2'h0; // @[Mux.scala 19:72:@2549.4]
  assign _T_1956 = _T_1583 ? btb_bj_type_47 : 2'h0; // @[Mux.scala 19:72:@2550.4]
  assign _T_1958 = _T_1584 ? btb_bj_type_48 : 2'h0; // @[Mux.scala 19:72:@2551.4]
  assign _T_1960 = _T_1585 ? btb_bj_type_49 : 2'h0; // @[Mux.scala 19:72:@2552.4]
  assign _T_1962 = _T_1586 ? btb_bj_type_50 : 2'h0; // @[Mux.scala 19:72:@2553.4]
  assign _T_1964 = _T_1587 ? btb_bj_type_51 : 2'h0; // @[Mux.scala 19:72:@2554.4]
  assign _T_1966 = _T_1588 ? btb_bj_type_52 : 2'h0; // @[Mux.scala 19:72:@2555.4]
  assign _T_1968 = _T_1589 ? btb_bj_type_53 : 2'h0; // @[Mux.scala 19:72:@2556.4]
  assign _T_1970 = _T_1590 ? btb_bj_type_54 : 2'h0; // @[Mux.scala 19:72:@2557.4]
  assign _T_1972 = _T_1591 ? btb_bj_type_55 : 2'h0; // @[Mux.scala 19:72:@2558.4]
  assign _T_1974 = _T_1592 ? btb_bj_type_56 : 2'h0; // @[Mux.scala 19:72:@2559.4]
  assign _T_1976 = _T_1593 ? btb_bj_type_57 : 2'h0; // @[Mux.scala 19:72:@2560.4]
  assign _T_1978 = _T_1594 ? btb_bj_type_58 : 2'h0; // @[Mux.scala 19:72:@2561.4]
  assign _T_1980 = _T_1595 ? btb_bj_type_59 : 2'h0; // @[Mux.scala 19:72:@2562.4]
  assign _T_1982 = _T_1596 ? btb_bj_type_60 : 2'h0; // @[Mux.scala 19:72:@2563.4]
  assign _T_1984 = _T_1597 ? btb_bj_type_61 : 2'h0; // @[Mux.scala 19:72:@2564.4]
  assign _T_1986 = _T_1598 ? btb_bj_type_62 : 2'h0; // @[Mux.scala 19:72:@2565.4]
  assign _T_1988 = _T_1599 ? btb_bj_type_63 : 2'h0; // @[Mux.scala 19:72:@2566.4]
  assign _T_1989 = _T_1862 | _T_1864; // @[Mux.scala 19:72:@2567.4]
  assign _T_1990 = _T_1989 | _T_1866; // @[Mux.scala 19:72:@2568.4]
  assign _T_1991 = _T_1990 | _T_1868; // @[Mux.scala 19:72:@2569.4]
  assign _T_1992 = _T_1991 | _T_1870; // @[Mux.scala 19:72:@2570.4]
  assign _T_1993 = _T_1992 | _T_1872; // @[Mux.scala 19:72:@2571.4]
  assign _T_1994 = _T_1993 | _T_1874; // @[Mux.scala 19:72:@2572.4]
  assign _T_1995 = _T_1994 | _T_1876; // @[Mux.scala 19:72:@2573.4]
  assign _T_1996 = _T_1995 | _T_1878; // @[Mux.scala 19:72:@2574.4]
  assign _T_1997 = _T_1996 | _T_1880; // @[Mux.scala 19:72:@2575.4]
  assign _T_1998 = _T_1997 | _T_1882; // @[Mux.scala 19:72:@2576.4]
  assign _T_1999 = _T_1998 | _T_1884; // @[Mux.scala 19:72:@2577.4]
  assign _T_2000 = _T_1999 | _T_1886; // @[Mux.scala 19:72:@2578.4]
  assign _T_2001 = _T_2000 | _T_1888; // @[Mux.scala 19:72:@2579.4]
  assign _T_2002 = _T_2001 | _T_1890; // @[Mux.scala 19:72:@2580.4]
  assign _T_2003 = _T_2002 | _T_1892; // @[Mux.scala 19:72:@2581.4]
  assign _T_2004 = _T_2003 | _T_1894; // @[Mux.scala 19:72:@2582.4]
  assign _T_2005 = _T_2004 | _T_1896; // @[Mux.scala 19:72:@2583.4]
  assign _T_2006 = _T_2005 | _T_1898; // @[Mux.scala 19:72:@2584.4]
  assign _T_2007 = _T_2006 | _T_1900; // @[Mux.scala 19:72:@2585.4]
  assign _T_2008 = _T_2007 | _T_1902; // @[Mux.scala 19:72:@2586.4]
  assign _T_2009 = _T_2008 | _T_1904; // @[Mux.scala 19:72:@2587.4]
  assign _T_2010 = _T_2009 | _T_1906; // @[Mux.scala 19:72:@2588.4]
  assign _T_2011 = _T_2010 | _T_1908; // @[Mux.scala 19:72:@2589.4]
  assign _T_2012 = _T_2011 | _T_1910; // @[Mux.scala 19:72:@2590.4]
  assign _T_2013 = _T_2012 | _T_1912; // @[Mux.scala 19:72:@2591.4]
  assign _T_2014 = _T_2013 | _T_1914; // @[Mux.scala 19:72:@2592.4]
  assign _T_2015 = _T_2014 | _T_1916; // @[Mux.scala 19:72:@2593.4]
  assign _T_2016 = _T_2015 | _T_1918; // @[Mux.scala 19:72:@2594.4]
  assign _T_2017 = _T_2016 | _T_1920; // @[Mux.scala 19:72:@2595.4]
  assign _T_2018 = _T_2017 | _T_1922; // @[Mux.scala 19:72:@2596.4]
  assign _T_2019 = _T_2018 | _T_1924; // @[Mux.scala 19:72:@2597.4]
  assign _T_2020 = _T_2019 | _T_1926; // @[Mux.scala 19:72:@2598.4]
  assign _T_2021 = _T_2020 | _T_1928; // @[Mux.scala 19:72:@2599.4]
  assign _T_2022 = _T_2021 | _T_1930; // @[Mux.scala 19:72:@2600.4]
  assign _T_2023 = _T_2022 | _T_1932; // @[Mux.scala 19:72:@2601.4]
  assign _T_2024 = _T_2023 | _T_1934; // @[Mux.scala 19:72:@2602.4]
  assign _T_2025 = _T_2024 | _T_1936; // @[Mux.scala 19:72:@2603.4]
  assign _T_2026 = _T_2025 | _T_1938; // @[Mux.scala 19:72:@2604.4]
  assign _T_2027 = _T_2026 | _T_1940; // @[Mux.scala 19:72:@2605.4]
  assign _T_2028 = _T_2027 | _T_1942; // @[Mux.scala 19:72:@2606.4]
  assign _T_2029 = _T_2028 | _T_1944; // @[Mux.scala 19:72:@2607.4]
  assign _T_2030 = _T_2029 | _T_1946; // @[Mux.scala 19:72:@2608.4]
  assign _T_2031 = _T_2030 | _T_1948; // @[Mux.scala 19:72:@2609.4]
  assign _T_2032 = _T_2031 | _T_1950; // @[Mux.scala 19:72:@2610.4]
  assign _T_2033 = _T_2032 | _T_1952; // @[Mux.scala 19:72:@2611.4]
  assign _T_2034 = _T_2033 | _T_1954; // @[Mux.scala 19:72:@2612.4]
  assign _T_2035 = _T_2034 | _T_1956; // @[Mux.scala 19:72:@2613.4]
  assign _T_2036 = _T_2035 | _T_1958; // @[Mux.scala 19:72:@2614.4]
  assign _T_2037 = _T_2036 | _T_1960; // @[Mux.scala 19:72:@2615.4]
  assign _T_2038 = _T_2037 | _T_1962; // @[Mux.scala 19:72:@2616.4]
  assign _T_2039 = _T_2038 | _T_1964; // @[Mux.scala 19:72:@2617.4]
  assign _T_2040 = _T_2039 | _T_1966; // @[Mux.scala 19:72:@2618.4]
  assign _T_2041 = _T_2040 | _T_1968; // @[Mux.scala 19:72:@2619.4]
  assign _T_2042 = _T_2041 | _T_1970; // @[Mux.scala 19:72:@2620.4]
  assign _T_2043 = _T_2042 | _T_1972; // @[Mux.scala 19:72:@2621.4]
  assign _T_2044 = _T_2043 | _T_1974; // @[Mux.scala 19:72:@2622.4]
  assign _T_2045 = _T_2044 | _T_1976; // @[Mux.scala 19:72:@2623.4]
  assign _T_2046 = _T_2045 | _T_1978; // @[Mux.scala 19:72:@2624.4]
  assign _T_2047 = _T_2046 | _T_1980; // @[Mux.scala 19:72:@2625.4]
  assign _T_2048 = _T_2047 | _T_1982; // @[Mux.scala 19:72:@2626.4]
  assign _T_2049 = _T_2048 | _T_1984; // @[Mux.scala 19:72:@2627.4]
  assign _T_2050 = _T_2049 | _T_1986; // @[Mux.scala 19:72:@2628.4]
  assign predict_1_bj_type = _T_2050 | _T_1988; // @[Mux.scala 19:72:@2629.4]
  assign _T_2120 = _T_1536 ? btb_h_count_0 : 2'h0; // @[Mux.scala 19:72:@2697.4]
  assign _T_2122 = _T_1537 ? btb_h_count_1 : 2'h0; // @[Mux.scala 19:72:@2698.4]
  assign _T_2124 = _T_1538 ? btb_h_count_2 : 2'h0; // @[Mux.scala 19:72:@2699.4]
  assign _T_2126 = _T_1539 ? btb_h_count_3 : 2'h0; // @[Mux.scala 19:72:@2700.4]
  assign _T_2128 = _T_1540 ? btb_h_count_4 : 2'h0; // @[Mux.scala 19:72:@2701.4]
  assign _T_2130 = _T_1541 ? btb_h_count_5 : 2'h0; // @[Mux.scala 19:72:@2702.4]
  assign _T_2132 = _T_1542 ? btb_h_count_6 : 2'h0; // @[Mux.scala 19:72:@2703.4]
  assign _T_2134 = _T_1543 ? btb_h_count_7 : 2'h0; // @[Mux.scala 19:72:@2704.4]
  assign _T_2136 = _T_1544 ? btb_h_count_8 : 2'h0; // @[Mux.scala 19:72:@2705.4]
  assign _T_2138 = _T_1545 ? btb_h_count_9 : 2'h0; // @[Mux.scala 19:72:@2706.4]
  assign _T_2140 = _T_1546 ? btb_h_count_10 : 2'h0; // @[Mux.scala 19:72:@2707.4]
  assign _T_2142 = _T_1547 ? btb_h_count_11 : 2'h0; // @[Mux.scala 19:72:@2708.4]
  assign _T_2144 = _T_1548 ? btb_h_count_12 : 2'h0; // @[Mux.scala 19:72:@2709.4]
  assign _T_2146 = _T_1549 ? btb_h_count_13 : 2'h0; // @[Mux.scala 19:72:@2710.4]
  assign _T_2148 = _T_1550 ? btb_h_count_14 : 2'h0; // @[Mux.scala 19:72:@2711.4]
  assign _T_2150 = _T_1551 ? btb_h_count_15 : 2'h0; // @[Mux.scala 19:72:@2712.4]
  assign _T_2152 = _T_1552 ? btb_h_count_16 : 2'h0; // @[Mux.scala 19:72:@2713.4]
  assign _T_2154 = _T_1553 ? btb_h_count_17 : 2'h0; // @[Mux.scala 19:72:@2714.4]
  assign _T_2156 = _T_1554 ? btb_h_count_18 : 2'h0; // @[Mux.scala 19:72:@2715.4]
  assign _T_2158 = _T_1555 ? btb_h_count_19 : 2'h0; // @[Mux.scala 19:72:@2716.4]
  assign _T_2160 = _T_1556 ? btb_h_count_20 : 2'h0; // @[Mux.scala 19:72:@2717.4]
  assign _T_2162 = _T_1557 ? btb_h_count_21 : 2'h0; // @[Mux.scala 19:72:@2718.4]
  assign _T_2164 = _T_1558 ? btb_h_count_22 : 2'h0; // @[Mux.scala 19:72:@2719.4]
  assign _T_2166 = _T_1559 ? btb_h_count_23 : 2'h0; // @[Mux.scala 19:72:@2720.4]
  assign _T_2168 = _T_1560 ? btb_h_count_24 : 2'h0; // @[Mux.scala 19:72:@2721.4]
  assign _T_2170 = _T_1561 ? btb_h_count_25 : 2'h0; // @[Mux.scala 19:72:@2722.4]
  assign _T_2172 = _T_1562 ? btb_h_count_26 : 2'h0; // @[Mux.scala 19:72:@2723.4]
  assign _T_2174 = _T_1563 ? btb_h_count_27 : 2'h0; // @[Mux.scala 19:72:@2724.4]
  assign _T_2176 = _T_1564 ? btb_h_count_28 : 2'h0; // @[Mux.scala 19:72:@2725.4]
  assign _T_2178 = _T_1565 ? btb_h_count_29 : 2'h0; // @[Mux.scala 19:72:@2726.4]
  assign _T_2180 = _T_1566 ? btb_h_count_30 : 2'h0; // @[Mux.scala 19:72:@2727.4]
  assign _T_2182 = _T_1567 ? btb_h_count_31 : 2'h0; // @[Mux.scala 19:72:@2728.4]
  assign _T_2184 = _T_1568 ? btb_h_count_32 : 2'h0; // @[Mux.scala 19:72:@2729.4]
  assign _T_2186 = _T_1569 ? btb_h_count_33 : 2'h0; // @[Mux.scala 19:72:@2730.4]
  assign _T_2188 = _T_1570 ? btb_h_count_34 : 2'h0; // @[Mux.scala 19:72:@2731.4]
  assign _T_2190 = _T_1571 ? btb_h_count_35 : 2'h0; // @[Mux.scala 19:72:@2732.4]
  assign _T_2192 = _T_1572 ? btb_h_count_36 : 2'h0; // @[Mux.scala 19:72:@2733.4]
  assign _T_2194 = _T_1573 ? btb_h_count_37 : 2'h0; // @[Mux.scala 19:72:@2734.4]
  assign _T_2196 = _T_1574 ? btb_h_count_38 : 2'h0; // @[Mux.scala 19:72:@2735.4]
  assign _T_2198 = _T_1575 ? btb_h_count_39 : 2'h0; // @[Mux.scala 19:72:@2736.4]
  assign _T_2200 = _T_1576 ? btb_h_count_40 : 2'h0; // @[Mux.scala 19:72:@2737.4]
  assign _T_2202 = _T_1577 ? btb_h_count_41 : 2'h0; // @[Mux.scala 19:72:@2738.4]
  assign _T_2204 = _T_1578 ? btb_h_count_42 : 2'h0; // @[Mux.scala 19:72:@2739.4]
  assign _T_2206 = _T_1579 ? btb_h_count_43 : 2'h0; // @[Mux.scala 19:72:@2740.4]
  assign _T_2208 = _T_1580 ? btb_h_count_44 : 2'h0; // @[Mux.scala 19:72:@2741.4]
  assign _T_2210 = _T_1581 ? btb_h_count_45 : 2'h0; // @[Mux.scala 19:72:@2742.4]
  assign _T_2212 = _T_1582 ? btb_h_count_46 : 2'h0; // @[Mux.scala 19:72:@2743.4]
  assign _T_2214 = _T_1583 ? btb_h_count_47 : 2'h0; // @[Mux.scala 19:72:@2744.4]
  assign _T_2216 = _T_1584 ? btb_h_count_48 : 2'h0; // @[Mux.scala 19:72:@2745.4]
  assign _T_2218 = _T_1585 ? btb_h_count_49 : 2'h0; // @[Mux.scala 19:72:@2746.4]
  assign _T_2220 = _T_1586 ? btb_h_count_50 : 2'h0; // @[Mux.scala 19:72:@2747.4]
  assign _T_2222 = _T_1587 ? btb_h_count_51 : 2'h0; // @[Mux.scala 19:72:@2748.4]
  assign _T_2224 = _T_1588 ? btb_h_count_52 : 2'h0; // @[Mux.scala 19:72:@2749.4]
  assign _T_2226 = _T_1589 ? btb_h_count_53 : 2'h0; // @[Mux.scala 19:72:@2750.4]
  assign _T_2228 = _T_1590 ? btb_h_count_54 : 2'h0; // @[Mux.scala 19:72:@2751.4]
  assign _T_2230 = _T_1591 ? btb_h_count_55 : 2'h0; // @[Mux.scala 19:72:@2752.4]
  assign _T_2232 = _T_1592 ? btb_h_count_56 : 2'h0; // @[Mux.scala 19:72:@2753.4]
  assign _T_2234 = _T_1593 ? btb_h_count_57 : 2'h0; // @[Mux.scala 19:72:@2754.4]
  assign _T_2236 = _T_1594 ? btb_h_count_58 : 2'h0; // @[Mux.scala 19:72:@2755.4]
  assign _T_2238 = _T_1595 ? btb_h_count_59 : 2'h0; // @[Mux.scala 19:72:@2756.4]
  assign _T_2240 = _T_1596 ? btb_h_count_60 : 2'h0; // @[Mux.scala 19:72:@2757.4]
  assign _T_2242 = _T_1597 ? btb_h_count_61 : 2'h0; // @[Mux.scala 19:72:@2758.4]
  assign _T_2244 = _T_1598 ? btb_h_count_62 : 2'h0; // @[Mux.scala 19:72:@2759.4]
  assign _T_2246 = _T_1599 ? btb_h_count_63 : 2'h0; // @[Mux.scala 19:72:@2760.4]
  assign _T_2247 = _T_2120 | _T_2122; // @[Mux.scala 19:72:@2761.4]
  assign _T_2248 = _T_2247 | _T_2124; // @[Mux.scala 19:72:@2762.4]
  assign _T_2249 = _T_2248 | _T_2126; // @[Mux.scala 19:72:@2763.4]
  assign _T_2250 = _T_2249 | _T_2128; // @[Mux.scala 19:72:@2764.4]
  assign _T_2251 = _T_2250 | _T_2130; // @[Mux.scala 19:72:@2765.4]
  assign _T_2252 = _T_2251 | _T_2132; // @[Mux.scala 19:72:@2766.4]
  assign _T_2253 = _T_2252 | _T_2134; // @[Mux.scala 19:72:@2767.4]
  assign _T_2254 = _T_2253 | _T_2136; // @[Mux.scala 19:72:@2768.4]
  assign _T_2255 = _T_2254 | _T_2138; // @[Mux.scala 19:72:@2769.4]
  assign _T_2256 = _T_2255 | _T_2140; // @[Mux.scala 19:72:@2770.4]
  assign _T_2257 = _T_2256 | _T_2142; // @[Mux.scala 19:72:@2771.4]
  assign _T_2258 = _T_2257 | _T_2144; // @[Mux.scala 19:72:@2772.4]
  assign _T_2259 = _T_2258 | _T_2146; // @[Mux.scala 19:72:@2773.4]
  assign _T_2260 = _T_2259 | _T_2148; // @[Mux.scala 19:72:@2774.4]
  assign _T_2261 = _T_2260 | _T_2150; // @[Mux.scala 19:72:@2775.4]
  assign _T_2262 = _T_2261 | _T_2152; // @[Mux.scala 19:72:@2776.4]
  assign _T_2263 = _T_2262 | _T_2154; // @[Mux.scala 19:72:@2777.4]
  assign _T_2264 = _T_2263 | _T_2156; // @[Mux.scala 19:72:@2778.4]
  assign _T_2265 = _T_2264 | _T_2158; // @[Mux.scala 19:72:@2779.4]
  assign _T_2266 = _T_2265 | _T_2160; // @[Mux.scala 19:72:@2780.4]
  assign _T_2267 = _T_2266 | _T_2162; // @[Mux.scala 19:72:@2781.4]
  assign _T_2268 = _T_2267 | _T_2164; // @[Mux.scala 19:72:@2782.4]
  assign _T_2269 = _T_2268 | _T_2166; // @[Mux.scala 19:72:@2783.4]
  assign _T_2270 = _T_2269 | _T_2168; // @[Mux.scala 19:72:@2784.4]
  assign _T_2271 = _T_2270 | _T_2170; // @[Mux.scala 19:72:@2785.4]
  assign _T_2272 = _T_2271 | _T_2172; // @[Mux.scala 19:72:@2786.4]
  assign _T_2273 = _T_2272 | _T_2174; // @[Mux.scala 19:72:@2787.4]
  assign _T_2274 = _T_2273 | _T_2176; // @[Mux.scala 19:72:@2788.4]
  assign _T_2275 = _T_2274 | _T_2178; // @[Mux.scala 19:72:@2789.4]
  assign _T_2276 = _T_2275 | _T_2180; // @[Mux.scala 19:72:@2790.4]
  assign _T_2277 = _T_2276 | _T_2182; // @[Mux.scala 19:72:@2791.4]
  assign _T_2278 = _T_2277 | _T_2184; // @[Mux.scala 19:72:@2792.4]
  assign _T_2279 = _T_2278 | _T_2186; // @[Mux.scala 19:72:@2793.4]
  assign _T_2280 = _T_2279 | _T_2188; // @[Mux.scala 19:72:@2794.4]
  assign _T_2281 = _T_2280 | _T_2190; // @[Mux.scala 19:72:@2795.4]
  assign _T_2282 = _T_2281 | _T_2192; // @[Mux.scala 19:72:@2796.4]
  assign _T_2283 = _T_2282 | _T_2194; // @[Mux.scala 19:72:@2797.4]
  assign _T_2284 = _T_2283 | _T_2196; // @[Mux.scala 19:72:@2798.4]
  assign _T_2285 = _T_2284 | _T_2198; // @[Mux.scala 19:72:@2799.4]
  assign _T_2286 = _T_2285 | _T_2200; // @[Mux.scala 19:72:@2800.4]
  assign _T_2287 = _T_2286 | _T_2202; // @[Mux.scala 19:72:@2801.4]
  assign _T_2288 = _T_2287 | _T_2204; // @[Mux.scala 19:72:@2802.4]
  assign _T_2289 = _T_2288 | _T_2206; // @[Mux.scala 19:72:@2803.4]
  assign _T_2290 = _T_2289 | _T_2208; // @[Mux.scala 19:72:@2804.4]
  assign _T_2291 = _T_2290 | _T_2210; // @[Mux.scala 19:72:@2805.4]
  assign _T_2292 = _T_2291 | _T_2212; // @[Mux.scala 19:72:@2806.4]
  assign _T_2293 = _T_2292 | _T_2214; // @[Mux.scala 19:72:@2807.4]
  assign _T_2294 = _T_2293 | _T_2216; // @[Mux.scala 19:72:@2808.4]
  assign _T_2295 = _T_2294 | _T_2218; // @[Mux.scala 19:72:@2809.4]
  assign _T_2296 = _T_2295 | _T_2220; // @[Mux.scala 19:72:@2810.4]
  assign _T_2297 = _T_2296 | _T_2222; // @[Mux.scala 19:72:@2811.4]
  assign _T_2298 = _T_2297 | _T_2224; // @[Mux.scala 19:72:@2812.4]
  assign _T_2299 = _T_2298 | _T_2226; // @[Mux.scala 19:72:@2813.4]
  assign _T_2300 = _T_2299 | _T_2228; // @[Mux.scala 19:72:@2814.4]
  assign _T_2301 = _T_2300 | _T_2230; // @[Mux.scala 19:72:@2815.4]
  assign _T_2302 = _T_2301 | _T_2232; // @[Mux.scala 19:72:@2816.4]
  assign _T_2303 = _T_2302 | _T_2234; // @[Mux.scala 19:72:@2817.4]
  assign _T_2304 = _T_2303 | _T_2236; // @[Mux.scala 19:72:@2818.4]
  assign _T_2305 = _T_2304 | _T_2238; // @[Mux.scala 19:72:@2819.4]
  assign _T_2306 = _T_2305 | _T_2240; // @[Mux.scala 19:72:@2820.4]
  assign _T_2307 = _T_2306 | _T_2242; // @[Mux.scala 19:72:@2821.4]
  assign _T_2308 = _T_2307 | _T_2244; // @[Mux.scala 19:72:@2822.4]
  assign predict_1_h_count = _T_2308 | _T_2246; // @[Mux.scala 19:72:@2823.4]
  assign _T_2313 = _T_178[9:0]; // @[BTB.scala 110:54:@2828.4]
  assign predict_1_gshxor = gb_history ^ _T_2313; // @[BTB.scala 110:44:@2829.4]
  assign predict_1_gshare = bht__T_2316_data; // @[BTB.scala 98:21:@1087.4 BTB.scala 112:25:@2834.4]
  assign _T_2318 = predict_1_gshare[1]; // @[BTB.scala 47:40:@2836.4]
  assign _T_2319 = predict_1_h_count[1]; // @[BTB.scala 47:52:@2837.4]
  assign predict_1_select = arb__T_2315_data; // @[BTB.scala 98:21:@1087.4 BTB.scala 111:25:@2832.4]
  assign _T_2320 = predict_1_select ? _T_2318 : _T_2319; // @[BTB.scala 47:25:@2838.4]
  assign predict_1_history = {_T_1240,_T_2320}; // @[Cat.scala 30:58:@2839.4]
  assign _T_2323 = predict_1_lookup != 64'h0; // @[BTB.scala 40:28:@2841.4]
  assign _T_2327 = predict_1_bj_type != 2'h2; // @[BTB.scala 49:42:@2844.4]
  assign _T_2331 = _T_2327 | _T_2320; // @[BTB.scala 49:63:@2848.4]
  assign _T_2332 = _T_2323 & _T_2331; // @[BTB.scala 49:30:@2849.4]
  assign _T_2337 = predict_1_bj_type == 2'h1; // @[BTB.scala 119:54:@2856.4]
  assign _T_2347 = _T_2332 ? predict_1_jump_tgt : predict_1_cont_tgt; // @[BTB.scala 120:34:@2864.4]
  assign shift_wire = io_branch & shift_reg; // @[BTB.scala 124:30:@2868.4]
  assign _T_2351 = io_fb_type == 2'h2; // @[BTB.scala 126:22:@2870.6]
  assign _T_2352 = io_feedBack_history[8:0]; // @[BTB.scala 127:44:@2872.8]
  assign _T_2353 = {_T_2352,io_feedBack_redirect}; // @[Cat.scala 30:58:@2873.8]
  assign _GEN_0 = _T_2351 ? _T_2353 : io_feedBack_history; // @[BTB.scala 126:44:@2871.6]
  assign _T_2355 = predict_0_bj_type == 2'h2; // @[BTB.scala 46:30:@2882.8]
  assign _T_2360 = _T_2355 & _T_186; // @[BTB.scala 132:38:@2886.8]
  assign _T_2362 = _T_2360 == 1'h0; // @[BTB.scala 132:18:@2887.8]
  assign _T_2364 = predict_1_bj_type == 2'h2; // @[BTB.scala 46:30:@2888.8]
  assign _T_2366 = _T_2364 == 1'h0; // @[BTB.scala 132:79:@2889.8]
  assign _T_2367 = _T_2362 & _T_2366; // @[BTB.scala 132:76:@2890.8]
  assign _T_2370 = {_T_1240,1'h0}; // @[Cat.scala 30:58:@2894.10]
  assign _T_2380 = predict_0_history[8:0]; // @[BTB.scala 137:45:@2906.14]
  assign _T_2384 = {_T_2380,_T_2320}; // @[Cat.scala 30:58:@2910.14]
  assign _GEN_1 = _T_2364 ? _T_2384 : predict_0_history; // @[BTB.scala 136:32:@2905.12]
  assign _GEN_2 = _T_2364 ? predict_1_history : gb_history; // @[BTB.scala 141:35:@2919.12]
  assign _GEN_3 = _T_2360 ? _GEN_1 : _GEN_2; // @[BTB.scala 135:72:@2903.10]
  assign _GEN_4 = shift_wire ? _T_2370 : _GEN_3; // @[BTB.scala 133:23:@2892.8]
  assign _GEN_5 = io_if_pc_valid ? _T_2367 : shift_reg; // @[BTB.scala 131:30:@2881.6]
  assign _GEN_6 = io_if_pc_valid ? _GEN_4 : gb_history; // @[BTB.scala 131:30:@2881.6]
  assign _GEN_7 = io_fb_pc_valid ? _GEN_0 : _GEN_6; // @[BTB.scala 125:25:@2869.4]
  assign _T_2393 = io_fb_pc_bits[31:2]; // @[BTB.scala 176:35:@2936.4]
  assign _T_2394 = io_feedBack_tgt[31:2]; // @[BTB.scala 177:37:@2938.4]
  assign _T_2396 = io_fb_pc_bits[11:2]; // @[BTB.scala 181:62:@2944.4]
  assign _T_2397 = io_feedBack_history ^ _T_2396; // @[BTB.scala 181:47:@2945.4]
  assign _T_2398 = fb_reg_lfsr[0]; // @[BTB.scala 160:22:@2947.4]
  assign _T_2399 = fb_reg_lfsr[1]; // @[BTB.scala 160:32:@2948.4]
  assign _T_2400 = _T_2398 ^ _T_2399; // @[BTB.scala 160:26:@2949.4]
  assign _T_2401 = fb_reg_lfsr[5:1]; // @[BTB.scala 160:41:@2950.4]
  assign _T_2402 = {_T_2400,_T_2401}; // @[Cat.scala 30:58:@2951.4]
  assign _T_2404 = btb_pc_0 == fb_reg_pc; // @[BTB.scala 192:44:@2954.4]
  assign _T_2405 = btb_pc_1 == fb_reg_pc; // @[BTB.scala 192:44:@2955.4]
  assign _T_2406 = btb_pc_2 == fb_reg_pc; // @[BTB.scala 192:44:@2956.4]
  assign _T_2407 = btb_pc_3 == fb_reg_pc; // @[BTB.scala 192:44:@2957.4]
  assign _T_2408 = btb_pc_4 == fb_reg_pc; // @[BTB.scala 192:44:@2958.4]
  assign _T_2409 = btb_pc_5 == fb_reg_pc; // @[BTB.scala 192:44:@2959.4]
  assign _T_2410 = btb_pc_6 == fb_reg_pc; // @[BTB.scala 192:44:@2960.4]
  assign _T_2411 = btb_pc_7 == fb_reg_pc; // @[BTB.scala 192:44:@2961.4]
  assign _T_2412 = btb_pc_8 == fb_reg_pc; // @[BTB.scala 192:44:@2962.4]
  assign _T_2413 = btb_pc_9 == fb_reg_pc; // @[BTB.scala 192:44:@2963.4]
  assign _T_2414 = btb_pc_10 == fb_reg_pc; // @[BTB.scala 192:44:@2964.4]
  assign _T_2415 = btb_pc_11 == fb_reg_pc; // @[BTB.scala 192:44:@2965.4]
  assign _T_2416 = btb_pc_12 == fb_reg_pc; // @[BTB.scala 192:44:@2966.4]
  assign _T_2417 = btb_pc_13 == fb_reg_pc; // @[BTB.scala 192:44:@2967.4]
  assign _T_2418 = btb_pc_14 == fb_reg_pc; // @[BTB.scala 192:44:@2968.4]
  assign _T_2419 = btb_pc_15 == fb_reg_pc; // @[BTB.scala 192:44:@2969.4]
  assign _T_2420 = btb_pc_16 == fb_reg_pc; // @[BTB.scala 192:44:@2970.4]
  assign _T_2421 = btb_pc_17 == fb_reg_pc; // @[BTB.scala 192:44:@2971.4]
  assign _T_2422 = btb_pc_18 == fb_reg_pc; // @[BTB.scala 192:44:@2972.4]
  assign _T_2423 = btb_pc_19 == fb_reg_pc; // @[BTB.scala 192:44:@2973.4]
  assign _T_2424 = btb_pc_20 == fb_reg_pc; // @[BTB.scala 192:44:@2974.4]
  assign _T_2425 = btb_pc_21 == fb_reg_pc; // @[BTB.scala 192:44:@2975.4]
  assign _T_2426 = btb_pc_22 == fb_reg_pc; // @[BTB.scala 192:44:@2976.4]
  assign _T_2427 = btb_pc_23 == fb_reg_pc; // @[BTB.scala 192:44:@2977.4]
  assign _T_2428 = btb_pc_24 == fb_reg_pc; // @[BTB.scala 192:44:@2978.4]
  assign _T_2429 = btb_pc_25 == fb_reg_pc; // @[BTB.scala 192:44:@2979.4]
  assign _T_2430 = btb_pc_26 == fb_reg_pc; // @[BTB.scala 192:44:@2980.4]
  assign _T_2431 = btb_pc_27 == fb_reg_pc; // @[BTB.scala 192:44:@2981.4]
  assign _T_2432 = btb_pc_28 == fb_reg_pc; // @[BTB.scala 192:44:@2982.4]
  assign _T_2433 = btb_pc_29 == fb_reg_pc; // @[BTB.scala 192:44:@2983.4]
  assign _T_2434 = btb_pc_30 == fb_reg_pc; // @[BTB.scala 192:44:@2984.4]
  assign _T_2435 = btb_pc_31 == fb_reg_pc; // @[BTB.scala 192:44:@2985.4]
  assign _T_2436 = btb_pc_32 == fb_reg_pc; // @[BTB.scala 192:44:@2986.4]
  assign _T_2437 = btb_pc_33 == fb_reg_pc; // @[BTB.scala 192:44:@2987.4]
  assign _T_2438 = btb_pc_34 == fb_reg_pc; // @[BTB.scala 192:44:@2988.4]
  assign _T_2439 = btb_pc_35 == fb_reg_pc; // @[BTB.scala 192:44:@2989.4]
  assign _T_2440 = btb_pc_36 == fb_reg_pc; // @[BTB.scala 192:44:@2990.4]
  assign _T_2441 = btb_pc_37 == fb_reg_pc; // @[BTB.scala 192:44:@2991.4]
  assign _T_2442 = btb_pc_38 == fb_reg_pc; // @[BTB.scala 192:44:@2992.4]
  assign _T_2443 = btb_pc_39 == fb_reg_pc; // @[BTB.scala 192:44:@2993.4]
  assign _T_2444 = btb_pc_40 == fb_reg_pc; // @[BTB.scala 192:44:@2994.4]
  assign _T_2445 = btb_pc_41 == fb_reg_pc; // @[BTB.scala 192:44:@2995.4]
  assign _T_2446 = btb_pc_42 == fb_reg_pc; // @[BTB.scala 192:44:@2996.4]
  assign _T_2447 = btb_pc_43 == fb_reg_pc; // @[BTB.scala 192:44:@2997.4]
  assign _T_2448 = btb_pc_44 == fb_reg_pc; // @[BTB.scala 192:44:@2998.4]
  assign _T_2449 = btb_pc_45 == fb_reg_pc; // @[BTB.scala 192:44:@2999.4]
  assign _T_2450 = btb_pc_46 == fb_reg_pc; // @[BTB.scala 192:44:@3000.4]
  assign _T_2451 = btb_pc_47 == fb_reg_pc; // @[BTB.scala 192:44:@3001.4]
  assign _T_2452 = btb_pc_48 == fb_reg_pc; // @[BTB.scala 192:44:@3002.4]
  assign _T_2453 = btb_pc_49 == fb_reg_pc; // @[BTB.scala 192:44:@3003.4]
  assign _T_2454 = btb_pc_50 == fb_reg_pc; // @[BTB.scala 192:44:@3004.4]
  assign _T_2455 = btb_pc_51 == fb_reg_pc; // @[BTB.scala 192:44:@3005.4]
  assign _T_2456 = btb_pc_52 == fb_reg_pc; // @[BTB.scala 192:44:@3006.4]
  assign _T_2457 = btb_pc_53 == fb_reg_pc; // @[BTB.scala 192:44:@3007.4]
  assign _T_2458 = btb_pc_54 == fb_reg_pc; // @[BTB.scala 192:44:@3008.4]
  assign _T_2459 = btb_pc_55 == fb_reg_pc; // @[BTB.scala 192:44:@3009.4]
  assign _T_2460 = btb_pc_56 == fb_reg_pc; // @[BTB.scala 192:44:@3010.4]
  assign _T_2461 = btb_pc_57 == fb_reg_pc; // @[BTB.scala 192:44:@3011.4]
  assign _T_2462 = btb_pc_58 == fb_reg_pc; // @[BTB.scala 192:44:@3012.4]
  assign _T_2463 = btb_pc_59 == fb_reg_pc; // @[BTB.scala 192:44:@3013.4]
  assign _T_2464 = btb_pc_60 == fb_reg_pc; // @[BTB.scala 192:44:@3014.4]
  assign _T_2465 = btb_pc_61 == fb_reg_pc; // @[BTB.scala 192:44:@3015.4]
  assign _T_2466 = btb_pc_62 == fb_reg_pc; // @[BTB.scala 192:44:@3016.4]
  assign _T_2467 = btb_pc_63 == fb_reg_pc; // @[BTB.scala 192:44:@3017.4]
  assign _T_2544 = {_T_2411,_T_2410,_T_2409,_T_2408,_T_2407,_T_2406,_T_2405,_T_2404}; // @[BTB.scala 192:60:@3089.4]
  assign _T_2552 = {_T_2419,_T_2418,_T_2417,_T_2416,_T_2415,_T_2414,_T_2413,_T_2412,_T_2544}; // @[BTB.scala 192:60:@3097.4]
  assign _T_2559 = {_T_2427,_T_2426,_T_2425,_T_2424,_T_2423,_T_2422,_T_2421,_T_2420}; // @[BTB.scala 192:60:@3104.4]
  assign _T_2568 = {_T_2435,_T_2434,_T_2433,_T_2432,_T_2431,_T_2430,_T_2429,_T_2428,_T_2559,_T_2552}; // @[BTB.scala 192:60:@3113.4]
  assign _T_2575 = {_T_2443,_T_2442,_T_2441,_T_2440,_T_2439,_T_2438,_T_2437,_T_2436}; // @[BTB.scala 192:60:@3120.4]
  assign _T_2583 = {_T_2451,_T_2450,_T_2449,_T_2448,_T_2447,_T_2446,_T_2445,_T_2444,_T_2575}; // @[BTB.scala 192:60:@3128.4]
  assign _T_2590 = {_T_2459,_T_2458,_T_2457,_T_2456,_T_2455,_T_2454,_T_2453,_T_2452}; // @[BTB.scala 192:60:@3135.4]
  assign _T_2599 = {_T_2467,_T_2466,_T_2465,_T_2464,_T_2463,_T_2462,_T_2461,_T_2460,_T_2590,_T_2583}; // @[BTB.scala 192:60:@3144.4]
  assign _T_2600 = {_T_2599,_T_2568}; // @[BTB.scala 192:60:@3145.4]
  assign feedback_lookup = _T_2600 & _T_457; // @[BTB.scala 192:67:@3209.4]
  assign _T_2665 = feedback_lookup[0]; // @[Mux.scala 21:36:@3211.4]
  assign _T_2666 = feedback_lookup[1]; // @[Mux.scala 21:36:@3212.4]
  assign _T_2667 = feedback_lookup[2]; // @[Mux.scala 21:36:@3213.4]
  assign _T_2668 = feedback_lookup[3]; // @[Mux.scala 21:36:@3214.4]
  assign _T_2669 = feedback_lookup[4]; // @[Mux.scala 21:36:@3215.4]
  assign _T_2670 = feedback_lookup[5]; // @[Mux.scala 21:36:@3216.4]
  assign _T_2671 = feedback_lookup[6]; // @[Mux.scala 21:36:@3217.4]
  assign _T_2672 = feedback_lookup[7]; // @[Mux.scala 21:36:@3218.4]
  assign _T_2673 = feedback_lookup[8]; // @[Mux.scala 21:36:@3219.4]
  assign _T_2674 = feedback_lookup[9]; // @[Mux.scala 21:36:@3220.4]
  assign _T_2675 = feedback_lookup[10]; // @[Mux.scala 21:36:@3221.4]
  assign _T_2676 = feedback_lookup[11]; // @[Mux.scala 21:36:@3222.4]
  assign _T_2677 = feedback_lookup[12]; // @[Mux.scala 21:36:@3223.4]
  assign _T_2678 = feedback_lookup[13]; // @[Mux.scala 21:36:@3224.4]
  assign _T_2679 = feedback_lookup[14]; // @[Mux.scala 21:36:@3225.4]
  assign _T_2680 = feedback_lookup[15]; // @[Mux.scala 21:36:@3226.4]
  assign _T_2681 = feedback_lookup[16]; // @[Mux.scala 21:36:@3227.4]
  assign _T_2682 = feedback_lookup[17]; // @[Mux.scala 21:36:@3228.4]
  assign _T_2683 = feedback_lookup[18]; // @[Mux.scala 21:36:@3229.4]
  assign _T_2684 = feedback_lookup[19]; // @[Mux.scala 21:36:@3230.4]
  assign _T_2685 = feedback_lookup[20]; // @[Mux.scala 21:36:@3231.4]
  assign _T_2686 = feedback_lookup[21]; // @[Mux.scala 21:36:@3232.4]
  assign _T_2687 = feedback_lookup[22]; // @[Mux.scala 21:36:@3233.4]
  assign _T_2688 = feedback_lookup[23]; // @[Mux.scala 21:36:@3234.4]
  assign _T_2689 = feedback_lookup[24]; // @[Mux.scala 21:36:@3235.4]
  assign _T_2690 = feedback_lookup[25]; // @[Mux.scala 21:36:@3236.4]
  assign _T_2691 = feedback_lookup[26]; // @[Mux.scala 21:36:@3237.4]
  assign _T_2692 = feedback_lookup[27]; // @[Mux.scala 21:36:@3238.4]
  assign _T_2693 = feedback_lookup[28]; // @[Mux.scala 21:36:@3239.4]
  assign _T_2694 = feedback_lookup[29]; // @[Mux.scala 21:36:@3240.4]
  assign _T_2695 = feedback_lookup[30]; // @[Mux.scala 21:36:@3241.4]
  assign _T_2696 = feedback_lookup[31]; // @[Mux.scala 21:36:@3242.4]
  assign _T_2697 = feedback_lookup[32]; // @[Mux.scala 21:36:@3243.4]
  assign _T_2698 = feedback_lookup[33]; // @[Mux.scala 21:36:@3244.4]
  assign _T_2699 = feedback_lookup[34]; // @[Mux.scala 21:36:@3245.4]
  assign _T_2700 = feedback_lookup[35]; // @[Mux.scala 21:36:@3246.4]
  assign _T_2701 = feedback_lookup[36]; // @[Mux.scala 21:36:@3247.4]
  assign _T_2702 = feedback_lookup[37]; // @[Mux.scala 21:36:@3248.4]
  assign _T_2703 = feedback_lookup[38]; // @[Mux.scala 21:36:@3249.4]
  assign _T_2704 = feedback_lookup[39]; // @[Mux.scala 21:36:@3250.4]
  assign _T_2705 = feedback_lookup[40]; // @[Mux.scala 21:36:@3251.4]
  assign _T_2706 = feedback_lookup[41]; // @[Mux.scala 21:36:@3252.4]
  assign _T_2707 = feedback_lookup[42]; // @[Mux.scala 21:36:@3253.4]
  assign _T_2708 = feedback_lookup[43]; // @[Mux.scala 21:36:@3254.4]
  assign _T_2709 = feedback_lookup[44]; // @[Mux.scala 21:36:@3255.4]
  assign _T_2710 = feedback_lookup[45]; // @[Mux.scala 21:36:@3256.4]
  assign _T_2711 = feedback_lookup[46]; // @[Mux.scala 21:36:@3257.4]
  assign _T_2712 = feedback_lookup[47]; // @[Mux.scala 21:36:@3258.4]
  assign _T_2713 = feedback_lookup[48]; // @[Mux.scala 21:36:@3259.4]
  assign _T_2714 = feedback_lookup[49]; // @[Mux.scala 21:36:@3260.4]
  assign _T_2715 = feedback_lookup[50]; // @[Mux.scala 21:36:@3261.4]
  assign _T_2716 = feedback_lookup[51]; // @[Mux.scala 21:36:@3262.4]
  assign _T_2717 = feedback_lookup[52]; // @[Mux.scala 21:36:@3263.4]
  assign _T_2718 = feedback_lookup[53]; // @[Mux.scala 21:36:@3264.4]
  assign _T_2719 = feedback_lookup[54]; // @[Mux.scala 21:36:@3265.4]
  assign _T_2720 = feedback_lookup[55]; // @[Mux.scala 21:36:@3266.4]
  assign _T_2721 = feedback_lookup[56]; // @[Mux.scala 21:36:@3267.4]
  assign _T_2722 = feedback_lookup[57]; // @[Mux.scala 21:36:@3268.4]
  assign _T_2723 = feedback_lookup[58]; // @[Mux.scala 21:36:@3269.4]
  assign _T_2724 = feedback_lookup[59]; // @[Mux.scala 21:36:@3270.4]
  assign _T_2725 = feedback_lookup[60]; // @[Mux.scala 21:36:@3271.4]
  assign _T_2726 = feedback_lookup[61]; // @[Mux.scala 21:36:@3272.4]
  assign _T_2727 = feedback_lookup[62]; // @[Mux.scala 21:36:@3273.4]
  assign _T_2728 = feedback_lookup[63]; // @[Mux.scala 21:36:@3274.4]
  assign _T_2731 = _T_2665 ? btb_h_count_0 : 2'h0; // @[Mux.scala 19:72:@3275.4]
  assign _T_2733 = _T_2666 ? btb_h_count_1 : 2'h0; // @[Mux.scala 19:72:@3276.4]
  assign _T_2735 = _T_2667 ? btb_h_count_2 : 2'h0; // @[Mux.scala 19:72:@3277.4]
  assign _T_2737 = _T_2668 ? btb_h_count_3 : 2'h0; // @[Mux.scala 19:72:@3278.4]
  assign _T_2739 = _T_2669 ? btb_h_count_4 : 2'h0; // @[Mux.scala 19:72:@3279.4]
  assign _T_2741 = _T_2670 ? btb_h_count_5 : 2'h0; // @[Mux.scala 19:72:@3280.4]
  assign _T_2743 = _T_2671 ? btb_h_count_6 : 2'h0; // @[Mux.scala 19:72:@3281.4]
  assign _T_2745 = _T_2672 ? btb_h_count_7 : 2'h0; // @[Mux.scala 19:72:@3282.4]
  assign _T_2747 = _T_2673 ? btb_h_count_8 : 2'h0; // @[Mux.scala 19:72:@3283.4]
  assign _T_2749 = _T_2674 ? btb_h_count_9 : 2'h0; // @[Mux.scala 19:72:@3284.4]
  assign _T_2751 = _T_2675 ? btb_h_count_10 : 2'h0; // @[Mux.scala 19:72:@3285.4]
  assign _T_2753 = _T_2676 ? btb_h_count_11 : 2'h0; // @[Mux.scala 19:72:@3286.4]
  assign _T_2755 = _T_2677 ? btb_h_count_12 : 2'h0; // @[Mux.scala 19:72:@3287.4]
  assign _T_2757 = _T_2678 ? btb_h_count_13 : 2'h0; // @[Mux.scala 19:72:@3288.4]
  assign _T_2759 = _T_2679 ? btb_h_count_14 : 2'h0; // @[Mux.scala 19:72:@3289.4]
  assign _T_2761 = _T_2680 ? btb_h_count_15 : 2'h0; // @[Mux.scala 19:72:@3290.4]
  assign _T_2763 = _T_2681 ? btb_h_count_16 : 2'h0; // @[Mux.scala 19:72:@3291.4]
  assign _T_2765 = _T_2682 ? btb_h_count_17 : 2'h0; // @[Mux.scala 19:72:@3292.4]
  assign _T_2767 = _T_2683 ? btb_h_count_18 : 2'h0; // @[Mux.scala 19:72:@3293.4]
  assign _T_2769 = _T_2684 ? btb_h_count_19 : 2'h0; // @[Mux.scala 19:72:@3294.4]
  assign _T_2771 = _T_2685 ? btb_h_count_20 : 2'h0; // @[Mux.scala 19:72:@3295.4]
  assign _T_2773 = _T_2686 ? btb_h_count_21 : 2'h0; // @[Mux.scala 19:72:@3296.4]
  assign _T_2775 = _T_2687 ? btb_h_count_22 : 2'h0; // @[Mux.scala 19:72:@3297.4]
  assign _T_2777 = _T_2688 ? btb_h_count_23 : 2'h0; // @[Mux.scala 19:72:@3298.4]
  assign _T_2779 = _T_2689 ? btb_h_count_24 : 2'h0; // @[Mux.scala 19:72:@3299.4]
  assign _T_2781 = _T_2690 ? btb_h_count_25 : 2'h0; // @[Mux.scala 19:72:@3300.4]
  assign _T_2783 = _T_2691 ? btb_h_count_26 : 2'h0; // @[Mux.scala 19:72:@3301.4]
  assign _T_2785 = _T_2692 ? btb_h_count_27 : 2'h0; // @[Mux.scala 19:72:@3302.4]
  assign _T_2787 = _T_2693 ? btb_h_count_28 : 2'h0; // @[Mux.scala 19:72:@3303.4]
  assign _T_2789 = _T_2694 ? btb_h_count_29 : 2'h0; // @[Mux.scala 19:72:@3304.4]
  assign _T_2791 = _T_2695 ? btb_h_count_30 : 2'h0; // @[Mux.scala 19:72:@3305.4]
  assign _T_2793 = _T_2696 ? btb_h_count_31 : 2'h0; // @[Mux.scala 19:72:@3306.4]
  assign _T_2795 = _T_2697 ? btb_h_count_32 : 2'h0; // @[Mux.scala 19:72:@3307.4]
  assign _T_2797 = _T_2698 ? btb_h_count_33 : 2'h0; // @[Mux.scala 19:72:@3308.4]
  assign _T_2799 = _T_2699 ? btb_h_count_34 : 2'h0; // @[Mux.scala 19:72:@3309.4]
  assign _T_2801 = _T_2700 ? btb_h_count_35 : 2'h0; // @[Mux.scala 19:72:@3310.4]
  assign _T_2803 = _T_2701 ? btb_h_count_36 : 2'h0; // @[Mux.scala 19:72:@3311.4]
  assign _T_2805 = _T_2702 ? btb_h_count_37 : 2'h0; // @[Mux.scala 19:72:@3312.4]
  assign _T_2807 = _T_2703 ? btb_h_count_38 : 2'h0; // @[Mux.scala 19:72:@3313.4]
  assign _T_2809 = _T_2704 ? btb_h_count_39 : 2'h0; // @[Mux.scala 19:72:@3314.4]
  assign _T_2811 = _T_2705 ? btb_h_count_40 : 2'h0; // @[Mux.scala 19:72:@3315.4]
  assign _T_2813 = _T_2706 ? btb_h_count_41 : 2'h0; // @[Mux.scala 19:72:@3316.4]
  assign _T_2815 = _T_2707 ? btb_h_count_42 : 2'h0; // @[Mux.scala 19:72:@3317.4]
  assign _T_2817 = _T_2708 ? btb_h_count_43 : 2'h0; // @[Mux.scala 19:72:@3318.4]
  assign _T_2819 = _T_2709 ? btb_h_count_44 : 2'h0; // @[Mux.scala 19:72:@3319.4]
  assign _T_2821 = _T_2710 ? btb_h_count_45 : 2'h0; // @[Mux.scala 19:72:@3320.4]
  assign _T_2823 = _T_2711 ? btb_h_count_46 : 2'h0; // @[Mux.scala 19:72:@3321.4]
  assign _T_2825 = _T_2712 ? btb_h_count_47 : 2'h0; // @[Mux.scala 19:72:@3322.4]
  assign _T_2827 = _T_2713 ? btb_h_count_48 : 2'h0; // @[Mux.scala 19:72:@3323.4]
  assign _T_2829 = _T_2714 ? btb_h_count_49 : 2'h0; // @[Mux.scala 19:72:@3324.4]
  assign _T_2831 = _T_2715 ? btb_h_count_50 : 2'h0; // @[Mux.scala 19:72:@3325.4]
  assign _T_2833 = _T_2716 ? btb_h_count_51 : 2'h0; // @[Mux.scala 19:72:@3326.4]
  assign _T_2835 = _T_2717 ? btb_h_count_52 : 2'h0; // @[Mux.scala 19:72:@3327.4]
  assign _T_2837 = _T_2718 ? btb_h_count_53 : 2'h0; // @[Mux.scala 19:72:@3328.4]
  assign _T_2839 = _T_2719 ? btb_h_count_54 : 2'h0; // @[Mux.scala 19:72:@3329.4]
  assign _T_2841 = _T_2720 ? btb_h_count_55 : 2'h0; // @[Mux.scala 19:72:@3330.4]
  assign _T_2843 = _T_2721 ? btb_h_count_56 : 2'h0; // @[Mux.scala 19:72:@3331.4]
  assign _T_2845 = _T_2722 ? btb_h_count_57 : 2'h0; // @[Mux.scala 19:72:@3332.4]
  assign _T_2847 = _T_2723 ? btb_h_count_58 : 2'h0; // @[Mux.scala 19:72:@3333.4]
  assign _T_2849 = _T_2724 ? btb_h_count_59 : 2'h0; // @[Mux.scala 19:72:@3334.4]
  assign _T_2851 = _T_2725 ? btb_h_count_60 : 2'h0; // @[Mux.scala 19:72:@3335.4]
  assign _T_2853 = _T_2726 ? btb_h_count_61 : 2'h0; // @[Mux.scala 19:72:@3336.4]
  assign _T_2855 = _T_2727 ? btb_h_count_62 : 2'h0; // @[Mux.scala 19:72:@3337.4]
  assign _T_2857 = _T_2728 ? btb_h_count_63 : 2'h0; // @[Mux.scala 19:72:@3338.4]
  assign _T_2858 = _T_2731 | _T_2733; // @[Mux.scala 19:72:@3339.4]
  assign _T_2859 = _T_2858 | _T_2735; // @[Mux.scala 19:72:@3340.4]
  assign _T_2860 = _T_2859 | _T_2737; // @[Mux.scala 19:72:@3341.4]
  assign _T_2861 = _T_2860 | _T_2739; // @[Mux.scala 19:72:@3342.4]
  assign _T_2862 = _T_2861 | _T_2741; // @[Mux.scala 19:72:@3343.4]
  assign _T_2863 = _T_2862 | _T_2743; // @[Mux.scala 19:72:@3344.4]
  assign _T_2864 = _T_2863 | _T_2745; // @[Mux.scala 19:72:@3345.4]
  assign _T_2865 = _T_2864 | _T_2747; // @[Mux.scala 19:72:@3346.4]
  assign _T_2866 = _T_2865 | _T_2749; // @[Mux.scala 19:72:@3347.4]
  assign _T_2867 = _T_2866 | _T_2751; // @[Mux.scala 19:72:@3348.4]
  assign _T_2868 = _T_2867 | _T_2753; // @[Mux.scala 19:72:@3349.4]
  assign _T_2869 = _T_2868 | _T_2755; // @[Mux.scala 19:72:@3350.4]
  assign _T_2870 = _T_2869 | _T_2757; // @[Mux.scala 19:72:@3351.4]
  assign _T_2871 = _T_2870 | _T_2759; // @[Mux.scala 19:72:@3352.4]
  assign _T_2872 = _T_2871 | _T_2761; // @[Mux.scala 19:72:@3353.4]
  assign _T_2873 = _T_2872 | _T_2763; // @[Mux.scala 19:72:@3354.4]
  assign _T_2874 = _T_2873 | _T_2765; // @[Mux.scala 19:72:@3355.4]
  assign _T_2875 = _T_2874 | _T_2767; // @[Mux.scala 19:72:@3356.4]
  assign _T_2876 = _T_2875 | _T_2769; // @[Mux.scala 19:72:@3357.4]
  assign _T_2877 = _T_2876 | _T_2771; // @[Mux.scala 19:72:@3358.4]
  assign _T_2878 = _T_2877 | _T_2773; // @[Mux.scala 19:72:@3359.4]
  assign _T_2879 = _T_2878 | _T_2775; // @[Mux.scala 19:72:@3360.4]
  assign _T_2880 = _T_2879 | _T_2777; // @[Mux.scala 19:72:@3361.4]
  assign _T_2881 = _T_2880 | _T_2779; // @[Mux.scala 19:72:@3362.4]
  assign _T_2882 = _T_2881 | _T_2781; // @[Mux.scala 19:72:@3363.4]
  assign _T_2883 = _T_2882 | _T_2783; // @[Mux.scala 19:72:@3364.4]
  assign _T_2884 = _T_2883 | _T_2785; // @[Mux.scala 19:72:@3365.4]
  assign _T_2885 = _T_2884 | _T_2787; // @[Mux.scala 19:72:@3366.4]
  assign _T_2886 = _T_2885 | _T_2789; // @[Mux.scala 19:72:@3367.4]
  assign _T_2887 = _T_2886 | _T_2791; // @[Mux.scala 19:72:@3368.4]
  assign _T_2888 = _T_2887 | _T_2793; // @[Mux.scala 19:72:@3369.4]
  assign _T_2889 = _T_2888 | _T_2795; // @[Mux.scala 19:72:@3370.4]
  assign _T_2890 = _T_2889 | _T_2797; // @[Mux.scala 19:72:@3371.4]
  assign _T_2891 = _T_2890 | _T_2799; // @[Mux.scala 19:72:@3372.4]
  assign _T_2892 = _T_2891 | _T_2801; // @[Mux.scala 19:72:@3373.4]
  assign _T_2893 = _T_2892 | _T_2803; // @[Mux.scala 19:72:@3374.4]
  assign _T_2894 = _T_2893 | _T_2805; // @[Mux.scala 19:72:@3375.4]
  assign _T_2895 = _T_2894 | _T_2807; // @[Mux.scala 19:72:@3376.4]
  assign _T_2896 = _T_2895 | _T_2809; // @[Mux.scala 19:72:@3377.4]
  assign _T_2897 = _T_2896 | _T_2811; // @[Mux.scala 19:72:@3378.4]
  assign _T_2898 = _T_2897 | _T_2813; // @[Mux.scala 19:72:@3379.4]
  assign _T_2899 = _T_2898 | _T_2815; // @[Mux.scala 19:72:@3380.4]
  assign _T_2900 = _T_2899 | _T_2817; // @[Mux.scala 19:72:@3381.4]
  assign _T_2901 = _T_2900 | _T_2819; // @[Mux.scala 19:72:@3382.4]
  assign _T_2902 = _T_2901 | _T_2821; // @[Mux.scala 19:72:@3383.4]
  assign _T_2903 = _T_2902 | _T_2823; // @[Mux.scala 19:72:@3384.4]
  assign _T_2904 = _T_2903 | _T_2825; // @[Mux.scala 19:72:@3385.4]
  assign _T_2905 = _T_2904 | _T_2827; // @[Mux.scala 19:72:@3386.4]
  assign _T_2906 = _T_2905 | _T_2829; // @[Mux.scala 19:72:@3387.4]
  assign _T_2907 = _T_2906 | _T_2831; // @[Mux.scala 19:72:@3388.4]
  assign _T_2908 = _T_2907 | _T_2833; // @[Mux.scala 19:72:@3389.4]
  assign _T_2909 = _T_2908 | _T_2835; // @[Mux.scala 19:72:@3390.4]
  assign _T_2910 = _T_2909 | _T_2837; // @[Mux.scala 19:72:@3391.4]
  assign _T_2911 = _T_2910 | _T_2839; // @[Mux.scala 19:72:@3392.4]
  assign _T_2912 = _T_2911 | _T_2841; // @[Mux.scala 19:72:@3393.4]
  assign _T_2913 = _T_2912 | _T_2843; // @[Mux.scala 19:72:@3394.4]
  assign _T_2914 = _T_2913 | _T_2845; // @[Mux.scala 19:72:@3395.4]
  assign _T_2915 = _T_2914 | _T_2847; // @[Mux.scala 19:72:@3396.4]
  assign _T_2916 = _T_2915 | _T_2849; // @[Mux.scala 19:72:@3397.4]
  assign _T_2917 = _T_2916 | _T_2851; // @[Mux.scala 19:72:@3398.4]
  assign _T_2918 = _T_2917 | _T_2853; // @[Mux.scala 19:72:@3399.4]
  assign _T_2919 = _T_2918 | _T_2855; // @[Mux.scala 19:72:@3400.4]
  assign feedback_h_count = _T_2919 | _T_2857; // @[Mux.scala 19:72:@3401.4]
  assign _T_2925 = feedback_lookup != 64'h0; // @[BTB.scala 186:30:@3407.4]
  assign _T_2926 = feedback_lookup[63:32]; // @[OneHot.scala 26:18:@3408.4]
  assign _T_2927 = feedback_lookup[31:0]; // @[OneHot.scala 27:18:@3409.4]
  assign _T_2929 = _T_2926 != 32'h0; // @[OneHot.scala 28:14:@3410.4]
  assign _T_2930 = _T_2926 | _T_2927; // @[OneHot.scala 28:28:@3411.4]
  assign _T_2931 = _T_2930[31:16]; // @[OneHot.scala 26:18:@3412.4]
  assign _T_2932 = _T_2930[15:0]; // @[OneHot.scala 27:18:@3413.4]
  assign _T_2934 = _T_2931 != 16'h0; // @[OneHot.scala 28:14:@3414.4]
  assign _T_2935 = _T_2931 | _T_2932; // @[OneHot.scala 28:28:@3415.4]
  assign _T_2936 = _T_2935[15:8]; // @[OneHot.scala 26:18:@3416.4]
  assign _T_2937 = _T_2935[7:0]; // @[OneHot.scala 27:18:@3417.4]
  assign _T_2939 = _T_2936 != 8'h0; // @[OneHot.scala 28:14:@3418.4]
  assign _T_2940 = _T_2936 | _T_2937; // @[OneHot.scala 28:28:@3419.4]
  assign _T_2941 = _T_2940[7:4]; // @[OneHot.scala 26:18:@3420.4]
  assign _T_2942 = _T_2940[3:0]; // @[OneHot.scala 27:18:@3421.4]
  assign _T_2944 = _T_2941 != 4'h0; // @[OneHot.scala 28:14:@3422.4]
  assign _T_2945 = _T_2941 | _T_2942; // @[OneHot.scala 28:28:@3423.4]
  assign _T_2946 = _T_2945[3:2]; // @[OneHot.scala 26:18:@3424.4]
  assign _T_2947 = _T_2945[1:0]; // @[OneHot.scala 27:18:@3425.4]
  assign _T_2949 = _T_2946 != 2'h0; // @[OneHot.scala 28:14:@3426.4]
  assign _T_2950 = _T_2946 | _T_2947; // @[OneHot.scala 28:28:@3427.4]
  assign _T_2951 = _T_2950[1]; // @[CircuitMath.scala 30:8:@3428.4]
  assign _T_2956 = {_T_2929,_T_2934,_T_2939,_T_2944,_T_2949,_T_2951}; // @[Cat.scala 30:58:@3433.4]
  assign _T_3020 = ~ _T_457; // @[BTB.scala 196:26:@3497.4]
  assign _T_3022 = _T_3020 == 64'h0; // @[BTB.scala 196:26:@3498.4]
  assign _T_3087 = _T_3020[0]; // @[OneHot.scala 39:40:@3563.4]
  assign _T_3088 = _T_3020[1]; // @[OneHot.scala 39:40:@3564.4]
  assign _T_3089 = _T_3020[2]; // @[OneHot.scala 39:40:@3565.4]
  assign _T_3090 = _T_3020[3]; // @[OneHot.scala 39:40:@3566.4]
  assign _T_3091 = _T_3020[4]; // @[OneHot.scala 39:40:@3567.4]
  assign _T_3092 = _T_3020[5]; // @[OneHot.scala 39:40:@3568.4]
  assign _T_3093 = _T_3020[6]; // @[OneHot.scala 39:40:@3569.4]
  assign _T_3094 = _T_3020[7]; // @[OneHot.scala 39:40:@3570.4]
  assign _T_3095 = _T_3020[8]; // @[OneHot.scala 39:40:@3571.4]
  assign _T_3096 = _T_3020[9]; // @[OneHot.scala 39:40:@3572.4]
  assign _T_3097 = _T_3020[10]; // @[OneHot.scala 39:40:@3573.4]
  assign _T_3098 = _T_3020[11]; // @[OneHot.scala 39:40:@3574.4]
  assign _T_3099 = _T_3020[12]; // @[OneHot.scala 39:40:@3575.4]
  assign _T_3100 = _T_3020[13]; // @[OneHot.scala 39:40:@3576.4]
  assign _T_3101 = _T_3020[14]; // @[OneHot.scala 39:40:@3577.4]
  assign _T_3102 = _T_3020[15]; // @[OneHot.scala 39:40:@3578.4]
  assign _T_3103 = _T_3020[16]; // @[OneHot.scala 39:40:@3579.4]
  assign _T_3104 = _T_3020[17]; // @[OneHot.scala 39:40:@3580.4]
  assign _T_3105 = _T_3020[18]; // @[OneHot.scala 39:40:@3581.4]
  assign _T_3106 = _T_3020[19]; // @[OneHot.scala 39:40:@3582.4]
  assign _T_3107 = _T_3020[20]; // @[OneHot.scala 39:40:@3583.4]
  assign _T_3108 = _T_3020[21]; // @[OneHot.scala 39:40:@3584.4]
  assign _T_3109 = _T_3020[22]; // @[OneHot.scala 39:40:@3585.4]
  assign _T_3110 = _T_3020[23]; // @[OneHot.scala 39:40:@3586.4]
  assign _T_3111 = _T_3020[24]; // @[OneHot.scala 39:40:@3587.4]
  assign _T_3112 = _T_3020[25]; // @[OneHot.scala 39:40:@3588.4]
  assign _T_3113 = _T_3020[26]; // @[OneHot.scala 39:40:@3589.4]
  assign _T_3114 = _T_3020[27]; // @[OneHot.scala 39:40:@3590.4]
  assign _T_3115 = _T_3020[28]; // @[OneHot.scala 39:40:@3591.4]
  assign _T_3116 = _T_3020[29]; // @[OneHot.scala 39:40:@3592.4]
  assign _T_3117 = _T_3020[30]; // @[OneHot.scala 39:40:@3593.4]
  assign _T_3118 = _T_3020[31]; // @[OneHot.scala 39:40:@3594.4]
  assign _T_3119 = _T_3020[32]; // @[OneHot.scala 39:40:@3595.4]
  assign _T_3120 = _T_3020[33]; // @[OneHot.scala 39:40:@3596.4]
  assign _T_3121 = _T_3020[34]; // @[OneHot.scala 39:40:@3597.4]
  assign _T_3122 = _T_3020[35]; // @[OneHot.scala 39:40:@3598.4]
  assign _T_3123 = _T_3020[36]; // @[OneHot.scala 39:40:@3599.4]
  assign _T_3124 = _T_3020[37]; // @[OneHot.scala 39:40:@3600.4]
  assign _T_3125 = _T_3020[38]; // @[OneHot.scala 39:40:@3601.4]
  assign _T_3126 = _T_3020[39]; // @[OneHot.scala 39:40:@3602.4]
  assign _T_3127 = _T_3020[40]; // @[OneHot.scala 39:40:@3603.4]
  assign _T_3128 = _T_3020[41]; // @[OneHot.scala 39:40:@3604.4]
  assign _T_3129 = _T_3020[42]; // @[OneHot.scala 39:40:@3605.4]
  assign _T_3130 = _T_3020[43]; // @[OneHot.scala 39:40:@3606.4]
  assign _T_3131 = _T_3020[44]; // @[OneHot.scala 39:40:@3607.4]
  assign _T_3132 = _T_3020[45]; // @[OneHot.scala 39:40:@3608.4]
  assign _T_3133 = _T_3020[46]; // @[OneHot.scala 39:40:@3609.4]
  assign _T_3134 = _T_3020[47]; // @[OneHot.scala 39:40:@3610.4]
  assign _T_3135 = _T_3020[48]; // @[OneHot.scala 39:40:@3611.4]
  assign _T_3136 = _T_3020[49]; // @[OneHot.scala 39:40:@3612.4]
  assign _T_3137 = _T_3020[50]; // @[OneHot.scala 39:40:@3613.4]
  assign _T_3138 = _T_3020[51]; // @[OneHot.scala 39:40:@3614.4]
  assign _T_3139 = _T_3020[52]; // @[OneHot.scala 39:40:@3615.4]
  assign _T_3140 = _T_3020[53]; // @[OneHot.scala 39:40:@3616.4]
  assign _T_3141 = _T_3020[54]; // @[OneHot.scala 39:40:@3617.4]
  assign _T_3142 = _T_3020[55]; // @[OneHot.scala 39:40:@3618.4]
  assign _T_3143 = _T_3020[56]; // @[OneHot.scala 39:40:@3619.4]
  assign _T_3144 = _T_3020[57]; // @[OneHot.scala 39:40:@3620.4]
  assign _T_3145 = _T_3020[58]; // @[OneHot.scala 39:40:@3621.4]
  assign _T_3146 = _T_3020[59]; // @[OneHot.scala 39:40:@3622.4]
  assign _T_3147 = _T_3020[60]; // @[OneHot.scala 39:40:@3623.4]
  assign _T_3148 = _T_3020[61]; // @[OneHot.scala 39:40:@3624.4]
  assign _T_3149 = _T_3020[62]; // @[OneHot.scala 39:40:@3625.4]
  assign _T_3215 = _T_3149 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@3627.4]
  assign _T_3216 = _T_3148 ? 6'h3d : _T_3215; // @[Mux.scala 31:69:@3628.4]
  assign _T_3217 = _T_3147 ? 6'h3c : _T_3216; // @[Mux.scala 31:69:@3629.4]
  assign _T_3218 = _T_3146 ? 6'h3b : _T_3217; // @[Mux.scala 31:69:@3630.4]
  assign _T_3219 = _T_3145 ? 6'h3a : _T_3218; // @[Mux.scala 31:69:@3631.4]
  assign _T_3220 = _T_3144 ? 6'h39 : _T_3219; // @[Mux.scala 31:69:@3632.4]
  assign _T_3221 = _T_3143 ? 6'h38 : _T_3220; // @[Mux.scala 31:69:@3633.4]
  assign _T_3222 = _T_3142 ? 6'h37 : _T_3221; // @[Mux.scala 31:69:@3634.4]
  assign _T_3223 = _T_3141 ? 6'h36 : _T_3222; // @[Mux.scala 31:69:@3635.4]
  assign _T_3224 = _T_3140 ? 6'h35 : _T_3223; // @[Mux.scala 31:69:@3636.4]
  assign _T_3225 = _T_3139 ? 6'h34 : _T_3224; // @[Mux.scala 31:69:@3637.4]
  assign _T_3226 = _T_3138 ? 6'h33 : _T_3225; // @[Mux.scala 31:69:@3638.4]
  assign _T_3227 = _T_3137 ? 6'h32 : _T_3226; // @[Mux.scala 31:69:@3639.4]
  assign _T_3228 = _T_3136 ? 6'h31 : _T_3227; // @[Mux.scala 31:69:@3640.4]
  assign _T_3229 = _T_3135 ? 6'h30 : _T_3228; // @[Mux.scala 31:69:@3641.4]
  assign _T_3230 = _T_3134 ? 6'h2f : _T_3229; // @[Mux.scala 31:69:@3642.4]
  assign _T_3231 = _T_3133 ? 6'h2e : _T_3230; // @[Mux.scala 31:69:@3643.4]
  assign _T_3232 = _T_3132 ? 6'h2d : _T_3231; // @[Mux.scala 31:69:@3644.4]
  assign _T_3233 = _T_3131 ? 6'h2c : _T_3232; // @[Mux.scala 31:69:@3645.4]
  assign _T_3234 = _T_3130 ? 6'h2b : _T_3233; // @[Mux.scala 31:69:@3646.4]
  assign _T_3235 = _T_3129 ? 6'h2a : _T_3234; // @[Mux.scala 31:69:@3647.4]
  assign _T_3236 = _T_3128 ? 6'h29 : _T_3235; // @[Mux.scala 31:69:@3648.4]
  assign _T_3237 = _T_3127 ? 6'h28 : _T_3236; // @[Mux.scala 31:69:@3649.4]
  assign _T_3238 = _T_3126 ? 6'h27 : _T_3237; // @[Mux.scala 31:69:@3650.4]
  assign _T_3239 = _T_3125 ? 6'h26 : _T_3238; // @[Mux.scala 31:69:@3651.4]
  assign _T_3240 = _T_3124 ? 6'h25 : _T_3239; // @[Mux.scala 31:69:@3652.4]
  assign _T_3241 = _T_3123 ? 6'h24 : _T_3240; // @[Mux.scala 31:69:@3653.4]
  assign _T_3242 = _T_3122 ? 6'h23 : _T_3241; // @[Mux.scala 31:69:@3654.4]
  assign _T_3243 = _T_3121 ? 6'h22 : _T_3242; // @[Mux.scala 31:69:@3655.4]
  assign _T_3244 = _T_3120 ? 6'h21 : _T_3243; // @[Mux.scala 31:69:@3656.4]
  assign _T_3245 = _T_3119 ? 6'h20 : _T_3244; // @[Mux.scala 31:69:@3657.4]
  assign _T_3246 = _T_3118 ? 6'h1f : _T_3245; // @[Mux.scala 31:69:@3658.4]
  assign _T_3247 = _T_3117 ? 6'h1e : _T_3246; // @[Mux.scala 31:69:@3659.4]
  assign _T_3248 = _T_3116 ? 6'h1d : _T_3247; // @[Mux.scala 31:69:@3660.4]
  assign _T_3249 = _T_3115 ? 6'h1c : _T_3248; // @[Mux.scala 31:69:@3661.4]
  assign _T_3250 = _T_3114 ? 6'h1b : _T_3249; // @[Mux.scala 31:69:@3662.4]
  assign _T_3251 = _T_3113 ? 6'h1a : _T_3250; // @[Mux.scala 31:69:@3663.4]
  assign _T_3252 = _T_3112 ? 6'h19 : _T_3251; // @[Mux.scala 31:69:@3664.4]
  assign _T_3253 = _T_3111 ? 6'h18 : _T_3252; // @[Mux.scala 31:69:@3665.4]
  assign _T_3254 = _T_3110 ? 6'h17 : _T_3253; // @[Mux.scala 31:69:@3666.4]
  assign _T_3255 = _T_3109 ? 6'h16 : _T_3254; // @[Mux.scala 31:69:@3667.4]
  assign _T_3256 = _T_3108 ? 6'h15 : _T_3255; // @[Mux.scala 31:69:@3668.4]
  assign _T_3257 = _T_3107 ? 6'h14 : _T_3256; // @[Mux.scala 31:69:@3669.4]
  assign _T_3258 = _T_3106 ? 6'h13 : _T_3257; // @[Mux.scala 31:69:@3670.4]
  assign _T_3259 = _T_3105 ? 6'h12 : _T_3258; // @[Mux.scala 31:69:@3671.4]
  assign _T_3260 = _T_3104 ? 6'h11 : _T_3259; // @[Mux.scala 31:69:@3672.4]
  assign _T_3261 = _T_3103 ? 6'h10 : _T_3260; // @[Mux.scala 31:69:@3673.4]
  assign _T_3262 = _T_3102 ? 6'hf : _T_3261; // @[Mux.scala 31:69:@3674.4]
  assign _T_3263 = _T_3101 ? 6'he : _T_3262; // @[Mux.scala 31:69:@3675.4]
  assign _T_3264 = _T_3100 ? 6'hd : _T_3263; // @[Mux.scala 31:69:@3676.4]
  assign _T_3265 = _T_3099 ? 6'hc : _T_3264; // @[Mux.scala 31:69:@3677.4]
  assign _T_3266 = _T_3098 ? 6'hb : _T_3265; // @[Mux.scala 31:69:@3678.4]
  assign _T_3267 = _T_3097 ? 6'ha : _T_3266; // @[Mux.scala 31:69:@3679.4]
  assign _T_3268 = _T_3096 ? 6'h9 : _T_3267; // @[Mux.scala 31:69:@3680.4]
  assign _T_3269 = _T_3095 ? 6'h8 : _T_3268; // @[Mux.scala 31:69:@3681.4]
  assign _T_3270 = _T_3094 ? 6'h7 : _T_3269; // @[Mux.scala 31:69:@3682.4]
  assign _T_3271 = _T_3093 ? 6'h6 : _T_3270; // @[Mux.scala 31:69:@3683.4]
  assign _T_3272 = _T_3092 ? 6'h5 : _T_3271; // @[Mux.scala 31:69:@3684.4]
  assign _T_3273 = _T_3091 ? 6'h4 : _T_3272; // @[Mux.scala 31:69:@3685.4]
  assign _T_3274 = _T_3090 ? 6'h3 : _T_3273; // @[Mux.scala 31:69:@3686.4]
  assign _T_3275 = _T_3089 ? 6'h2 : _T_3274; // @[Mux.scala 31:69:@3687.4]
  assign _T_3276 = _T_3088 ? 6'h1 : _T_3275; // @[Mux.scala 31:69:@3688.4]
  assign _T_3277 = _T_3087 ? 6'h0 : _T_3276; // @[Mux.scala 31:69:@3689.4]
  assign _T_3278 = _T_3022 ? fb_reg_lfsr : _T_3277; // @[BTB.scala 196:8:@3690.4]
  assign feedback_idx = _T_2925 ? _T_2956 : _T_3278; // @[BTB.scala 195:26:@3691.4]
  assign _GEN_9 = 6'h0 == feedback_idx ? 1'h1 : btb_valid_0; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_10 = 6'h1 == feedback_idx ? 1'h1 : btb_valid_1; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_11 = 6'h2 == feedback_idx ? 1'h1 : btb_valid_2; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_12 = 6'h3 == feedback_idx ? 1'h1 : btb_valid_3; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_13 = 6'h4 == feedback_idx ? 1'h1 : btb_valid_4; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_14 = 6'h5 == feedback_idx ? 1'h1 : btb_valid_5; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_15 = 6'h6 == feedback_idx ? 1'h1 : btb_valid_6; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_16 = 6'h7 == feedback_idx ? 1'h1 : btb_valid_7; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_17 = 6'h8 == feedback_idx ? 1'h1 : btb_valid_8; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_18 = 6'h9 == feedback_idx ? 1'h1 : btb_valid_9; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_19 = 6'ha == feedback_idx ? 1'h1 : btb_valid_10; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_20 = 6'hb == feedback_idx ? 1'h1 : btb_valid_11; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_21 = 6'hc == feedback_idx ? 1'h1 : btb_valid_12; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_22 = 6'hd == feedback_idx ? 1'h1 : btb_valid_13; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_23 = 6'he == feedback_idx ? 1'h1 : btb_valid_14; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_24 = 6'hf == feedback_idx ? 1'h1 : btb_valid_15; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_25 = 6'h10 == feedback_idx ? 1'h1 : btb_valid_16; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_26 = 6'h11 == feedback_idx ? 1'h1 : btb_valid_17; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_27 = 6'h12 == feedback_idx ? 1'h1 : btb_valid_18; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_28 = 6'h13 == feedback_idx ? 1'h1 : btb_valid_19; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_29 = 6'h14 == feedback_idx ? 1'h1 : btb_valid_20; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_30 = 6'h15 == feedback_idx ? 1'h1 : btb_valid_21; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_31 = 6'h16 == feedback_idx ? 1'h1 : btb_valid_22; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_32 = 6'h17 == feedback_idx ? 1'h1 : btb_valid_23; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_33 = 6'h18 == feedback_idx ? 1'h1 : btb_valid_24; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_34 = 6'h19 == feedback_idx ? 1'h1 : btb_valid_25; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_35 = 6'h1a == feedback_idx ? 1'h1 : btb_valid_26; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_36 = 6'h1b == feedback_idx ? 1'h1 : btb_valid_27; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_37 = 6'h1c == feedback_idx ? 1'h1 : btb_valid_28; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_38 = 6'h1d == feedback_idx ? 1'h1 : btb_valid_29; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_39 = 6'h1e == feedback_idx ? 1'h1 : btb_valid_30; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_40 = 6'h1f == feedback_idx ? 1'h1 : btb_valid_31; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_41 = 6'h20 == feedback_idx ? 1'h1 : btb_valid_32; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_42 = 6'h21 == feedback_idx ? 1'h1 : btb_valid_33; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_43 = 6'h22 == feedback_idx ? 1'h1 : btb_valid_34; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_44 = 6'h23 == feedback_idx ? 1'h1 : btb_valid_35; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_45 = 6'h24 == feedback_idx ? 1'h1 : btb_valid_36; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_46 = 6'h25 == feedback_idx ? 1'h1 : btb_valid_37; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_47 = 6'h26 == feedback_idx ? 1'h1 : btb_valid_38; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_48 = 6'h27 == feedback_idx ? 1'h1 : btb_valid_39; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_49 = 6'h28 == feedback_idx ? 1'h1 : btb_valid_40; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_50 = 6'h29 == feedback_idx ? 1'h1 : btb_valid_41; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_51 = 6'h2a == feedback_idx ? 1'h1 : btb_valid_42; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_52 = 6'h2b == feedback_idx ? 1'h1 : btb_valid_43; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_53 = 6'h2c == feedback_idx ? 1'h1 : btb_valid_44; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_54 = 6'h2d == feedback_idx ? 1'h1 : btb_valid_45; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_55 = 6'h2e == feedback_idx ? 1'h1 : btb_valid_46; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_56 = 6'h2f == feedback_idx ? 1'h1 : btb_valid_47; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_57 = 6'h30 == feedback_idx ? 1'h1 : btb_valid_48; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_58 = 6'h31 == feedback_idx ? 1'h1 : btb_valid_49; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_59 = 6'h32 == feedback_idx ? 1'h1 : btb_valid_50; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_60 = 6'h33 == feedback_idx ? 1'h1 : btb_valid_51; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_61 = 6'h34 == feedback_idx ? 1'h1 : btb_valid_52; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_62 = 6'h35 == feedback_idx ? 1'h1 : btb_valid_53; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_63 = 6'h36 == feedback_idx ? 1'h1 : btb_valid_54; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_64 = 6'h37 == feedback_idx ? 1'h1 : btb_valid_55; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_65 = 6'h38 == feedback_idx ? 1'h1 : btb_valid_56; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_66 = 6'h39 == feedback_idx ? 1'h1 : btb_valid_57; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_67 = 6'h3a == feedback_idx ? 1'h1 : btb_valid_58; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_68 = 6'h3b == feedback_idx ? 1'h1 : btb_valid_59; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_69 = 6'h3c == feedback_idx ? 1'h1 : btb_valid_60; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_70 = 6'h3d == feedback_idx ? 1'h1 : btb_valid_61; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_71 = 6'h3e == feedback_idx ? 1'h1 : btb_valid_62; // @[BTB.scala 201:32:@3697.8]
  assign _GEN_72 = 6'h3f == feedback_idx ? 1'h1 : btb_valid_63; // @[BTB.scala 201:32:@3697.8]
  assign _T_3285 = fb_reg_btb_type == 2'h2; // @[BTB.scala 203:51:@3702.10]
  assign _GEN_73 = 6'h0 == feedback_idx ? _T_3285 : btb_valid_0; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_74 = 6'h1 == feedback_idx ? _T_3285 : btb_valid_1; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_75 = 6'h2 == feedback_idx ? _T_3285 : btb_valid_2; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_76 = 6'h3 == feedback_idx ? _T_3285 : btb_valid_3; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_77 = 6'h4 == feedback_idx ? _T_3285 : btb_valid_4; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_78 = 6'h5 == feedback_idx ? _T_3285 : btb_valid_5; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_79 = 6'h6 == feedback_idx ? _T_3285 : btb_valid_6; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_80 = 6'h7 == feedback_idx ? _T_3285 : btb_valid_7; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_81 = 6'h8 == feedback_idx ? _T_3285 : btb_valid_8; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_82 = 6'h9 == feedback_idx ? _T_3285 : btb_valid_9; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_83 = 6'ha == feedback_idx ? _T_3285 : btb_valid_10; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_84 = 6'hb == feedback_idx ? _T_3285 : btb_valid_11; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_85 = 6'hc == feedback_idx ? _T_3285 : btb_valid_12; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_86 = 6'hd == feedback_idx ? _T_3285 : btb_valid_13; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_87 = 6'he == feedback_idx ? _T_3285 : btb_valid_14; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_88 = 6'hf == feedback_idx ? _T_3285 : btb_valid_15; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_89 = 6'h10 == feedback_idx ? _T_3285 : btb_valid_16; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_90 = 6'h11 == feedback_idx ? _T_3285 : btb_valid_17; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_91 = 6'h12 == feedback_idx ? _T_3285 : btb_valid_18; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_92 = 6'h13 == feedback_idx ? _T_3285 : btb_valid_19; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_93 = 6'h14 == feedback_idx ? _T_3285 : btb_valid_20; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_94 = 6'h15 == feedback_idx ? _T_3285 : btb_valid_21; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_95 = 6'h16 == feedback_idx ? _T_3285 : btb_valid_22; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_96 = 6'h17 == feedback_idx ? _T_3285 : btb_valid_23; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_97 = 6'h18 == feedback_idx ? _T_3285 : btb_valid_24; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_98 = 6'h19 == feedback_idx ? _T_3285 : btb_valid_25; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_99 = 6'h1a == feedback_idx ? _T_3285 : btb_valid_26; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_100 = 6'h1b == feedback_idx ? _T_3285 : btb_valid_27; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_101 = 6'h1c == feedback_idx ? _T_3285 : btb_valid_28; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_102 = 6'h1d == feedback_idx ? _T_3285 : btb_valid_29; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_103 = 6'h1e == feedback_idx ? _T_3285 : btb_valid_30; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_104 = 6'h1f == feedback_idx ? _T_3285 : btb_valid_31; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_105 = 6'h20 == feedback_idx ? _T_3285 : btb_valid_32; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_106 = 6'h21 == feedback_idx ? _T_3285 : btb_valid_33; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_107 = 6'h22 == feedback_idx ? _T_3285 : btb_valid_34; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_108 = 6'h23 == feedback_idx ? _T_3285 : btb_valid_35; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_109 = 6'h24 == feedback_idx ? _T_3285 : btb_valid_36; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_110 = 6'h25 == feedback_idx ? _T_3285 : btb_valid_37; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_111 = 6'h26 == feedback_idx ? _T_3285 : btb_valid_38; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_112 = 6'h27 == feedback_idx ? _T_3285 : btb_valid_39; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_113 = 6'h28 == feedback_idx ? _T_3285 : btb_valid_40; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_114 = 6'h29 == feedback_idx ? _T_3285 : btb_valid_41; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_115 = 6'h2a == feedback_idx ? _T_3285 : btb_valid_42; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_116 = 6'h2b == feedback_idx ? _T_3285 : btb_valid_43; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_117 = 6'h2c == feedback_idx ? _T_3285 : btb_valid_44; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_118 = 6'h2d == feedback_idx ? _T_3285 : btb_valid_45; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_119 = 6'h2e == feedback_idx ? _T_3285 : btb_valid_46; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_120 = 6'h2f == feedback_idx ? _T_3285 : btb_valid_47; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_121 = 6'h30 == feedback_idx ? _T_3285 : btb_valid_48; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_122 = 6'h31 == feedback_idx ? _T_3285 : btb_valid_49; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_123 = 6'h32 == feedback_idx ? _T_3285 : btb_valid_50; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_124 = 6'h33 == feedback_idx ? _T_3285 : btb_valid_51; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_125 = 6'h34 == feedback_idx ? _T_3285 : btb_valid_52; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_126 = 6'h35 == feedback_idx ? _T_3285 : btb_valid_53; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_127 = 6'h36 == feedback_idx ? _T_3285 : btb_valid_54; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_128 = 6'h37 == feedback_idx ? _T_3285 : btb_valid_55; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_129 = 6'h38 == feedback_idx ? _T_3285 : btb_valid_56; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_130 = 6'h39 == feedback_idx ? _T_3285 : btb_valid_57; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_131 = 6'h3a == feedback_idx ? _T_3285 : btb_valid_58; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_132 = 6'h3b == feedback_idx ? _T_3285 : btb_valid_59; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_133 = 6'h3c == feedback_idx ? _T_3285 : btb_valid_60; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_134 = 6'h3d == feedback_idx ? _T_3285 : btb_valid_61; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_135 = 6'h3e == feedback_idx ? _T_3285 : btb_valid_62; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_136 = 6'h3f == feedback_idx ? _T_3285 : btb_valid_63; // @[BTB.scala 203:32:@3703.10]
  assign _GEN_137 = _T_2925 ? _GEN_73 : btb_valid_0; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_138 = _T_2925 ? _GEN_74 : btb_valid_1; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_139 = _T_2925 ? _GEN_75 : btb_valid_2; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_140 = _T_2925 ? _GEN_76 : btb_valid_3; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_141 = _T_2925 ? _GEN_77 : btb_valid_4; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_142 = _T_2925 ? _GEN_78 : btb_valid_5; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_143 = _T_2925 ? _GEN_79 : btb_valid_6; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_144 = _T_2925 ? _GEN_80 : btb_valid_7; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_145 = _T_2925 ? _GEN_81 : btb_valid_8; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_146 = _T_2925 ? _GEN_82 : btb_valid_9; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_147 = _T_2925 ? _GEN_83 : btb_valid_10; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_148 = _T_2925 ? _GEN_84 : btb_valid_11; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_149 = _T_2925 ? _GEN_85 : btb_valid_12; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_150 = _T_2925 ? _GEN_86 : btb_valid_13; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_151 = _T_2925 ? _GEN_87 : btb_valid_14; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_152 = _T_2925 ? _GEN_88 : btb_valid_15; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_153 = _T_2925 ? _GEN_89 : btb_valid_16; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_154 = _T_2925 ? _GEN_90 : btb_valid_17; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_155 = _T_2925 ? _GEN_91 : btb_valid_18; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_156 = _T_2925 ? _GEN_92 : btb_valid_19; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_157 = _T_2925 ? _GEN_93 : btb_valid_20; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_158 = _T_2925 ? _GEN_94 : btb_valid_21; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_159 = _T_2925 ? _GEN_95 : btb_valid_22; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_160 = _T_2925 ? _GEN_96 : btb_valid_23; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_161 = _T_2925 ? _GEN_97 : btb_valid_24; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_162 = _T_2925 ? _GEN_98 : btb_valid_25; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_163 = _T_2925 ? _GEN_99 : btb_valid_26; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_164 = _T_2925 ? _GEN_100 : btb_valid_27; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_165 = _T_2925 ? _GEN_101 : btb_valid_28; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_166 = _T_2925 ? _GEN_102 : btb_valid_29; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_167 = _T_2925 ? _GEN_103 : btb_valid_30; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_168 = _T_2925 ? _GEN_104 : btb_valid_31; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_169 = _T_2925 ? _GEN_105 : btb_valid_32; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_170 = _T_2925 ? _GEN_106 : btb_valid_33; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_171 = _T_2925 ? _GEN_107 : btb_valid_34; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_172 = _T_2925 ? _GEN_108 : btb_valid_35; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_173 = _T_2925 ? _GEN_109 : btb_valid_36; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_174 = _T_2925 ? _GEN_110 : btb_valid_37; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_175 = _T_2925 ? _GEN_111 : btb_valid_38; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_176 = _T_2925 ? _GEN_112 : btb_valid_39; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_177 = _T_2925 ? _GEN_113 : btb_valid_40; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_178 = _T_2925 ? _GEN_114 : btb_valid_41; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_179 = _T_2925 ? _GEN_115 : btb_valid_42; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_180 = _T_2925 ? _GEN_116 : btb_valid_43; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_181 = _T_2925 ? _GEN_117 : btb_valid_44; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_182 = _T_2925 ? _GEN_118 : btb_valid_45; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_183 = _T_2925 ? _GEN_119 : btb_valid_46; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_184 = _T_2925 ? _GEN_120 : btb_valid_47; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_185 = _T_2925 ? _GEN_121 : btb_valid_48; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_186 = _T_2925 ? _GEN_122 : btb_valid_49; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_187 = _T_2925 ? _GEN_123 : btb_valid_50; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_188 = _T_2925 ? _GEN_124 : btb_valid_51; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_189 = _T_2925 ? _GEN_125 : btb_valid_52; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_190 = _T_2925 ? _GEN_126 : btb_valid_53; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_191 = _T_2925 ? _GEN_127 : btb_valid_54; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_192 = _T_2925 ? _GEN_128 : btb_valid_55; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_193 = _T_2925 ? _GEN_129 : btb_valid_56; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_194 = _T_2925 ? _GEN_130 : btb_valid_57; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_195 = _T_2925 ? _GEN_131 : btb_valid_58; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_196 = _T_2925 ? _GEN_132 : btb_valid_59; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_197 = _T_2925 ? _GEN_133 : btb_valid_60; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_198 = _T_2925 ? _GEN_134 : btb_valid_61; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_199 = _T_2925 ? _GEN_135 : btb_valid_62; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_200 = _T_2925 ? _GEN_136 : btb_valid_63; // @[BTB.scala 202:32:@3701.8]
  assign _GEN_201 = fb_reg_redirect ? _GEN_9 : _GEN_137; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_202 = fb_reg_redirect ? _GEN_10 : _GEN_138; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_203 = fb_reg_redirect ? _GEN_11 : _GEN_139; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_204 = fb_reg_redirect ? _GEN_12 : _GEN_140; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_205 = fb_reg_redirect ? _GEN_13 : _GEN_141; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_206 = fb_reg_redirect ? _GEN_14 : _GEN_142; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_207 = fb_reg_redirect ? _GEN_15 : _GEN_143; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_208 = fb_reg_redirect ? _GEN_16 : _GEN_144; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_209 = fb_reg_redirect ? _GEN_17 : _GEN_145; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_210 = fb_reg_redirect ? _GEN_18 : _GEN_146; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_211 = fb_reg_redirect ? _GEN_19 : _GEN_147; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_212 = fb_reg_redirect ? _GEN_20 : _GEN_148; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_213 = fb_reg_redirect ? _GEN_21 : _GEN_149; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_214 = fb_reg_redirect ? _GEN_22 : _GEN_150; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_215 = fb_reg_redirect ? _GEN_23 : _GEN_151; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_216 = fb_reg_redirect ? _GEN_24 : _GEN_152; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_217 = fb_reg_redirect ? _GEN_25 : _GEN_153; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_218 = fb_reg_redirect ? _GEN_26 : _GEN_154; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_219 = fb_reg_redirect ? _GEN_27 : _GEN_155; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_220 = fb_reg_redirect ? _GEN_28 : _GEN_156; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_221 = fb_reg_redirect ? _GEN_29 : _GEN_157; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_222 = fb_reg_redirect ? _GEN_30 : _GEN_158; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_223 = fb_reg_redirect ? _GEN_31 : _GEN_159; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_224 = fb_reg_redirect ? _GEN_32 : _GEN_160; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_225 = fb_reg_redirect ? _GEN_33 : _GEN_161; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_226 = fb_reg_redirect ? _GEN_34 : _GEN_162; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_227 = fb_reg_redirect ? _GEN_35 : _GEN_163; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_228 = fb_reg_redirect ? _GEN_36 : _GEN_164; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_229 = fb_reg_redirect ? _GEN_37 : _GEN_165; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_230 = fb_reg_redirect ? _GEN_38 : _GEN_166; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_231 = fb_reg_redirect ? _GEN_39 : _GEN_167; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_232 = fb_reg_redirect ? _GEN_40 : _GEN_168; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_233 = fb_reg_redirect ? _GEN_41 : _GEN_169; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_234 = fb_reg_redirect ? _GEN_42 : _GEN_170; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_235 = fb_reg_redirect ? _GEN_43 : _GEN_171; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_236 = fb_reg_redirect ? _GEN_44 : _GEN_172; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_237 = fb_reg_redirect ? _GEN_45 : _GEN_173; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_238 = fb_reg_redirect ? _GEN_46 : _GEN_174; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_239 = fb_reg_redirect ? _GEN_47 : _GEN_175; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_240 = fb_reg_redirect ? _GEN_48 : _GEN_176; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_241 = fb_reg_redirect ? _GEN_49 : _GEN_177; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_242 = fb_reg_redirect ? _GEN_50 : _GEN_178; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_243 = fb_reg_redirect ? _GEN_51 : _GEN_179; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_244 = fb_reg_redirect ? _GEN_52 : _GEN_180; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_245 = fb_reg_redirect ? _GEN_53 : _GEN_181; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_246 = fb_reg_redirect ? _GEN_54 : _GEN_182; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_247 = fb_reg_redirect ? _GEN_55 : _GEN_183; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_248 = fb_reg_redirect ? _GEN_56 : _GEN_184; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_249 = fb_reg_redirect ? _GEN_57 : _GEN_185; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_250 = fb_reg_redirect ? _GEN_58 : _GEN_186; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_251 = fb_reg_redirect ? _GEN_59 : _GEN_187; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_252 = fb_reg_redirect ? _GEN_60 : _GEN_188; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_253 = fb_reg_redirect ? _GEN_61 : _GEN_189; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_254 = fb_reg_redirect ? _GEN_62 : _GEN_190; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_255 = fb_reg_redirect ? _GEN_63 : _GEN_191; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_256 = fb_reg_redirect ? _GEN_64 : _GEN_192; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_257 = fb_reg_redirect ? _GEN_65 : _GEN_193; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_258 = fb_reg_redirect ? _GEN_66 : _GEN_194; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_259 = fb_reg_redirect ? _GEN_67 : _GEN_195; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_260 = fb_reg_redirect ? _GEN_68 : _GEN_196; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_261 = fb_reg_redirect ? _GEN_69 : _GEN_197; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_262 = fb_reg_redirect ? _GEN_70 : _GEN_198; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_263 = fb_reg_redirect ? _GEN_71 : _GEN_199; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_264 = fb_reg_redirect ? _GEN_72 : _GEN_200; // @[BTB.scala 200:28:@3696.6]
  assign _GEN_265 = 6'h0 == feedback_idx ? fb_reg_pc : btb_pc_0; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_266 = 6'h1 == feedback_idx ? fb_reg_pc : btb_pc_1; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_267 = 6'h2 == feedback_idx ? fb_reg_pc : btb_pc_2; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_268 = 6'h3 == feedback_idx ? fb_reg_pc : btb_pc_3; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_269 = 6'h4 == feedback_idx ? fb_reg_pc : btb_pc_4; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_270 = 6'h5 == feedback_idx ? fb_reg_pc : btb_pc_5; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_271 = 6'h6 == feedback_idx ? fb_reg_pc : btb_pc_6; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_272 = 6'h7 == feedback_idx ? fb_reg_pc : btb_pc_7; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_273 = 6'h8 == feedback_idx ? fb_reg_pc : btb_pc_8; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_274 = 6'h9 == feedback_idx ? fb_reg_pc : btb_pc_9; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_275 = 6'ha == feedback_idx ? fb_reg_pc : btb_pc_10; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_276 = 6'hb == feedback_idx ? fb_reg_pc : btb_pc_11; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_277 = 6'hc == feedback_idx ? fb_reg_pc : btb_pc_12; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_278 = 6'hd == feedback_idx ? fb_reg_pc : btb_pc_13; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_279 = 6'he == feedback_idx ? fb_reg_pc : btb_pc_14; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_280 = 6'hf == feedback_idx ? fb_reg_pc : btb_pc_15; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_281 = 6'h10 == feedback_idx ? fb_reg_pc : btb_pc_16; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_282 = 6'h11 == feedback_idx ? fb_reg_pc : btb_pc_17; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_283 = 6'h12 == feedback_idx ? fb_reg_pc : btb_pc_18; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_284 = 6'h13 == feedback_idx ? fb_reg_pc : btb_pc_19; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_285 = 6'h14 == feedback_idx ? fb_reg_pc : btb_pc_20; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_286 = 6'h15 == feedback_idx ? fb_reg_pc : btb_pc_21; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_287 = 6'h16 == feedback_idx ? fb_reg_pc : btb_pc_22; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_288 = 6'h17 == feedback_idx ? fb_reg_pc : btb_pc_23; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_289 = 6'h18 == feedback_idx ? fb_reg_pc : btb_pc_24; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_290 = 6'h19 == feedback_idx ? fb_reg_pc : btb_pc_25; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_291 = 6'h1a == feedback_idx ? fb_reg_pc : btb_pc_26; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_292 = 6'h1b == feedback_idx ? fb_reg_pc : btb_pc_27; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_293 = 6'h1c == feedback_idx ? fb_reg_pc : btb_pc_28; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_294 = 6'h1d == feedback_idx ? fb_reg_pc : btb_pc_29; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_295 = 6'h1e == feedback_idx ? fb_reg_pc : btb_pc_30; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_296 = 6'h1f == feedback_idx ? fb_reg_pc : btb_pc_31; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_297 = 6'h20 == feedback_idx ? fb_reg_pc : btb_pc_32; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_298 = 6'h21 == feedback_idx ? fb_reg_pc : btb_pc_33; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_299 = 6'h22 == feedback_idx ? fb_reg_pc : btb_pc_34; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_300 = 6'h23 == feedback_idx ? fb_reg_pc : btb_pc_35; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_301 = 6'h24 == feedback_idx ? fb_reg_pc : btb_pc_36; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_302 = 6'h25 == feedback_idx ? fb_reg_pc : btb_pc_37; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_303 = 6'h26 == feedback_idx ? fb_reg_pc : btb_pc_38; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_304 = 6'h27 == feedback_idx ? fb_reg_pc : btb_pc_39; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_305 = 6'h28 == feedback_idx ? fb_reg_pc : btb_pc_40; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_306 = 6'h29 == feedback_idx ? fb_reg_pc : btb_pc_41; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_307 = 6'h2a == feedback_idx ? fb_reg_pc : btb_pc_42; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_308 = 6'h2b == feedback_idx ? fb_reg_pc : btb_pc_43; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_309 = 6'h2c == feedback_idx ? fb_reg_pc : btb_pc_44; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_310 = 6'h2d == feedback_idx ? fb_reg_pc : btb_pc_45; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_311 = 6'h2e == feedback_idx ? fb_reg_pc : btb_pc_46; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_312 = 6'h2f == feedback_idx ? fb_reg_pc : btb_pc_47; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_313 = 6'h30 == feedback_idx ? fb_reg_pc : btb_pc_48; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_314 = 6'h31 == feedback_idx ? fb_reg_pc : btb_pc_49; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_315 = 6'h32 == feedback_idx ? fb_reg_pc : btb_pc_50; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_316 = 6'h33 == feedback_idx ? fb_reg_pc : btb_pc_51; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_317 = 6'h34 == feedback_idx ? fb_reg_pc : btb_pc_52; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_318 = 6'h35 == feedback_idx ? fb_reg_pc : btb_pc_53; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_319 = 6'h36 == feedback_idx ? fb_reg_pc : btb_pc_54; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_320 = 6'h37 == feedback_idx ? fb_reg_pc : btb_pc_55; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_321 = 6'h38 == feedback_idx ? fb_reg_pc : btb_pc_56; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_322 = 6'h39 == feedback_idx ? fb_reg_pc : btb_pc_57; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_323 = 6'h3a == feedback_idx ? fb_reg_pc : btb_pc_58; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_324 = 6'h3b == feedback_idx ? fb_reg_pc : btb_pc_59; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_325 = 6'h3c == feedback_idx ? fb_reg_pc : btb_pc_60; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_326 = 6'h3d == feedback_idx ? fb_reg_pc : btb_pc_61; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_327 = 6'h3e == feedback_idx ? fb_reg_pc : btb_pc_62; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_328 = 6'h3f == feedback_idx ? fb_reg_pc : btb_pc_63; // @[BTB.scala 206:33:@3706.8]
  assign _GEN_329 = 6'h0 == feedback_idx ? fb_reg_tgt : btb_tgt_0; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_330 = 6'h1 == feedback_idx ? fb_reg_tgt : btb_tgt_1; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_331 = 6'h2 == feedback_idx ? fb_reg_tgt : btb_tgt_2; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_332 = 6'h3 == feedback_idx ? fb_reg_tgt : btb_tgt_3; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_333 = 6'h4 == feedback_idx ? fb_reg_tgt : btb_tgt_4; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_334 = 6'h5 == feedback_idx ? fb_reg_tgt : btb_tgt_5; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_335 = 6'h6 == feedback_idx ? fb_reg_tgt : btb_tgt_6; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_336 = 6'h7 == feedback_idx ? fb_reg_tgt : btb_tgt_7; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_337 = 6'h8 == feedback_idx ? fb_reg_tgt : btb_tgt_8; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_338 = 6'h9 == feedback_idx ? fb_reg_tgt : btb_tgt_9; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_339 = 6'ha == feedback_idx ? fb_reg_tgt : btb_tgt_10; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_340 = 6'hb == feedback_idx ? fb_reg_tgt : btb_tgt_11; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_341 = 6'hc == feedback_idx ? fb_reg_tgt : btb_tgt_12; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_342 = 6'hd == feedback_idx ? fb_reg_tgt : btb_tgt_13; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_343 = 6'he == feedback_idx ? fb_reg_tgt : btb_tgt_14; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_344 = 6'hf == feedback_idx ? fb_reg_tgt : btb_tgt_15; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_345 = 6'h10 == feedback_idx ? fb_reg_tgt : btb_tgt_16; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_346 = 6'h11 == feedback_idx ? fb_reg_tgt : btb_tgt_17; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_347 = 6'h12 == feedback_idx ? fb_reg_tgt : btb_tgt_18; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_348 = 6'h13 == feedback_idx ? fb_reg_tgt : btb_tgt_19; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_349 = 6'h14 == feedback_idx ? fb_reg_tgt : btb_tgt_20; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_350 = 6'h15 == feedback_idx ? fb_reg_tgt : btb_tgt_21; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_351 = 6'h16 == feedback_idx ? fb_reg_tgt : btb_tgt_22; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_352 = 6'h17 == feedback_idx ? fb_reg_tgt : btb_tgt_23; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_353 = 6'h18 == feedback_idx ? fb_reg_tgt : btb_tgt_24; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_354 = 6'h19 == feedback_idx ? fb_reg_tgt : btb_tgt_25; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_355 = 6'h1a == feedback_idx ? fb_reg_tgt : btb_tgt_26; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_356 = 6'h1b == feedback_idx ? fb_reg_tgt : btb_tgt_27; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_357 = 6'h1c == feedback_idx ? fb_reg_tgt : btb_tgt_28; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_358 = 6'h1d == feedback_idx ? fb_reg_tgt : btb_tgt_29; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_359 = 6'h1e == feedback_idx ? fb_reg_tgt : btb_tgt_30; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_360 = 6'h1f == feedback_idx ? fb_reg_tgt : btb_tgt_31; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_361 = 6'h20 == feedback_idx ? fb_reg_tgt : btb_tgt_32; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_362 = 6'h21 == feedback_idx ? fb_reg_tgt : btb_tgt_33; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_363 = 6'h22 == feedback_idx ? fb_reg_tgt : btb_tgt_34; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_364 = 6'h23 == feedback_idx ? fb_reg_tgt : btb_tgt_35; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_365 = 6'h24 == feedback_idx ? fb_reg_tgt : btb_tgt_36; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_366 = 6'h25 == feedback_idx ? fb_reg_tgt : btb_tgt_37; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_367 = 6'h26 == feedback_idx ? fb_reg_tgt : btb_tgt_38; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_368 = 6'h27 == feedback_idx ? fb_reg_tgt : btb_tgt_39; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_369 = 6'h28 == feedback_idx ? fb_reg_tgt : btb_tgt_40; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_370 = 6'h29 == feedback_idx ? fb_reg_tgt : btb_tgt_41; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_371 = 6'h2a == feedback_idx ? fb_reg_tgt : btb_tgt_42; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_372 = 6'h2b == feedback_idx ? fb_reg_tgt : btb_tgt_43; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_373 = 6'h2c == feedback_idx ? fb_reg_tgt : btb_tgt_44; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_374 = 6'h2d == feedback_idx ? fb_reg_tgt : btb_tgt_45; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_375 = 6'h2e == feedback_idx ? fb_reg_tgt : btb_tgt_46; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_376 = 6'h2f == feedback_idx ? fb_reg_tgt : btb_tgt_47; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_377 = 6'h30 == feedback_idx ? fb_reg_tgt : btb_tgt_48; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_378 = 6'h31 == feedback_idx ? fb_reg_tgt : btb_tgt_49; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_379 = 6'h32 == feedback_idx ? fb_reg_tgt : btb_tgt_50; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_380 = 6'h33 == feedback_idx ? fb_reg_tgt : btb_tgt_51; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_381 = 6'h34 == feedback_idx ? fb_reg_tgt : btb_tgt_52; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_382 = 6'h35 == feedback_idx ? fb_reg_tgt : btb_tgt_53; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_383 = 6'h36 == feedback_idx ? fb_reg_tgt : btb_tgt_54; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_384 = 6'h37 == feedback_idx ? fb_reg_tgt : btb_tgt_55; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_385 = 6'h38 == feedback_idx ? fb_reg_tgt : btb_tgt_56; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_386 = 6'h39 == feedback_idx ? fb_reg_tgt : btb_tgt_57; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_387 = 6'h3a == feedback_idx ? fb_reg_tgt : btb_tgt_58; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_388 = 6'h3b == feedback_idx ? fb_reg_tgt : btb_tgt_59; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_389 = 6'h3c == feedback_idx ? fb_reg_tgt : btb_tgt_60; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_390 = 6'h3d == feedback_idx ? fb_reg_tgt : btb_tgt_61; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_391 = 6'h3e == feedback_idx ? fb_reg_tgt : btb_tgt_62; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_392 = 6'h3f == feedback_idx ? fb_reg_tgt : btb_tgt_63; // @[BTB.scala 207:33:@3707.8]
  assign _GEN_393 = 6'h0 == feedback_idx ? fb_reg_btb_type : btb_bj_type_0; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_394 = 6'h1 == feedback_idx ? fb_reg_btb_type : btb_bj_type_1; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_395 = 6'h2 == feedback_idx ? fb_reg_btb_type : btb_bj_type_2; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_396 = 6'h3 == feedback_idx ? fb_reg_btb_type : btb_bj_type_3; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_397 = 6'h4 == feedback_idx ? fb_reg_btb_type : btb_bj_type_4; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_398 = 6'h5 == feedback_idx ? fb_reg_btb_type : btb_bj_type_5; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_399 = 6'h6 == feedback_idx ? fb_reg_btb_type : btb_bj_type_6; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_400 = 6'h7 == feedback_idx ? fb_reg_btb_type : btb_bj_type_7; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_401 = 6'h8 == feedback_idx ? fb_reg_btb_type : btb_bj_type_8; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_402 = 6'h9 == feedback_idx ? fb_reg_btb_type : btb_bj_type_9; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_403 = 6'ha == feedback_idx ? fb_reg_btb_type : btb_bj_type_10; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_404 = 6'hb == feedback_idx ? fb_reg_btb_type : btb_bj_type_11; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_405 = 6'hc == feedback_idx ? fb_reg_btb_type : btb_bj_type_12; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_406 = 6'hd == feedback_idx ? fb_reg_btb_type : btb_bj_type_13; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_407 = 6'he == feedback_idx ? fb_reg_btb_type : btb_bj_type_14; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_408 = 6'hf == feedback_idx ? fb_reg_btb_type : btb_bj_type_15; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_409 = 6'h10 == feedback_idx ? fb_reg_btb_type : btb_bj_type_16; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_410 = 6'h11 == feedback_idx ? fb_reg_btb_type : btb_bj_type_17; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_411 = 6'h12 == feedback_idx ? fb_reg_btb_type : btb_bj_type_18; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_412 = 6'h13 == feedback_idx ? fb_reg_btb_type : btb_bj_type_19; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_413 = 6'h14 == feedback_idx ? fb_reg_btb_type : btb_bj_type_20; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_414 = 6'h15 == feedback_idx ? fb_reg_btb_type : btb_bj_type_21; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_415 = 6'h16 == feedback_idx ? fb_reg_btb_type : btb_bj_type_22; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_416 = 6'h17 == feedback_idx ? fb_reg_btb_type : btb_bj_type_23; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_417 = 6'h18 == feedback_idx ? fb_reg_btb_type : btb_bj_type_24; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_418 = 6'h19 == feedback_idx ? fb_reg_btb_type : btb_bj_type_25; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_419 = 6'h1a == feedback_idx ? fb_reg_btb_type : btb_bj_type_26; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_420 = 6'h1b == feedback_idx ? fb_reg_btb_type : btb_bj_type_27; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_421 = 6'h1c == feedback_idx ? fb_reg_btb_type : btb_bj_type_28; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_422 = 6'h1d == feedback_idx ? fb_reg_btb_type : btb_bj_type_29; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_423 = 6'h1e == feedback_idx ? fb_reg_btb_type : btb_bj_type_30; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_424 = 6'h1f == feedback_idx ? fb_reg_btb_type : btb_bj_type_31; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_425 = 6'h20 == feedback_idx ? fb_reg_btb_type : btb_bj_type_32; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_426 = 6'h21 == feedback_idx ? fb_reg_btb_type : btb_bj_type_33; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_427 = 6'h22 == feedback_idx ? fb_reg_btb_type : btb_bj_type_34; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_428 = 6'h23 == feedback_idx ? fb_reg_btb_type : btb_bj_type_35; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_429 = 6'h24 == feedback_idx ? fb_reg_btb_type : btb_bj_type_36; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_430 = 6'h25 == feedback_idx ? fb_reg_btb_type : btb_bj_type_37; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_431 = 6'h26 == feedback_idx ? fb_reg_btb_type : btb_bj_type_38; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_432 = 6'h27 == feedback_idx ? fb_reg_btb_type : btb_bj_type_39; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_433 = 6'h28 == feedback_idx ? fb_reg_btb_type : btb_bj_type_40; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_434 = 6'h29 == feedback_idx ? fb_reg_btb_type : btb_bj_type_41; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_435 = 6'h2a == feedback_idx ? fb_reg_btb_type : btb_bj_type_42; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_436 = 6'h2b == feedback_idx ? fb_reg_btb_type : btb_bj_type_43; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_437 = 6'h2c == feedback_idx ? fb_reg_btb_type : btb_bj_type_44; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_438 = 6'h2d == feedback_idx ? fb_reg_btb_type : btb_bj_type_45; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_439 = 6'h2e == feedback_idx ? fb_reg_btb_type : btb_bj_type_46; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_440 = 6'h2f == feedback_idx ? fb_reg_btb_type : btb_bj_type_47; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_441 = 6'h30 == feedback_idx ? fb_reg_btb_type : btb_bj_type_48; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_442 = 6'h31 == feedback_idx ? fb_reg_btb_type : btb_bj_type_49; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_443 = 6'h32 == feedback_idx ? fb_reg_btb_type : btb_bj_type_50; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_444 = 6'h33 == feedback_idx ? fb_reg_btb_type : btb_bj_type_51; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_445 = 6'h34 == feedback_idx ? fb_reg_btb_type : btb_bj_type_52; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_446 = 6'h35 == feedback_idx ? fb_reg_btb_type : btb_bj_type_53; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_447 = 6'h36 == feedback_idx ? fb_reg_btb_type : btb_bj_type_54; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_448 = 6'h37 == feedback_idx ? fb_reg_btb_type : btb_bj_type_55; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_449 = 6'h38 == feedback_idx ? fb_reg_btb_type : btb_bj_type_56; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_450 = 6'h39 == feedback_idx ? fb_reg_btb_type : btb_bj_type_57; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_451 = 6'h3a == feedback_idx ? fb_reg_btb_type : btb_bj_type_58; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_452 = 6'h3b == feedback_idx ? fb_reg_btb_type : btb_bj_type_59; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_453 = 6'h3c == feedback_idx ? fb_reg_btb_type : btb_bj_type_60; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_454 = 6'h3d == feedback_idx ? fb_reg_btb_type : btb_bj_type_61; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_455 = 6'h3e == feedback_idx ? fb_reg_btb_type : btb_bj_type_62; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_456 = 6'h3f == feedback_idx ? fb_reg_btb_type : btb_bj_type_63; // @[BTB.scala 208:33:@3708.8]
  assign _GEN_457 = fb_reg_redirect ? _GEN_265 : btb_pc_0; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_458 = fb_reg_redirect ? _GEN_266 : btb_pc_1; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_459 = fb_reg_redirect ? _GEN_267 : btb_pc_2; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_460 = fb_reg_redirect ? _GEN_268 : btb_pc_3; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_461 = fb_reg_redirect ? _GEN_269 : btb_pc_4; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_462 = fb_reg_redirect ? _GEN_270 : btb_pc_5; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_463 = fb_reg_redirect ? _GEN_271 : btb_pc_6; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_464 = fb_reg_redirect ? _GEN_272 : btb_pc_7; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_465 = fb_reg_redirect ? _GEN_273 : btb_pc_8; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_466 = fb_reg_redirect ? _GEN_274 : btb_pc_9; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_467 = fb_reg_redirect ? _GEN_275 : btb_pc_10; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_468 = fb_reg_redirect ? _GEN_276 : btb_pc_11; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_469 = fb_reg_redirect ? _GEN_277 : btb_pc_12; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_470 = fb_reg_redirect ? _GEN_278 : btb_pc_13; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_471 = fb_reg_redirect ? _GEN_279 : btb_pc_14; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_472 = fb_reg_redirect ? _GEN_280 : btb_pc_15; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_473 = fb_reg_redirect ? _GEN_281 : btb_pc_16; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_474 = fb_reg_redirect ? _GEN_282 : btb_pc_17; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_475 = fb_reg_redirect ? _GEN_283 : btb_pc_18; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_476 = fb_reg_redirect ? _GEN_284 : btb_pc_19; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_477 = fb_reg_redirect ? _GEN_285 : btb_pc_20; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_478 = fb_reg_redirect ? _GEN_286 : btb_pc_21; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_479 = fb_reg_redirect ? _GEN_287 : btb_pc_22; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_480 = fb_reg_redirect ? _GEN_288 : btb_pc_23; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_481 = fb_reg_redirect ? _GEN_289 : btb_pc_24; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_482 = fb_reg_redirect ? _GEN_290 : btb_pc_25; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_483 = fb_reg_redirect ? _GEN_291 : btb_pc_26; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_484 = fb_reg_redirect ? _GEN_292 : btb_pc_27; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_485 = fb_reg_redirect ? _GEN_293 : btb_pc_28; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_486 = fb_reg_redirect ? _GEN_294 : btb_pc_29; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_487 = fb_reg_redirect ? _GEN_295 : btb_pc_30; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_488 = fb_reg_redirect ? _GEN_296 : btb_pc_31; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_489 = fb_reg_redirect ? _GEN_297 : btb_pc_32; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_490 = fb_reg_redirect ? _GEN_298 : btb_pc_33; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_491 = fb_reg_redirect ? _GEN_299 : btb_pc_34; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_492 = fb_reg_redirect ? _GEN_300 : btb_pc_35; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_493 = fb_reg_redirect ? _GEN_301 : btb_pc_36; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_494 = fb_reg_redirect ? _GEN_302 : btb_pc_37; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_495 = fb_reg_redirect ? _GEN_303 : btb_pc_38; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_496 = fb_reg_redirect ? _GEN_304 : btb_pc_39; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_497 = fb_reg_redirect ? _GEN_305 : btb_pc_40; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_498 = fb_reg_redirect ? _GEN_306 : btb_pc_41; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_499 = fb_reg_redirect ? _GEN_307 : btb_pc_42; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_500 = fb_reg_redirect ? _GEN_308 : btb_pc_43; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_501 = fb_reg_redirect ? _GEN_309 : btb_pc_44; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_502 = fb_reg_redirect ? _GEN_310 : btb_pc_45; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_503 = fb_reg_redirect ? _GEN_311 : btb_pc_46; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_504 = fb_reg_redirect ? _GEN_312 : btb_pc_47; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_505 = fb_reg_redirect ? _GEN_313 : btb_pc_48; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_506 = fb_reg_redirect ? _GEN_314 : btb_pc_49; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_507 = fb_reg_redirect ? _GEN_315 : btb_pc_50; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_508 = fb_reg_redirect ? _GEN_316 : btb_pc_51; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_509 = fb_reg_redirect ? _GEN_317 : btb_pc_52; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_510 = fb_reg_redirect ? _GEN_318 : btb_pc_53; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_511 = fb_reg_redirect ? _GEN_319 : btb_pc_54; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_512 = fb_reg_redirect ? _GEN_320 : btb_pc_55; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_513 = fb_reg_redirect ? _GEN_321 : btb_pc_56; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_514 = fb_reg_redirect ? _GEN_322 : btb_pc_57; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_515 = fb_reg_redirect ? _GEN_323 : btb_pc_58; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_516 = fb_reg_redirect ? _GEN_324 : btb_pc_59; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_517 = fb_reg_redirect ? _GEN_325 : btb_pc_60; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_518 = fb_reg_redirect ? _GEN_326 : btb_pc_61; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_519 = fb_reg_redirect ? _GEN_327 : btb_pc_62; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_520 = fb_reg_redirect ? _GEN_328 : btb_pc_63; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_521 = fb_reg_redirect ? _GEN_329 : btb_tgt_0; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_522 = fb_reg_redirect ? _GEN_330 : btb_tgt_1; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_523 = fb_reg_redirect ? _GEN_331 : btb_tgt_2; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_524 = fb_reg_redirect ? _GEN_332 : btb_tgt_3; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_525 = fb_reg_redirect ? _GEN_333 : btb_tgt_4; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_526 = fb_reg_redirect ? _GEN_334 : btb_tgt_5; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_527 = fb_reg_redirect ? _GEN_335 : btb_tgt_6; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_528 = fb_reg_redirect ? _GEN_336 : btb_tgt_7; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_529 = fb_reg_redirect ? _GEN_337 : btb_tgt_8; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_530 = fb_reg_redirect ? _GEN_338 : btb_tgt_9; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_531 = fb_reg_redirect ? _GEN_339 : btb_tgt_10; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_532 = fb_reg_redirect ? _GEN_340 : btb_tgt_11; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_533 = fb_reg_redirect ? _GEN_341 : btb_tgt_12; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_534 = fb_reg_redirect ? _GEN_342 : btb_tgt_13; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_535 = fb_reg_redirect ? _GEN_343 : btb_tgt_14; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_536 = fb_reg_redirect ? _GEN_344 : btb_tgt_15; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_537 = fb_reg_redirect ? _GEN_345 : btb_tgt_16; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_538 = fb_reg_redirect ? _GEN_346 : btb_tgt_17; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_539 = fb_reg_redirect ? _GEN_347 : btb_tgt_18; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_540 = fb_reg_redirect ? _GEN_348 : btb_tgt_19; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_541 = fb_reg_redirect ? _GEN_349 : btb_tgt_20; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_542 = fb_reg_redirect ? _GEN_350 : btb_tgt_21; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_543 = fb_reg_redirect ? _GEN_351 : btb_tgt_22; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_544 = fb_reg_redirect ? _GEN_352 : btb_tgt_23; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_545 = fb_reg_redirect ? _GEN_353 : btb_tgt_24; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_546 = fb_reg_redirect ? _GEN_354 : btb_tgt_25; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_547 = fb_reg_redirect ? _GEN_355 : btb_tgt_26; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_548 = fb_reg_redirect ? _GEN_356 : btb_tgt_27; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_549 = fb_reg_redirect ? _GEN_357 : btb_tgt_28; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_550 = fb_reg_redirect ? _GEN_358 : btb_tgt_29; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_551 = fb_reg_redirect ? _GEN_359 : btb_tgt_30; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_552 = fb_reg_redirect ? _GEN_360 : btb_tgt_31; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_553 = fb_reg_redirect ? _GEN_361 : btb_tgt_32; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_554 = fb_reg_redirect ? _GEN_362 : btb_tgt_33; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_555 = fb_reg_redirect ? _GEN_363 : btb_tgt_34; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_556 = fb_reg_redirect ? _GEN_364 : btb_tgt_35; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_557 = fb_reg_redirect ? _GEN_365 : btb_tgt_36; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_558 = fb_reg_redirect ? _GEN_366 : btb_tgt_37; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_559 = fb_reg_redirect ? _GEN_367 : btb_tgt_38; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_560 = fb_reg_redirect ? _GEN_368 : btb_tgt_39; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_561 = fb_reg_redirect ? _GEN_369 : btb_tgt_40; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_562 = fb_reg_redirect ? _GEN_370 : btb_tgt_41; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_563 = fb_reg_redirect ? _GEN_371 : btb_tgt_42; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_564 = fb_reg_redirect ? _GEN_372 : btb_tgt_43; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_565 = fb_reg_redirect ? _GEN_373 : btb_tgt_44; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_566 = fb_reg_redirect ? _GEN_374 : btb_tgt_45; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_567 = fb_reg_redirect ? _GEN_375 : btb_tgt_46; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_568 = fb_reg_redirect ? _GEN_376 : btb_tgt_47; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_569 = fb_reg_redirect ? _GEN_377 : btb_tgt_48; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_570 = fb_reg_redirect ? _GEN_378 : btb_tgt_49; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_571 = fb_reg_redirect ? _GEN_379 : btb_tgt_50; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_572 = fb_reg_redirect ? _GEN_380 : btb_tgt_51; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_573 = fb_reg_redirect ? _GEN_381 : btb_tgt_52; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_574 = fb_reg_redirect ? _GEN_382 : btb_tgt_53; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_575 = fb_reg_redirect ? _GEN_383 : btb_tgt_54; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_576 = fb_reg_redirect ? _GEN_384 : btb_tgt_55; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_577 = fb_reg_redirect ? _GEN_385 : btb_tgt_56; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_578 = fb_reg_redirect ? _GEN_386 : btb_tgt_57; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_579 = fb_reg_redirect ? _GEN_387 : btb_tgt_58; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_580 = fb_reg_redirect ? _GEN_388 : btb_tgt_59; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_581 = fb_reg_redirect ? _GEN_389 : btb_tgt_60; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_582 = fb_reg_redirect ? _GEN_390 : btb_tgt_61; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_583 = fb_reg_redirect ? _GEN_391 : btb_tgt_62; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_584 = fb_reg_redirect ? _GEN_392 : btb_tgt_63; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_585 = fb_reg_redirect ? _GEN_393 : btb_bj_type_0; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_586 = fb_reg_redirect ? _GEN_394 : btb_bj_type_1; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_587 = fb_reg_redirect ? _GEN_395 : btb_bj_type_2; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_588 = fb_reg_redirect ? _GEN_396 : btb_bj_type_3; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_589 = fb_reg_redirect ? _GEN_397 : btb_bj_type_4; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_590 = fb_reg_redirect ? _GEN_398 : btb_bj_type_5; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_591 = fb_reg_redirect ? _GEN_399 : btb_bj_type_6; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_592 = fb_reg_redirect ? _GEN_400 : btb_bj_type_7; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_593 = fb_reg_redirect ? _GEN_401 : btb_bj_type_8; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_594 = fb_reg_redirect ? _GEN_402 : btb_bj_type_9; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_595 = fb_reg_redirect ? _GEN_403 : btb_bj_type_10; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_596 = fb_reg_redirect ? _GEN_404 : btb_bj_type_11; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_597 = fb_reg_redirect ? _GEN_405 : btb_bj_type_12; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_598 = fb_reg_redirect ? _GEN_406 : btb_bj_type_13; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_599 = fb_reg_redirect ? _GEN_407 : btb_bj_type_14; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_600 = fb_reg_redirect ? _GEN_408 : btb_bj_type_15; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_601 = fb_reg_redirect ? _GEN_409 : btb_bj_type_16; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_602 = fb_reg_redirect ? _GEN_410 : btb_bj_type_17; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_603 = fb_reg_redirect ? _GEN_411 : btb_bj_type_18; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_604 = fb_reg_redirect ? _GEN_412 : btb_bj_type_19; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_605 = fb_reg_redirect ? _GEN_413 : btb_bj_type_20; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_606 = fb_reg_redirect ? _GEN_414 : btb_bj_type_21; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_607 = fb_reg_redirect ? _GEN_415 : btb_bj_type_22; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_608 = fb_reg_redirect ? _GEN_416 : btb_bj_type_23; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_609 = fb_reg_redirect ? _GEN_417 : btb_bj_type_24; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_610 = fb_reg_redirect ? _GEN_418 : btb_bj_type_25; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_611 = fb_reg_redirect ? _GEN_419 : btb_bj_type_26; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_612 = fb_reg_redirect ? _GEN_420 : btb_bj_type_27; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_613 = fb_reg_redirect ? _GEN_421 : btb_bj_type_28; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_614 = fb_reg_redirect ? _GEN_422 : btb_bj_type_29; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_615 = fb_reg_redirect ? _GEN_423 : btb_bj_type_30; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_616 = fb_reg_redirect ? _GEN_424 : btb_bj_type_31; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_617 = fb_reg_redirect ? _GEN_425 : btb_bj_type_32; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_618 = fb_reg_redirect ? _GEN_426 : btb_bj_type_33; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_619 = fb_reg_redirect ? _GEN_427 : btb_bj_type_34; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_620 = fb_reg_redirect ? _GEN_428 : btb_bj_type_35; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_621 = fb_reg_redirect ? _GEN_429 : btb_bj_type_36; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_622 = fb_reg_redirect ? _GEN_430 : btb_bj_type_37; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_623 = fb_reg_redirect ? _GEN_431 : btb_bj_type_38; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_624 = fb_reg_redirect ? _GEN_432 : btb_bj_type_39; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_625 = fb_reg_redirect ? _GEN_433 : btb_bj_type_40; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_626 = fb_reg_redirect ? _GEN_434 : btb_bj_type_41; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_627 = fb_reg_redirect ? _GEN_435 : btb_bj_type_42; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_628 = fb_reg_redirect ? _GEN_436 : btb_bj_type_43; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_629 = fb_reg_redirect ? _GEN_437 : btb_bj_type_44; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_630 = fb_reg_redirect ? _GEN_438 : btb_bj_type_45; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_631 = fb_reg_redirect ? _GEN_439 : btb_bj_type_46; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_632 = fb_reg_redirect ? _GEN_440 : btb_bj_type_47; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_633 = fb_reg_redirect ? _GEN_441 : btb_bj_type_48; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_634 = fb_reg_redirect ? _GEN_442 : btb_bj_type_49; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_635 = fb_reg_redirect ? _GEN_443 : btb_bj_type_50; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_636 = fb_reg_redirect ? _GEN_444 : btb_bj_type_51; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_637 = fb_reg_redirect ? _GEN_445 : btb_bj_type_52; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_638 = fb_reg_redirect ? _GEN_446 : btb_bj_type_53; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_639 = fb_reg_redirect ? _GEN_447 : btb_bj_type_54; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_640 = fb_reg_redirect ? _GEN_448 : btb_bj_type_55; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_641 = fb_reg_redirect ? _GEN_449 : btb_bj_type_56; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_642 = fb_reg_redirect ? _GEN_450 : btb_bj_type_57; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_643 = fb_reg_redirect ? _GEN_451 : btb_bj_type_58; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_644 = fb_reg_redirect ? _GEN_452 : btb_bj_type_59; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_645 = fb_reg_redirect ? _GEN_453 : btb_bj_type_60; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_646 = fb_reg_redirect ? _GEN_454 : btb_bj_type_61; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_647 = fb_reg_redirect ? _GEN_455 : btb_bj_type_62; // @[BTB.scala 205:28:@3705.6]
  assign _GEN_648 = fb_reg_redirect ? _GEN_456 : btb_bj_type_63; // @[BTB.scala 205:28:@3705.6]
  assign _T_3291 = feedback_h_count != 2'h0; // @[BTB.scala 72:38:@3715.12]
  assign _T_3292 = feedback_h_count[1]; // @[BTB.scala 72:45:@3716.12]
  assign _T_3293 = feedback_h_count[0]; // @[BTB.scala 72:54:@3717.12]
  assign _T_3295 = _T_3293 == 1'h0; // @[BTB.scala 72:52:@3718.12]
  assign _T_3296 = _T_3292 | _T_3295; // @[BTB.scala 72:49:@3719.12]
  assign _T_3297 = {_T_3291,_T_3296}; // @[Cat.scala 30:58:@3720.12]
  assign _GEN_649 = 6'h0 == feedback_idx ? _T_3297 : btb_h_count_0; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_650 = 6'h1 == feedback_idx ? _T_3297 : btb_h_count_1; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_651 = 6'h2 == feedback_idx ? _T_3297 : btb_h_count_2; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_652 = 6'h3 == feedback_idx ? _T_3297 : btb_h_count_3; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_653 = 6'h4 == feedback_idx ? _T_3297 : btb_h_count_4; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_654 = 6'h5 == feedback_idx ? _T_3297 : btb_h_count_5; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_655 = 6'h6 == feedback_idx ? _T_3297 : btb_h_count_6; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_656 = 6'h7 == feedback_idx ? _T_3297 : btb_h_count_7; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_657 = 6'h8 == feedback_idx ? _T_3297 : btb_h_count_8; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_658 = 6'h9 == feedback_idx ? _T_3297 : btb_h_count_9; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_659 = 6'ha == feedback_idx ? _T_3297 : btb_h_count_10; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_660 = 6'hb == feedback_idx ? _T_3297 : btb_h_count_11; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_661 = 6'hc == feedback_idx ? _T_3297 : btb_h_count_12; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_662 = 6'hd == feedback_idx ? _T_3297 : btb_h_count_13; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_663 = 6'he == feedback_idx ? _T_3297 : btb_h_count_14; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_664 = 6'hf == feedback_idx ? _T_3297 : btb_h_count_15; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_665 = 6'h10 == feedback_idx ? _T_3297 : btb_h_count_16; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_666 = 6'h11 == feedback_idx ? _T_3297 : btb_h_count_17; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_667 = 6'h12 == feedback_idx ? _T_3297 : btb_h_count_18; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_668 = 6'h13 == feedback_idx ? _T_3297 : btb_h_count_19; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_669 = 6'h14 == feedback_idx ? _T_3297 : btb_h_count_20; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_670 = 6'h15 == feedback_idx ? _T_3297 : btb_h_count_21; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_671 = 6'h16 == feedback_idx ? _T_3297 : btb_h_count_22; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_672 = 6'h17 == feedback_idx ? _T_3297 : btb_h_count_23; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_673 = 6'h18 == feedback_idx ? _T_3297 : btb_h_count_24; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_674 = 6'h19 == feedback_idx ? _T_3297 : btb_h_count_25; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_675 = 6'h1a == feedback_idx ? _T_3297 : btb_h_count_26; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_676 = 6'h1b == feedback_idx ? _T_3297 : btb_h_count_27; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_677 = 6'h1c == feedback_idx ? _T_3297 : btb_h_count_28; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_678 = 6'h1d == feedback_idx ? _T_3297 : btb_h_count_29; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_679 = 6'h1e == feedback_idx ? _T_3297 : btb_h_count_30; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_680 = 6'h1f == feedback_idx ? _T_3297 : btb_h_count_31; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_681 = 6'h20 == feedback_idx ? _T_3297 : btb_h_count_32; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_682 = 6'h21 == feedback_idx ? _T_3297 : btb_h_count_33; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_683 = 6'h22 == feedback_idx ? _T_3297 : btb_h_count_34; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_684 = 6'h23 == feedback_idx ? _T_3297 : btb_h_count_35; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_685 = 6'h24 == feedback_idx ? _T_3297 : btb_h_count_36; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_686 = 6'h25 == feedback_idx ? _T_3297 : btb_h_count_37; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_687 = 6'h26 == feedback_idx ? _T_3297 : btb_h_count_38; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_688 = 6'h27 == feedback_idx ? _T_3297 : btb_h_count_39; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_689 = 6'h28 == feedback_idx ? _T_3297 : btb_h_count_40; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_690 = 6'h29 == feedback_idx ? _T_3297 : btb_h_count_41; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_691 = 6'h2a == feedback_idx ? _T_3297 : btb_h_count_42; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_692 = 6'h2b == feedback_idx ? _T_3297 : btb_h_count_43; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_693 = 6'h2c == feedback_idx ? _T_3297 : btb_h_count_44; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_694 = 6'h2d == feedback_idx ? _T_3297 : btb_h_count_45; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_695 = 6'h2e == feedback_idx ? _T_3297 : btb_h_count_46; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_696 = 6'h2f == feedback_idx ? _T_3297 : btb_h_count_47; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_697 = 6'h30 == feedback_idx ? _T_3297 : btb_h_count_48; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_698 = 6'h31 == feedback_idx ? _T_3297 : btb_h_count_49; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_699 = 6'h32 == feedback_idx ? _T_3297 : btb_h_count_50; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_700 = 6'h33 == feedback_idx ? _T_3297 : btb_h_count_51; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_701 = 6'h34 == feedback_idx ? _T_3297 : btb_h_count_52; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_702 = 6'h35 == feedback_idx ? _T_3297 : btb_h_count_53; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_703 = 6'h36 == feedback_idx ? _T_3297 : btb_h_count_54; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_704 = 6'h37 == feedback_idx ? _T_3297 : btb_h_count_55; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_705 = 6'h38 == feedback_idx ? _T_3297 : btb_h_count_56; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_706 = 6'h39 == feedback_idx ? _T_3297 : btb_h_count_57; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_707 = 6'h3a == feedback_idx ? _T_3297 : btb_h_count_58; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_708 = 6'h3b == feedback_idx ? _T_3297 : btb_h_count_59; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_709 = 6'h3c == feedback_idx ? _T_3297 : btb_h_count_60; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_710 = 6'h3d == feedback_idx ? _T_3297 : btb_h_count_61; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_711 = 6'h3e == feedback_idx ? _T_3297 : btb_h_count_62; // @[BTB.scala 214:37:@3721.12]
  assign _GEN_712 = 6'h3f == feedback_idx ? _T_3297 : btb_h_count_63; // @[BTB.scala 214:37:@3721.12]
  assign feedback_gshare = bht__T_2923_data; // @[BTB.scala 184:22:@2953.4 BTB.scala 194:20:@3406.4]
  assign _T_3300 = feedback_gshare != 2'h0; // @[BTB.scala 72:38:@3723.12]
  assign _T_3301 = feedback_gshare[1]; // @[BTB.scala 72:45:@3724.12]
  assign _T_3302 = feedback_gshare[0]; // @[BTB.scala 72:54:@3725.12]
  assign _T_3304 = _T_3302 == 1'h0; // @[BTB.scala 72:52:@3726.12]
  assign _T_3305 = _T_3301 | _T_3304; // @[BTB.scala 72:49:@3727.12]
  assign _T_3307 = ~ feedback_h_count; // @[BTB.scala 74:38:@3732.12]
  assign _T_3309 = _T_3307 == 2'h0; // @[BTB.scala 74:38:@3733.12]
  assign _T_3314 = _T_3292 & _T_3295; // @[BTB.scala 74:49:@3737.12]
  assign _T_3315 = {_T_3309,_T_3314}; // @[Cat.scala 30:58:@3738.12]
  assign _GEN_713 = 6'h0 == feedback_idx ? _T_3315 : btb_h_count_0; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_714 = 6'h1 == feedback_idx ? _T_3315 : btb_h_count_1; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_715 = 6'h2 == feedback_idx ? _T_3315 : btb_h_count_2; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_716 = 6'h3 == feedback_idx ? _T_3315 : btb_h_count_3; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_717 = 6'h4 == feedback_idx ? _T_3315 : btb_h_count_4; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_718 = 6'h5 == feedback_idx ? _T_3315 : btb_h_count_5; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_719 = 6'h6 == feedback_idx ? _T_3315 : btb_h_count_6; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_720 = 6'h7 == feedback_idx ? _T_3315 : btb_h_count_7; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_721 = 6'h8 == feedback_idx ? _T_3315 : btb_h_count_8; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_722 = 6'h9 == feedback_idx ? _T_3315 : btb_h_count_9; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_723 = 6'ha == feedback_idx ? _T_3315 : btb_h_count_10; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_724 = 6'hb == feedback_idx ? _T_3315 : btb_h_count_11; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_725 = 6'hc == feedback_idx ? _T_3315 : btb_h_count_12; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_726 = 6'hd == feedback_idx ? _T_3315 : btb_h_count_13; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_727 = 6'he == feedback_idx ? _T_3315 : btb_h_count_14; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_728 = 6'hf == feedback_idx ? _T_3315 : btb_h_count_15; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_729 = 6'h10 == feedback_idx ? _T_3315 : btb_h_count_16; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_730 = 6'h11 == feedback_idx ? _T_3315 : btb_h_count_17; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_731 = 6'h12 == feedback_idx ? _T_3315 : btb_h_count_18; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_732 = 6'h13 == feedback_idx ? _T_3315 : btb_h_count_19; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_733 = 6'h14 == feedback_idx ? _T_3315 : btb_h_count_20; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_734 = 6'h15 == feedback_idx ? _T_3315 : btb_h_count_21; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_735 = 6'h16 == feedback_idx ? _T_3315 : btb_h_count_22; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_736 = 6'h17 == feedback_idx ? _T_3315 : btb_h_count_23; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_737 = 6'h18 == feedback_idx ? _T_3315 : btb_h_count_24; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_738 = 6'h19 == feedback_idx ? _T_3315 : btb_h_count_25; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_739 = 6'h1a == feedback_idx ? _T_3315 : btb_h_count_26; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_740 = 6'h1b == feedback_idx ? _T_3315 : btb_h_count_27; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_741 = 6'h1c == feedback_idx ? _T_3315 : btb_h_count_28; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_742 = 6'h1d == feedback_idx ? _T_3315 : btb_h_count_29; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_743 = 6'h1e == feedback_idx ? _T_3315 : btb_h_count_30; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_744 = 6'h1f == feedback_idx ? _T_3315 : btb_h_count_31; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_745 = 6'h20 == feedback_idx ? _T_3315 : btb_h_count_32; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_746 = 6'h21 == feedback_idx ? _T_3315 : btb_h_count_33; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_747 = 6'h22 == feedback_idx ? _T_3315 : btb_h_count_34; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_748 = 6'h23 == feedback_idx ? _T_3315 : btb_h_count_35; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_749 = 6'h24 == feedback_idx ? _T_3315 : btb_h_count_36; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_750 = 6'h25 == feedback_idx ? _T_3315 : btb_h_count_37; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_751 = 6'h26 == feedback_idx ? _T_3315 : btb_h_count_38; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_752 = 6'h27 == feedback_idx ? _T_3315 : btb_h_count_39; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_753 = 6'h28 == feedback_idx ? _T_3315 : btb_h_count_40; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_754 = 6'h29 == feedback_idx ? _T_3315 : btb_h_count_41; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_755 = 6'h2a == feedback_idx ? _T_3315 : btb_h_count_42; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_756 = 6'h2b == feedback_idx ? _T_3315 : btb_h_count_43; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_757 = 6'h2c == feedback_idx ? _T_3315 : btb_h_count_44; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_758 = 6'h2d == feedback_idx ? _T_3315 : btb_h_count_45; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_759 = 6'h2e == feedback_idx ? _T_3315 : btb_h_count_46; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_760 = 6'h2f == feedback_idx ? _T_3315 : btb_h_count_47; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_761 = 6'h30 == feedback_idx ? _T_3315 : btb_h_count_48; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_762 = 6'h31 == feedback_idx ? _T_3315 : btb_h_count_49; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_763 = 6'h32 == feedback_idx ? _T_3315 : btb_h_count_50; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_764 = 6'h33 == feedback_idx ? _T_3315 : btb_h_count_51; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_765 = 6'h34 == feedback_idx ? _T_3315 : btb_h_count_52; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_766 = 6'h35 == feedback_idx ? _T_3315 : btb_h_count_53; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_767 = 6'h36 == feedback_idx ? _T_3315 : btb_h_count_54; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_768 = 6'h37 == feedback_idx ? _T_3315 : btb_h_count_55; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_769 = 6'h38 == feedback_idx ? _T_3315 : btb_h_count_56; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_770 = 6'h39 == feedback_idx ? _T_3315 : btb_h_count_57; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_771 = 6'h3a == feedback_idx ? _T_3315 : btb_h_count_58; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_772 = 6'h3b == feedback_idx ? _T_3315 : btb_h_count_59; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_773 = 6'h3c == feedback_idx ? _T_3315 : btb_h_count_60; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_774 = 6'h3d == feedback_idx ? _T_3315 : btb_h_count_61; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_775 = 6'h3e == feedback_idx ? _T_3315 : btb_h_count_62; // @[BTB.scala 217:37:@3739.12]
  assign _GEN_776 = 6'h3f == feedback_idx ? _T_3315 : btb_h_count_63; // @[BTB.scala 217:37:@3739.12]
  assign _T_3317 = ~ feedback_gshare; // @[BTB.scala 74:38:@3741.12]
  assign _T_3319 = _T_3317 == 2'h0; // @[BTB.scala 74:38:@3742.12]
  assign _T_3324 = _T_3301 & _T_3304; // @[BTB.scala 74:49:@3746.12]
  assign _GEN_777 = fb_reg_redirect ? _GEN_649 : _GEN_713; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_778 = fb_reg_redirect ? _GEN_650 : _GEN_714; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_779 = fb_reg_redirect ? _GEN_651 : _GEN_715; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_780 = fb_reg_redirect ? _GEN_652 : _GEN_716; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_781 = fb_reg_redirect ? _GEN_653 : _GEN_717; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_782 = fb_reg_redirect ? _GEN_654 : _GEN_718; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_783 = fb_reg_redirect ? _GEN_655 : _GEN_719; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_784 = fb_reg_redirect ? _GEN_656 : _GEN_720; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_785 = fb_reg_redirect ? _GEN_657 : _GEN_721; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_786 = fb_reg_redirect ? _GEN_658 : _GEN_722; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_787 = fb_reg_redirect ? _GEN_659 : _GEN_723; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_788 = fb_reg_redirect ? _GEN_660 : _GEN_724; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_789 = fb_reg_redirect ? _GEN_661 : _GEN_725; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_790 = fb_reg_redirect ? _GEN_662 : _GEN_726; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_791 = fb_reg_redirect ? _GEN_663 : _GEN_727; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_792 = fb_reg_redirect ? _GEN_664 : _GEN_728; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_793 = fb_reg_redirect ? _GEN_665 : _GEN_729; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_794 = fb_reg_redirect ? _GEN_666 : _GEN_730; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_795 = fb_reg_redirect ? _GEN_667 : _GEN_731; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_796 = fb_reg_redirect ? _GEN_668 : _GEN_732; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_797 = fb_reg_redirect ? _GEN_669 : _GEN_733; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_798 = fb_reg_redirect ? _GEN_670 : _GEN_734; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_799 = fb_reg_redirect ? _GEN_671 : _GEN_735; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_800 = fb_reg_redirect ? _GEN_672 : _GEN_736; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_801 = fb_reg_redirect ? _GEN_673 : _GEN_737; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_802 = fb_reg_redirect ? _GEN_674 : _GEN_738; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_803 = fb_reg_redirect ? _GEN_675 : _GEN_739; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_804 = fb_reg_redirect ? _GEN_676 : _GEN_740; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_805 = fb_reg_redirect ? _GEN_677 : _GEN_741; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_806 = fb_reg_redirect ? _GEN_678 : _GEN_742; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_807 = fb_reg_redirect ? _GEN_679 : _GEN_743; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_808 = fb_reg_redirect ? _GEN_680 : _GEN_744; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_809 = fb_reg_redirect ? _GEN_681 : _GEN_745; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_810 = fb_reg_redirect ? _GEN_682 : _GEN_746; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_811 = fb_reg_redirect ? _GEN_683 : _GEN_747; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_812 = fb_reg_redirect ? _GEN_684 : _GEN_748; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_813 = fb_reg_redirect ? _GEN_685 : _GEN_749; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_814 = fb_reg_redirect ? _GEN_686 : _GEN_750; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_815 = fb_reg_redirect ? _GEN_687 : _GEN_751; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_816 = fb_reg_redirect ? _GEN_688 : _GEN_752; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_817 = fb_reg_redirect ? _GEN_689 : _GEN_753; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_818 = fb_reg_redirect ? _GEN_690 : _GEN_754; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_819 = fb_reg_redirect ? _GEN_691 : _GEN_755; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_820 = fb_reg_redirect ? _GEN_692 : _GEN_756; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_821 = fb_reg_redirect ? _GEN_693 : _GEN_757; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_822 = fb_reg_redirect ? _GEN_694 : _GEN_758; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_823 = fb_reg_redirect ? _GEN_695 : _GEN_759; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_824 = fb_reg_redirect ? _GEN_696 : _GEN_760; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_825 = fb_reg_redirect ? _GEN_697 : _GEN_761; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_826 = fb_reg_redirect ? _GEN_698 : _GEN_762; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_827 = fb_reg_redirect ? _GEN_699 : _GEN_763; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_828 = fb_reg_redirect ? _GEN_700 : _GEN_764; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_829 = fb_reg_redirect ? _GEN_701 : _GEN_765; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_830 = fb_reg_redirect ? _GEN_702 : _GEN_766; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_831 = fb_reg_redirect ? _GEN_703 : _GEN_767; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_832 = fb_reg_redirect ? _GEN_704 : _GEN_768; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_833 = fb_reg_redirect ? _GEN_705 : _GEN_769; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_834 = fb_reg_redirect ? _GEN_706 : _GEN_770; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_835 = fb_reg_redirect ? _GEN_707 : _GEN_771; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_836 = fb_reg_redirect ? _GEN_708 : _GEN_772; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_837 = fb_reg_redirect ? _GEN_709 : _GEN_773; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_838 = fb_reg_redirect ? _GEN_710 : _GEN_774; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_839 = fb_reg_redirect ? _GEN_711 : _GEN_775; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_840 = fb_reg_redirect ? _GEN_712 : _GEN_776; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_848 = fb_reg_redirect ? 1'h0 : 1'h1; // @[BTB.scala 213:32:@3714.10]
  assign _GEN_851 = 6'h0 == feedback_idx ? 2'h2 : btb_h_count_0; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_852 = 6'h1 == feedback_idx ? 2'h2 : btb_h_count_1; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_853 = 6'h2 == feedback_idx ? 2'h2 : btb_h_count_2; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_854 = 6'h3 == feedback_idx ? 2'h2 : btb_h_count_3; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_855 = 6'h4 == feedback_idx ? 2'h2 : btb_h_count_4; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_856 = 6'h5 == feedback_idx ? 2'h2 : btb_h_count_5; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_857 = 6'h6 == feedback_idx ? 2'h2 : btb_h_count_6; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_858 = 6'h7 == feedback_idx ? 2'h2 : btb_h_count_7; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_859 = 6'h8 == feedback_idx ? 2'h2 : btb_h_count_8; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_860 = 6'h9 == feedback_idx ? 2'h2 : btb_h_count_9; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_861 = 6'ha == feedback_idx ? 2'h2 : btb_h_count_10; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_862 = 6'hb == feedback_idx ? 2'h2 : btb_h_count_11; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_863 = 6'hc == feedback_idx ? 2'h2 : btb_h_count_12; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_864 = 6'hd == feedback_idx ? 2'h2 : btb_h_count_13; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_865 = 6'he == feedback_idx ? 2'h2 : btb_h_count_14; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_866 = 6'hf == feedback_idx ? 2'h2 : btb_h_count_15; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_867 = 6'h10 == feedback_idx ? 2'h2 : btb_h_count_16; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_868 = 6'h11 == feedback_idx ? 2'h2 : btb_h_count_17; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_869 = 6'h12 == feedback_idx ? 2'h2 : btb_h_count_18; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_870 = 6'h13 == feedback_idx ? 2'h2 : btb_h_count_19; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_871 = 6'h14 == feedback_idx ? 2'h2 : btb_h_count_20; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_872 = 6'h15 == feedback_idx ? 2'h2 : btb_h_count_21; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_873 = 6'h16 == feedback_idx ? 2'h2 : btb_h_count_22; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_874 = 6'h17 == feedback_idx ? 2'h2 : btb_h_count_23; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_875 = 6'h18 == feedback_idx ? 2'h2 : btb_h_count_24; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_876 = 6'h19 == feedback_idx ? 2'h2 : btb_h_count_25; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_877 = 6'h1a == feedback_idx ? 2'h2 : btb_h_count_26; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_878 = 6'h1b == feedback_idx ? 2'h2 : btb_h_count_27; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_879 = 6'h1c == feedback_idx ? 2'h2 : btb_h_count_28; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_880 = 6'h1d == feedback_idx ? 2'h2 : btb_h_count_29; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_881 = 6'h1e == feedback_idx ? 2'h2 : btb_h_count_30; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_882 = 6'h1f == feedback_idx ? 2'h2 : btb_h_count_31; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_883 = 6'h20 == feedback_idx ? 2'h2 : btb_h_count_32; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_884 = 6'h21 == feedback_idx ? 2'h2 : btb_h_count_33; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_885 = 6'h22 == feedback_idx ? 2'h2 : btb_h_count_34; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_886 = 6'h23 == feedback_idx ? 2'h2 : btb_h_count_35; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_887 = 6'h24 == feedback_idx ? 2'h2 : btb_h_count_36; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_888 = 6'h25 == feedback_idx ? 2'h2 : btb_h_count_37; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_889 = 6'h26 == feedback_idx ? 2'h2 : btb_h_count_38; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_890 = 6'h27 == feedback_idx ? 2'h2 : btb_h_count_39; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_891 = 6'h28 == feedback_idx ? 2'h2 : btb_h_count_40; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_892 = 6'h29 == feedback_idx ? 2'h2 : btb_h_count_41; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_893 = 6'h2a == feedback_idx ? 2'h2 : btb_h_count_42; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_894 = 6'h2b == feedback_idx ? 2'h2 : btb_h_count_43; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_895 = 6'h2c == feedback_idx ? 2'h2 : btb_h_count_44; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_896 = 6'h2d == feedback_idx ? 2'h2 : btb_h_count_45; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_897 = 6'h2e == feedback_idx ? 2'h2 : btb_h_count_46; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_898 = 6'h2f == feedback_idx ? 2'h2 : btb_h_count_47; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_899 = 6'h30 == feedback_idx ? 2'h2 : btb_h_count_48; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_900 = 6'h31 == feedback_idx ? 2'h2 : btb_h_count_49; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_901 = 6'h32 == feedback_idx ? 2'h2 : btb_h_count_50; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_902 = 6'h33 == feedback_idx ? 2'h2 : btb_h_count_51; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_903 = 6'h34 == feedback_idx ? 2'h2 : btb_h_count_52; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_904 = 6'h35 == feedback_idx ? 2'h2 : btb_h_count_53; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_905 = 6'h36 == feedback_idx ? 2'h2 : btb_h_count_54; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_906 = 6'h37 == feedback_idx ? 2'h2 : btb_h_count_55; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_907 = 6'h38 == feedback_idx ? 2'h2 : btb_h_count_56; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_908 = 6'h39 == feedback_idx ? 2'h2 : btb_h_count_57; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_909 = 6'h3a == feedback_idx ? 2'h2 : btb_h_count_58; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_910 = 6'h3b == feedback_idx ? 2'h2 : btb_h_count_59; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_911 = 6'h3c == feedback_idx ? 2'h2 : btb_h_count_60; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_912 = 6'h3d == feedback_idx ? 2'h2 : btb_h_count_61; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_913 = 6'h3e == feedback_idx ? 2'h2 : btb_h_count_62; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_914 = 6'h3f == feedback_idx ? 2'h2 : btb_h_count_63; // @[BTB.scala 221:35:@3753.12]
  assign _GEN_915 = fb_reg_redirect ? _GEN_851 : btb_h_count_0; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_916 = fb_reg_redirect ? _GEN_852 : btb_h_count_1; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_917 = fb_reg_redirect ? _GEN_853 : btb_h_count_2; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_918 = fb_reg_redirect ? _GEN_854 : btb_h_count_3; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_919 = fb_reg_redirect ? _GEN_855 : btb_h_count_4; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_920 = fb_reg_redirect ? _GEN_856 : btb_h_count_5; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_921 = fb_reg_redirect ? _GEN_857 : btb_h_count_6; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_922 = fb_reg_redirect ? _GEN_858 : btb_h_count_7; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_923 = fb_reg_redirect ? _GEN_859 : btb_h_count_8; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_924 = fb_reg_redirect ? _GEN_860 : btb_h_count_9; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_925 = fb_reg_redirect ? _GEN_861 : btb_h_count_10; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_926 = fb_reg_redirect ? _GEN_862 : btb_h_count_11; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_927 = fb_reg_redirect ? _GEN_863 : btb_h_count_12; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_928 = fb_reg_redirect ? _GEN_864 : btb_h_count_13; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_929 = fb_reg_redirect ? _GEN_865 : btb_h_count_14; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_930 = fb_reg_redirect ? _GEN_866 : btb_h_count_15; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_931 = fb_reg_redirect ? _GEN_867 : btb_h_count_16; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_932 = fb_reg_redirect ? _GEN_868 : btb_h_count_17; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_933 = fb_reg_redirect ? _GEN_869 : btb_h_count_18; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_934 = fb_reg_redirect ? _GEN_870 : btb_h_count_19; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_935 = fb_reg_redirect ? _GEN_871 : btb_h_count_20; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_936 = fb_reg_redirect ? _GEN_872 : btb_h_count_21; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_937 = fb_reg_redirect ? _GEN_873 : btb_h_count_22; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_938 = fb_reg_redirect ? _GEN_874 : btb_h_count_23; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_939 = fb_reg_redirect ? _GEN_875 : btb_h_count_24; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_940 = fb_reg_redirect ? _GEN_876 : btb_h_count_25; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_941 = fb_reg_redirect ? _GEN_877 : btb_h_count_26; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_942 = fb_reg_redirect ? _GEN_878 : btb_h_count_27; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_943 = fb_reg_redirect ? _GEN_879 : btb_h_count_28; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_944 = fb_reg_redirect ? _GEN_880 : btb_h_count_29; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_945 = fb_reg_redirect ? _GEN_881 : btb_h_count_30; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_946 = fb_reg_redirect ? _GEN_882 : btb_h_count_31; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_947 = fb_reg_redirect ? _GEN_883 : btb_h_count_32; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_948 = fb_reg_redirect ? _GEN_884 : btb_h_count_33; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_949 = fb_reg_redirect ? _GEN_885 : btb_h_count_34; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_950 = fb_reg_redirect ? _GEN_886 : btb_h_count_35; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_951 = fb_reg_redirect ? _GEN_887 : btb_h_count_36; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_952 = fb_reg_redirect ? _GEN_888 : btb_h_count_37; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_953 = fb_reg_redirect ? _GEN_889 : btb_h_count_38; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_954 = fb_reg_redirect ? _GEN_890 : btb_h_count_39; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_955 = fb_reg_redirect ? _GEN_891 : btb_h_count_40; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_956 = fb_reg_redirect ? _GEN_892 : btb_h_count_41; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_957 = fb_reg_redirect ? _GEN_893 : btb_h_count_42; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_958 = fb_reg_redirect ? _GEN_894 : btb_h_count_43; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_959 = fb_reg_redirect ? _GEN_895 : btb_h_count_44; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_960 = fb_reg_redirect ? _GEN_896 : btb_h_count_45; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_961 = fb_reg_redirect ? _GEN_897 : btb_h_count_46; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_962 = fb_reg_redirect ? _GEN_898 : btb_h_count_47; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_963 = fb_reg_redirect ? _GEN_899 : btb_h_count_48; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_964 = fb_reg_redirect ? _GEN_900 : btb_h_count_49; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_965 = fb_reg_redirect ? _GEN_901 : btb_h_count_50; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_966 = fb_reg_redirect ? _GEN_902 : btb_h_count_51; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_967 = fb_reg_redirect ? _GEN_903 : btb_h_count_52; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_968 = fb_reg_redirect ? _GEN_904 : btb_h_count_53; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_969 = fb_reg_redirect ? _GEN_905 : btb_h_count_54; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_970 = fb_reg_redirect ? _GEN_906 : btb_h_count_55; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_971 = fb_reg_redirect ? _GEN_907 : btb_h_count_56; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_972 = fb_reg_redirect ? _GEN_908 : btb_h_count_57; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_973 = fb_reg_redirect ? _GEN_909 : btb_h_count_58; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_974 = fb_reg_redirect ? _GEN_910 : btb_h_count_59; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_975 = fb_reg_redirect ? _GEN_911 : btb_h_count_60; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_976 = fb_reg_redirect ? _GEN_912 : btb_h_count_61; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_977 = fb_reg_redirect ? _GEN_913 : btb_h_count_62; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_978 = fb_reg_redirect ? _GEN_914 : btb_h_count_63; // @[BTB.scala 220:35:@3752.10]
  assign _GEN_980 = _T_2925 ? _GEN_777 : _GEN_915; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_981 = _T_2925 ? _GEN_778 : _GEN_916; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_982 = _T_2925 ? _GEN_779 : _GEN_917; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_983 = _T_2925 ? _GEN_780 : _GEN_918; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_984 = _T_2925 ? _GEN_781 : _GEN_919; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_985 = _T_2925 ? _GEN_782 : _GEN_920; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_986 = _T_2925 ? _GEN_783 : _GEN_921; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_987 = _T_2925 ? _GEN_784 : _GEN_922; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_988 = _T_2925 ? _GEN_785 : _GEN_923; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_989 = _T_2925 ? _GEN_786 : _GEN_924; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_990 = _T_2925 ? _GEN_787 : _GEN_925; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_991 = _T_2925 ? _GEN_788 : _GEN_926; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_992 = _T_2925 ? _GEN_789 : _GEN_927; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_993 = _T_2925 ? _GEN_790 : _GEN_928; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_994 = _T_2925 ? _GEN_791 : _GEN_929; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_995 = _T_2925 ? _GEN_792 : _GEN_930; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_996 = _T_2925 ? _GEN_793 : _GEN_931; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_997 = _T_2925 ? _GEN_794 : _GEN_932; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_998 = _T_2925 ? _GEN_795 : _GEN_933; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_999 = _T_2925 ? _GEN_796 : _GEN_934; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1000 = _T_2925 ? _GEN_797 : _GEN_935; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1001 = _T_2925 ? _GEN_798 : _GEN_936; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1002 = _T_2925 ? _GEN_799 : _GEN_937; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1003 = _T_2925 ? _GEN_800 : _GEN_938; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1004 = _T_2925 ? _GEN_801 : _GEN_939; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1005 = _T_2925 ? _GEN_802 : _GEN_940; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1006 = _T_2925 ? _GEN_803 : _GEN_941; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1007 = _T_2925 ? _GEN_804 : _GEN_942; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1008 = _T_2925 ? _GEN_805 : _GEN_943; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1009 = _T_2925 ? _GEN_806 : _GEN_944; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1010 = _T_2925 ? _GEN_807 : _GEN_945; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1011 = _T_2925 ? _GEN_808 : _GEN_946; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1012 = _T_2925 ? _GEN_809 : _GEN_947; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1013 = _T_2925 ? _GEN_810 : _GEN_948; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1014 = _T_2925 ? _GEN_811 : _GEN_949; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1015 = _T_2925 ? _GEN_812 : _GEN_950; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1016 = _T_2925 ? _GEN_813 : _GEN_951; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1017 = _T_2925 ? _GEN_814 : _GEN_952; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1018 = _T_2925 ? _GEN_815 : _GEN_953; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1019 = _T_2925 ? _GEN_816 : _GEN_954; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1020 = _T_2925 ? _GEN_817 : _GEN_955; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1021 = _T_2925 ? _GEN_818 : _GEN_956; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1022 = _T_2925 ? _GEN_819 : _GEN_957; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1023 = _T_2925 ? _GEN_820 : _GEN_958; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1024 = _T_2925 ? _GEN_821 : _GEN_959; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1025 = _T_2925 ? _GEN_822 : _GEN_960; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1026 = _T_2925 ? _GEN_823 : _GEN_961; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1027 = _T_2925 ? _GEN_824 : _GEN_962; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1028 = _T_2925 ? _GEN_825 : _GEN_963; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1029 = _T_2925 ? _GEN_826 : _GEN_964; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1030 = _T_2925 ? _GEN_827 : _GEN_965; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1031 = _T_2925 ? _GEN_828 : _GEN_966; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1032 = _T_2925 ? _GEN_829 : _GEN_967; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1033 = _T_2925 ? _GEN_830 : _GEN_968; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1034 = _T_2925 ? _GEN_831 : _GEN_969; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1035 = _T_2925 ? _GEN_832 : _GEN_970; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1036 = _T_2925 ? _GEN_833 : _GEN_971; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1037 = _T_2925 ? _GEN_834 : _GEN_972; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1038 = _T_2925 ? _GEN_835 : _GEN_973; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1039 = _T_2925 ? _GEN_836 : _GEN_974; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1040 = _T_2925 ? _GEN_837 : _GEN_975; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1041 = _T_2925 ? _GEN_838 : _GEN_976; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1042 = _T_2925 ? _GEN_839 : _GEN_977; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1043 = _T_2925 ? _GEN_840 : _GEN_978; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1046 = _T_2925 ? fb_reg_redirect : 1'h0; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1051 = _T_2925 ? _GEN_848 : 1'h0; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1056 = _T_2925 ? 1'h0 : fb_reg_redirect; // @[BTB.scala 212:29:@3713.8]
  assign _GEN_1059 = _T_3285 ? _GEN_980 : btb_h_count_0; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1060 = _T_3285 ? _GEN_981 : btb_h_count_1; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1061 = _T_3285 ? _GEN_982 : btb_h_count_2; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1062 = _T_3285 ? _GEN_983 : btb_h_count_3; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1063 = _T_3285 ? _GEN_984 : btb_h_count_4; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1064 = _T_3285 ? _GEN_985 : btb_h_count_5; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1065 = _T_3285 ? _GEN_986 : btb_h_count_6; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1066 = _T_3285 ? _GEN_987 : btb_h_count_7; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1067 = _T_3285 ? _GEN_988 : btb_h_count_8; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1068 = _T_3285 ? _GEN_989 : btb_h_count_9; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1069 = _T_3285 ? _GEN_990 : btb_h_count_10; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1070 = _T_3285 ? _GEN_991 : btb_h_count_11; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1071 = _T_3285 ? _GEN_992 : btb_h_count_12; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1072 = _T_3285 ? _GEN_993 : btb_h_count_13; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1073 = _T_3285 ? _GEN_994 : btb_h_count_14; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1074 = _T_3285 ? _GEN_995 : btb_h_count_15; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1075 = _T_3285 ? _GEN_996 : btb_h_count_16; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1076 = _T_3285 ? _GEN_997 : btb_h_count_17; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1077 = _T_3285 ? _GEN_998 : btb_h_count_18; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1078 = _T_3285 ? _GEN_999 : btb_h_count_19; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1079 = _T_3285 ? _GEN_1000 : btb_h_count_20; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1080 = _T_3285 ? _GEN_1001 : btb_h_count_21; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1081 = _T_3285 ? _GEN_1002 : btb_h_count_22; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1082 = _T_3285 ? _GEN_1003 : btb_h_count_23; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1083 = _T_3285 ? _GEN_1004 : btb_h_count_24; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1084 = _T_3285 ? _GEN_1005 : btb_h_count_25; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1085 = _T_3285 ? _GEN_1006 : btb_h_count_26; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1086 = _T_3285 ? _GEN_1007 : btb_h_count_27; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1087 = _T_3285 ? _GEN_1008 : btb_h_count_28; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1088 = _T_3285 ? _GEN_1009 : btb_h_count_29; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1089 = _T_3285 ? _GEN_1010 : btb_h_count_30; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1090 = _T_3285 ? _GEN_1011 : btb_h_count_31; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1091 = _T_3285 ? _GEN_1012 : btb_h_count_32; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1092 = _T_3285 ? _GEN_1013 : btb_h_count_33; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1093 = _T_3285 ? _GEN_1014 : btb_h_count_34; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1094 = _T_3285 ? _GEN_1015 : btb_h_count_35; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1095 = _T_3285 ? _GEN_1016 : btb_h_count_36; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1096 = _T_3285 ? _GEN_1017 : btb_h_count_37; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1097 = _T_3285 ? _GEN_1018 : btb_h_count_38; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1098 = _T_3285 ? _GEN_1019 : btb_h_count_39; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1099 = _T_3285 ? _GEN_1020 : btb_h_count_40; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1100 = _T_3285 ? _GEN_1021 : btb_h_count_41; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1101 = _T_3285 ? _GEN_1022 : btb_h_count_42; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1102 = _T_3285 ? _GEN_1023 : btb_h_count_43; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1103 = _T_3285 ? _GEN_1024 : btb_h_count_44; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1104 = _T_3285 ? _GEN_1025 : btb_h_count_45; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1105 = _T_3285 ? _GEN_1026 : btb_h_count_46; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1106 = _T_3285 ? _GEN_1027 : btb_h_count_47; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1107 = _T_3285 ? _GEN_1028 : btb_h_count_48; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1108 = _T_3285 ? _GEN_1029 : btb_h_count_49; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1109 = _T_3285 ? _GEN_1030 : btb_h_count_50; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1110 = _T_3285 ? _GEN_1031 : btb_h_count_51; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1111 = _T_3285 ? _GEN_1032 : btb_h_count_52; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1112 = _T_3285 ? _GEN_1033 : btb_h_count_53; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1113 = _T_3285 ? _GEN_1034 : btb_h_count_54; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1114 = _T_3285 ? _GEN_1035 : btb_h_count_55; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1115 = _T_3285 ? _GEN_1036 : btb_h_count_56; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1116 = _T_3285 ? _GEN_1037 : btb_h_count_57; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1117 = _T_3285 ? _GEN_1038 : btb_h_count_58; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1118 = _T_3285 ? _GEN_1039 : btb_h_count_59; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1119 = _T_3285 ? _GEN_1040 : btb_h_count_60; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1120 = _T_3285 ? _GEN_1041 : btb_h_count_61; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1121 = _T_3285 ? _GEN_1042 : btb_h_count_62; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1122 = _T_3285 ? _GEN_1043 : btb_h_count_63; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1125 = _T_3285 ? _GEN_1046 : 1'h0; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1130 = _T_3285 ? _GEN_1051 : 1'h0; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1135 = _T_3285 ? _GEN_1056 : 1'h0; // @[BTB.scala 211:49:@3711.6]
  assign _GEN_1138 = fb_reg_valid ? _GEN_201 : btb_valid_0; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1139 = fb_reg_valid ? _GEN_202 : btb_valid_1; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1140 = fb_reg_valid ? _GEN_203 : btb_valid_2; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1141 = fb_reg_valid ? _GEN_204 : btb_valid_3; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1142 = fb_reg_valid ? _GEN_205 : btb_valid_4; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1143 = fb_reg_valid ? _GEN_206 : btb_valid_5; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1144 = fb_reg_valid ? _GEN_207 : btb_valid_6; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1145 = fb_reg_valid ? _GEN_208 : btb_valid_7; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1146 = fb_reg_valid ? _GEN_209 : btb_valid_8; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1147 = fb_reg_valid ? _GEN_210 : btb_valid_9; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1148 = fb_reg_valid ? _GEN_211 : btb_valid_10; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1149 = fb_reg_valid ? _GEN_212 : btb_valid_11; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1150 = fb_reg_valid ? _GEN_213 : btb_valid_12; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1151 = fb_reg_valid ? _GEN_214 : btb_valid_13; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1152 = fb_reg_valid ? _GEN_215 : btb_valid_14; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1153 = fb_reg_valid ? _GEN_216 : btb_valid_15; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1154 = fb_reg_valid ? _GEN_217 : btb_valid_16; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1155 = fb_reg_valid ? _GEN_218 : btb_valid_17; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1156 = fb_reg_valid ? _GEN_219 : btb_valid_18; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1157 = fb_reg_valid ? _GEN_220 : btb_valid_19; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1158 = fb_reg_valid ? _GEN_221 : btb_valid_20; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1159 = fb_reg_valid ? _GEN_222 : btb_valid_21; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1160 = fb_reg_valid ? _GEN_223 : btb_valid_22; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1161 = fb_reg_valid ? _GEN_224 : btb_valid_23; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1162 = fb_reg_valid ? _GEN_225 : btb_valid_24; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1163 = fb_reg_valid ? _GEN_226 : btb_valid_25; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1164 = fb_reg_valid ? _GEN_227 : btb_valid_26; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1165 = fb_reg_valid ? _GEN_228 : btb_valid_27; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1166 = fb_reg_valid ? _GEN_229 : btb_valid_28; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1167 = fb_reg_valid ? _GEN_230 : btb_valid_29; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1168 = fb_reg_valid ? _GEN_231 : btb_valid_30; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1169 = fb_reg_valid ? _GEN_232 : btb_valid_31; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1170 = fb_reg_valid ? _GEN_233 : btb_valid_32; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1171 = fb_reg_valid ? _GEN_234 : btb_valid_33; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1172 = fb_reg_valid ? _GEN_235 : btb_valid_34; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1173 = fb_reg_valid ? _GEN_236 : btb_valid_35; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1174 = fb_reg_valid ? _GEN_237 : btb_valid_36; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1175 = fb_reg_valid ? _GEN_238 : btb_valid_37; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1176 = fb_reg_valid ? _GEN_239 : btb_valid_38; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1177 = fb_reg_valid ? _GEN_240 : btb_valid_39; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1178 = fb_reg_valid ? _GEN_241 : btb_valid_40; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1179 = fb_reg_valid ? _GEN_242 : btb_valid_41; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1180 = fb_reg_valid ? _GEN_243 : btb_valid_42; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1181 = fb_reg_valid ? _GEN_244 : btb_valid_43; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1182 = fb_reg_valid ? _GEN_245 : btb_valid_44; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1183 = fb_reg_valid ? _GEN_246 : btb_valid_45; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1184 = fb_reg_valid ? _GEN_247 : btb_valid_46; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1185 = fb_reg_valid ? _GEN_248 : btb_valid_47; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1186 = fb_reg_valid ? _GEN_249 : btb_valid_48; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1187 = fb_reg_valid ? _GEN_250 : btb_valid_49; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1188 = fb_reg_valid ? _GEN_251 : btb_valid_50; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1189 = fb_reg_valid ? _GEN_252 : btb_valid_51; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1190 = fb_reg_valid ? _GEN_253 : btb_valid_52; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1191 = fb_reg_valid ? _GEN_254 : btb_valid_53; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1192 = fb_reg_valid ? _GEN_255 : btb_valid_54; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1193 = fb_reg_valid ? _GEN_256 : btb_valid_55; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1194 = fb_reg_valid ? _GEN_257 : btb_valid_56; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1195 = fb_reg_valid ? _GEN_258 : btb_valid_57; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1196 = fb_reg_valid ? _GEN_259 : btb_valid_58; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1197 = fb_reg_valid ? _GEN_260 : btb_valid_59; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1198 = fb_reg_valid ? _GEN_261 : btb_valid_60; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1199 = fb_reg_valid ? _GEN_262 : btb_valid_61; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1200 = fb_reg_valid ? _GEN_263 : btb_valid_62; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1201 = fb_reg_valid ? _GEN_264 : btb_valid_63; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1202 = fb_reg_valid ? _GEN_457 : btb_pc_0; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1203 = fb_reg_valid ? _GEN_458 : btb_pc_1; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1204 = fb_reg_valid ? _GEN_459 : btb_pc_2; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1205 = fb_reg_valid ? _GEN_460 : btb_pc_3; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1206 = fb_reg_valid ? _GEN_461 : btb_pc_4; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1207 = fb_reg_valid ? _GEN_462 : btb_pc_5; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1208 = fb_reg_valid ? _GEN_463 : btb_pc_6; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1209 = fb_reg_valid ? _GEN_464 : btb_pc_7; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1210 = fb_reg_valid ? _GEN_465 : btb_pc_8; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1211 = fb_reg_valid ? _GEN_466 : btb_pc_9; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1212 = fb_reg_valid ? _GEN_467 : btb_pc_10; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1213 = fb_reg_valid ? _GEN_468 : btb_pc_11; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1214 = fb_reg_valid ? _GEN_469 : btb_pc_12; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1215 = fb_reg_valid ? _GEN_470 : btb_pc_13; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1216 = fb_reg_valid ? _GEN_471 : btb_pc_14; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1217 = fb_reg_valid ? _GEN_472 : btb_pc_15; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1218 = fb_reg_valid ? _GEN_473 : btb_pc_16; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1219 = fb_reg_valid ? _GEN_474 : btb_pc_17; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1220 = fb_reg_valid ? _GEN_475 : btb_pc_18; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1221 = fb_reg_valid ? _GEN_476 : btb_pc_19; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1222 = fb_reg_valid ? _GEN_477 : btb_pc_20; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1223 = fb_reg_valid ? _GEN_478 : btb_pc_21; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1224 = fb_reg_valid ? _GEN_479 : btb_pc_22; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1225 = fb_reg_valid ? _GEN_480 : btb_pc_23; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1226 = fb_reg_valid ? _GEN_481 : btb_pc_24; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1227 = fb_reg_valid ? _GEN_482 : btb_pc_25; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1228 = fb_reg_valid ? _GEN_483 : btb_pc_26; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1229 = fb_reg_valid ? _GEN_484 : btb_pc_27; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1230 = fb_reg_valid ? _GEN_485 : btb_pc_28; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1231 = fb_reg_valid ? _GEN_486 : btb_pc_29; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1232 = fb_reg_valid ? _GEN_487 : btb_pc_30; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1233 = fb_reg_valid ? _GEN_488 : btb_pc_31; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1234 = fb_reg_valid ? _GEN_489 : btb_pc_32; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1235 = fb_reg_valid ? _GEN_490 : btb_pc_33; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1236 = fb_reg_valid ? _GEN_491 : btb_pc_34; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1237 = fb_reg_valid ? _GEN_492 : btb_pc_35; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1238 = fb_reg_valid ? _GEN_493 : btb_pc_36; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1239 = fb_reg_valid ? _GEN_494 : btb_pc_37; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1240 = fb_reg_valid ? _GEN_495 : btb_pc_38; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1241 = fb_reg_valid ? _GEN_496 : btb_pc_39; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1242 = fb_reg_valid ? _GEN_497 : btb_pc_40; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1243 = fb_reg_valid ? _GEN_498 : btb_pc_41; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1244 = fb_reg_valid ? _GEN_499 : btb_pc_42; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1245 = fb_reg_valid ? _GEN_500 : btb_pc_43; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1246 = fb_reg_valid ? _GEN_501 : btb_pc_44; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1247 = fb_reg_valid ? _GEN_502 : btb_pc_45; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1248 = fb_reg_valid ? _GEN_503 : btb_pc_46; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1249 = fb_reg_valid ? _GEN_504 : btb_pc_47; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1250 = fb_reg_valid ? _GEN_505 : btb_pc_48; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1251 = fb_reg_valid ? _GEN_506 : btb_pc_49; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1252 = fb_reg_valid ? _GEN_507 : btb_pc_50; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1253 = fb_reg_valid ? _GEN_508 : btb_pc_51; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1254 = fb_reg_valid ? _GEN_509 : btb_pc_52; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1255 = fb_reg_valid ? _GEN_510 : btb_pc_53; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1256 = fb_reg_valid ? _GEN_511 : btb_pc_54; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1257 = fb_reg_valid ? _GEN_512 : btb_pc_55; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1258 = fb_reg_valid ? _GEN_513 : btb_pc_56; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1259 = fb_reg_valid ? _GEN_514 : btb_pc_57; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1260 = fb_reg_valid ? _GEN_515 : btb_pc_58; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1261 = fb_reg_valid ? _GEN_516 : btb_pc_59; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1262 = fb_reg_valid ? _GEN_517 : btb_pc_60; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1263 = fb_reg_valid ? _GEN_518 : btb_pc_61; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1264 = fb_reg_valid ? _GEN_519 : btb_pc_62; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1265 = fb_reg_valid ? _GEN_520 : btb_pc_63; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1266 = fb_reg_valid ? _GEN_521 : btb_tgt_0; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1267 = fb_reg_valid ? _GEN_522 : btb_tgt_1; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1268 = fb_reg_valid ? _GEN_523 : btb_tgt_2; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1269 = fb_reg_valid ? _GEN_524 : btb_tgt_3; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1270 = fb_reg_valid ? _GEN_525 : btb_tgt_4; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1271 = fb_reg_valid ? _GEN_526 : btb_tgt_5; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1272 = fb_reg_valid ? _GEN_527 : btb_tgt_6; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1273 = fb_reg_valid ? _GEN_528 : btb_tgt_7; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1274 = fb_reg_valid ? _GEN_529 : btb_tgt_8; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1275 = fb_reg_valid ? _GEN_530 : btb_tgt_9; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1276 = fb_reg_valid ? _GEN_531 : btb_tgt_10; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1277 = fb_reg_valid ? _GEN_532 : btb_tgt_11; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1278 = fb_reg_valid ? _GEN_533 : btb_tgt_12; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1279 = fb_reg_valid ? _GEN_534 : btb_tgt_13; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1280 = fb_reg_valid ? _GEN_535 : btb_tgt_14; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1281 = fb_reg_valid ? _GEN_536 : btb_tgt_15; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1282 = fb_reg_valid ? _GEN_537 : btb_tgt_16; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1283 = fb_reg_valid ? _GEN_538 : btb_tgt_17; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1284 = fb_reg_valid ? _GEN_539 : btb_tgt_18; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1285 = fb_reg_valid ? _GEN_540 : btb_tgt_19; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1286 = fb_reg_valid ? _GEN_541 : btb_tgt_20; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1287 = fb_reg_valid ? _GEN_542 : btb_tgt_21; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1288 = fb_reg_valid ? _GEN_543 : btb_tgt_22; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1289 = fb_reg_valid ? _GEN_544 : btb_tgt_23; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1290 = fb_reg_valid ? _GEN_545 : btb_tgt_24; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1291 = fb_reg_valid ? _GEN_546 : btb_tgt_25; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1292 = fb_reg_valid ? _GEN_547 : btb_tgt_26; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1293 = fb_reg_valid ? _GEN_548 : btb_tgt_27; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1294 = fb_reg_valid ? _GEN_549 : btb_tgt_28; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1295 = fb_reg_valid ? _GEN_550 : btb_tgt_29; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1296 = fb_reg_valid ? _GEN_551 : btb_tgt_30; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1297 = fb_reg_valid ? _GEN_552 : btb_tgt_31; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1298 = fb_reg_valid ? _GEN_553 : btb_tgt_32; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1299 = fb_reg_valid ? _GEN_554 : btb_tgt_33; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1300 = fb_reg_valid ? _GEN_555 : btb_tgt_34; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1301 = fb_reg_valid ? _GEN_556 : btb_tgt_35; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1302 = fb_reg_valid ? _GEN_557 : btb_tgt_36; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1303 = fb_reg_valid ? _GEN_558 : btb_tgt_37; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1304 = fb_reg_valid ? _GEN_559 : btb_tgt_38; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1305 = fb_reg_valid ? _GEN_560 : btb_tgt_39; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1306 = fb_reg_valid ? _GEN_561 : btb_tgt_40; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1307 = fb_reg_valid ? _GEN_562 : btb_tgt_41; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1308 = fb_reg_valid ? _GEN_563 : btb_tgt_42; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1309 = fb_reg_valid ? _GEN_564 : btb_tgt_43; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1310 = fb_reg_valid ? _GEN_565 : btb_tgt_44; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1311 = fb_reg_valid ? _GEN_566 : btb_tgt_45; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1312 = fb_reg_valid ? _GEN_567 : btb_tgt_46; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1313 = fb_reg_valid ? _GEN_568 : btb_tgt_47; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1314 = fb_reg_valid ? _GEN_569 : btb_tgt_48; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1315 = fb_reg_valid ? _GEN_570 : btb_tgt_49; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1316 = fb_reg_valid ? _GEN_571 : btb_tgt_50; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1317 = fb_reg_valid ? _GEN_572 : btb_tgt_51; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1318 = fb_reg_valid ? _GEN_573 : btb_tgt_52; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1319 = fb_reg_valid ? _GEN_574 : btb_tgt_53; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1320 = fb_reg_valid ? _GEN_575 : btb_tgt_54; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1321 = fb_reg_valid ? _GEN_576 : btb_tgt_55; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1322 = fb_reg_valid ? _GEN_577 : btb_tgt_56; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1323 = fb_reg_valid ? _GEN_578 : btb_tgt_57; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1324 = fb_reg_valid ? _GEN_579 : btb_tgt_58; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1325 = fb_reg_valid ? _GEN_580 : btb_tgt_59; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1326 = fb_reg_valid ? _GEN_581 : btb_tgt_60; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1327 = fb_reg_valid ? _GEN_582 : btb_tgt_61; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1328 = fb_reg_valid ? _GEN_583 : btb_tgt_62; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1329 = fb_reg_valid ? _GEN_584 : btb_tgt_63; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1330 = fb_reg_valid ? _GEN_585 : btb_bj_type_0; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1331 = fb_reg_valid ? _GEN_586 : btb_bj_type_1; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1332 = fb_reg_valid ? _GEN_587 : btb_bj_type_2; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1333 = fb_reg_valid ? _GEN_588 : btb_bj_type_3; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1334 = fb_reg_valid ? _GEN_589 : btb_bj_type_4; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1335 = fb_reg_valid ? _GEN_590 : btb_bj_type_5; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1336 = fb_reg_valid ? _GEN_591 : btb_bj_type_6; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1337 = fb_reg_valid ? _GEN_592 : btb_bj_type_7; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1338 = fb_reg_valid ? _GEN_593 : btb_bj_type_8; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1339 = fb_reg_valid ? _GEN_594 : btb_bj_type_9; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1340 = fb_reg_valid ? _GEN_595 : btb_bj_type_10; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1341 = fb_reg_valid ? _GEN_596 : btb_bj_type_11; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1342 = fb_reg_valid ? _GEN_597 : btb_bj_type_12; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1343 = fb_reg_valid ? _GEN_598 : btb_bj_type_13; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1344 = fb_reg_valid ? _GEN_599 : btb_bj_type_14; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1345 = fb_reg_valid ? _GEN_600 : btb_bj_type_15; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1346 = fb_reg_valid ? _GEN_601 : btb_bj_type_16; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1347 = fb_reg_valid ? _GEN_602 : btb_bj_type_17; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1348 = fb_reg_valid ? _GEN_603 : btb_bj_type_18; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1349 = fb_reg_valid ? _GEN_604 : btb_bj_type_19; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1350 = fb_reg_valid ? _GEN_605 : btb_bj_type_20; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1351 = fb_reg_valid ? _GEN_606 : btb_bj_type_21; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1352 = fb_reg_valid ? _GEN_607 : btb_bj_type_22; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1353 = fb_reg_valid ? _GEN_608 : btb_bj_type_23; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1354 = fb_reg_valid ? _GEN_609 : btb_bj_type_24; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1355 = fb_reg_valid ? _GEN_610 : btb_bj_type_25; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1356 = fb_reg_valid ? _GEN_611 : btb_bj_type_26; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1357 = fb_reg_valid ? _GEN_612 : btb_bj_type_27; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1358 = fb_reg_valid ? _GEN_613 : btb_bj_type_28; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1359 = fb_reg_valid ? _GEN_614 : btb_bj_type_29; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1360 = fb_reg_valid ? _GEN_615 : btb_bj_type_30; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1361 = fb_reg_valid ? _GEN_616 : btb_bj_type_31; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1362 = fb_reg_valid ? _GEN_617 : btb_bj_type_32; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1363 = fb_reg_valid ? _GEN_618 : btb_bj_type_33; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1364 = fb_reg_valid ? _GEN_619 : btb_bj_type_34; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1365 = fb_reg_valid ? _GEN_620 : btb_bj_type_35; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1366 = fb_reg_valid ? _GEN_621 : btb_bj_type_36; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1367 = fb_reg_valid ? _GEN_622 : btb_bj_type_37; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1368 = fb_reg_valid ? _GEN_623 : btb_bj_type_38; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1369 = fb_reg_valid ? _GEN_624 : btb_bj_type_39; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1370 = fb_reg_valid ? _GEN_625 : btb_bj_type_40; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1371 = fb_reg_valid ? _GEN_626 : btb_bj_type_41; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1372 = fb_reg_valid ? _GEN_627 : btb_bj_type_42; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1373 = fb_reg_valid ? _GEN_628 : btb_bj_type_43; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1374 = fb_reg_valid ? _GEN_629 : btb_bj_type_44; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1375 = fb_reg_valid ? _GEN_630 : btb_bj_type_45; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1376 = fb_reg_valid ? _GEN_631 : btb_bj_type_46; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1377 = fb_reg_valid ? _GEN_632 : btb_bj_type_47; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1378 = fb_reg_valid ? _GEN_633 : btb_bj_type_48; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1379 = fb_reg_valid ? _GEN_634 : btb_bj_type_49; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1380 = fb_reg_valid ? _GEN_635 : btb_bj_type_50; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1381 = fb_reg_valid ? _GEN_636 : btb_bj_type_51; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1382 = fb_reg_valid ? _GEN_637 : btb_bj_type_52; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1383 = fb_reg_valid ? _GEN_638 : btb_bj_type_53; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1384 = fb_reg_valid ? _GEN_639 : btb_bj_type_54; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1385 = fb_reg_valid ? _GEN_640 : btb_bj_type_55; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1386 = fb_reg_valid ? _GEN_641 : btb_bj_type_56; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1387 = fb_reg_valid ? _GEN_642 : btb_bj_type_57; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1388 = fb_reg_valid ? _GEN_643 : btb_bj_type_58; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1389 = fb_reg_valid ? _GEN_644 : btb_bj_type_59; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1390 = fb_reg_valid ? _GEN_645 : btb_bj_type_60; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1391 = fb_reg_valid ? _GEN_646 : btb_bj_type_61; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1392 = fb_reg_valid ? _GEN_647 : btb_bj_type_62; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1393 = fb_reg_valid ? _GEN_648 : btb_bj_type_63; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1394 = fb_reg_valid ? _GEN_1059 : btb_h_count_0; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1395 = fb_reg_valid ? _GEN_1060 : btb_h_count_1; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1396 = fb_reg_valid ? _GEN_1061 : btb_h_count_2; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1397 = fb_reg_valid ? _GEN_1062 : btb_h_count_3; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1398 = fb_reg_valid ? _GEN_1063 : btb_h_count_4; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1399 = fb_reg_valid ? _GEN_1064 : btb_h_count_5; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1400 = fb_reg_valid ? _GEN_1065 : btb_h_count_6; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1401 = fb_reg_valid ? _GEN_1066 : btb_h_count_7; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1402 = fb_reg_valid ? _GEN_1067 : btb_h_count_8; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1403 = fb_reg_valid ? _GEN_1068 : btb_h_count_9; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1404 = fb_reg_valid ? _GEN_1069 : btb_h_count_10; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1405 = fb_reg_valid ? _GEN_1070 : btb_h_count_11; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1406 = fb_reg_valid ? _GEN_1071 : btb_h_count_12; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1407 = fb_reg_valid ? _GEN_1072 : btb_h_count_13; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1408 = fb_reg_valid ? _GEN_1073 : btb_h_count_14; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1409 = fb_reg_valid ? _GEN_1074 : btb_h_count_15; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1410 = fb_reg_valid ? _GEN_1075 : btb_h_count_16; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1411 = fb_reg_valid ? _GEN_1076 : btb_h_count_17; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1412 = fb_reg_valid ? _GEN_1077 : btb_h_count_18; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1413 = fb_reg_valid ? _GEN_1078 : btb_h_count_19; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1414 = fb_reg_valid ? _GEN_1079 : btb_h_count_20; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1415 = fb_reg_valid ? _GEN_1080 : btb_h_count_21; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1416 = fb_reg_valid ? _GEN_1081 : btb_h_count_22; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1417 = fb_reg_valid ? _GEN_1082 : btb_h_count_23; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1418 = fb_reg_valid ? _GEN_1083 : btb_h_count_24; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1419 = fb_reg_valid ? _GEN_1084 : btb_h_count_25; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1420 = fb_reg_valid ? _GEN_1085 : btb_h_count_26; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1421 = fb_reg_valid ? _GEN_1086 : btb_h_count_27; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1422 = fb_reg_valid ? _GEN_1087 : btb_h_count_28; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1423 = fb_reg_valid ? _GEN_1088 : btb_h_count_29; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1424 = fb_reg_valid ? _GEN_1089 : btb_h_count_30; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1425 = fb_reg_valid ? _GEN_1090 : btb_h_count_31; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1426 = fb_reg_valid ? _GEN_1091 : btb_h_count_32; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1427 = fb_reg_valid ? _GEN_1092 : btb_h_count_33; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1428 = fb_reg_valid ? _GEN_1093 : btb_h_count_34; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1429 = fb_reg_valid ? _GEN_1094 : btb_h_count_35; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1430 = fb_reg_valid ? _GEN_1095 : btb_h_count_36; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1431 = fb_reg_valid ? _GEN_1096 : btb_h_count_37; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1432 = fb_reg_valid ? _GEN_1097 : btb_h_count_38; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1433 = fb_reg_valid ? _GEN_1098 : btb_h_count_39; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1434 = fb_reg_valid ? _GEN_1099 : btb_h_count_40; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1435 = fb_reg_valid ? _GEN_1100 : btb_h_count_41; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1436 = fb_reg_valid ? _GEN_1101 : btb_h_count_42; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1437 = fb_reg_valid ? _GEN_1102 : btb_h_count_43; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1438 = fb_reg_valid ? _GEN_1103 : btb_h_count_44; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1439 = fb_reg_valid ? _GEN_1104 : btb_h_count_45; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1440 = fb_reg_valid ? _GEN_1105 : btb_h_count_46; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1441 = fb_reg_valid ? _GEN_1106 : btb_h_count_47; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1442 = fb_reg_valid ? _GEN_1107 : btb_h_count_48; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1443 = fb_reg_valid ? _GEN_1108 : btb_h_count_49; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1444 = fb_reg_valid ? _GEN_1109 : btb_h_count_50; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1445 = fb_reg_valid ? _GEN_1110 : btb_h_count_51; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1446 = fb_reg_valid ? _GEN_1111 : btb_h_count_52; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1447 = fb_reg_valid ? _GEN_1112 : btb_h_count_53; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1448 = fb_reg_valid ? _GEN_1113 : btb_h_count_54; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1449 = fb_reg_valid ? _GEN_1114 : btb_h_count_55; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1450 = fb_reg_valid ? _GEN_1115 : btb_h_count_56; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1451 = fb_reg_valid ? _GEN_1116 : btb_h_count_57; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1452 = fb_reg_valid ? _GEN_1117 : btb_h_count_58; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1453 = fb_reg_valid ? _GEN_1118 : btb_h_count_59; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1454 = fb_reg_valid ? _GEN_1119 : btb_h_count_60; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1455 = fb_reg_valid ? _GEN_1120 : btb_h_count_61; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1456 = fb_reg_valid ? _GEN_1121 : btb_h_count_62; // @[BTB.scala 199:23:@3695.4]
  assign _GEN_1457 = fb_reg_valid ? _GEN_1122 : btb_h_count_63; // @[BTB.scala 199:23:@3695.4]
  assign _T_3331 = fb_reg_miss & _T_2925; // @[BTB.scala 227:21:@3760.4]
  assign feedback_select = arb__T_3280_data; // @[BTB.scala 184:22:@2953.4 BTB.scala 197:20:@3694.4]
  assign _T_3333 = feedback_select == 1'h0; // @[BTB.scala 228:26:@3762.6]
  assign _T_3334 = fb_reg_diff & _T_3333; // @[BTB.scala 228:23:@3763.6]
  assign _GEN_1479 = _T_3334 ? 1'h0 : 1'h1; // @[BTB.scala 228:44:@3764.6]
  assign _T_3342 = {_T_175,1'h0,2'h0}; // @[Cat.scala 30:58:@3775.6]
  assign _T_3352 = predict_0_lookup[63:32]; // @[OneHot.scala 26:18:@3783.6]
  assign _T_3353 = predict_0_lookup[31:0]; // @[OneHot.scala 27:18:@3784.6]
  assign _T_3355 = _T_3352 != 32'h0; // @[OneHot.scala 28:14:@3785.6]
  assign _T_3356 = _T_3352 | _T_3353; // @[OneHot.scala 28:28:@3786.6]
  assign _T_3357 = _T_3356[31:16]; // @[OneHot.scala 26:18:@3787.6]
  assign _T_3358 = _T_3356[15:0]; // @[OneHot.scala 27:18:@3788.6]
  assign _T_3360 = _T_3357 != 16'h0; // @[OneHot.scala 28:14:@3789.6]
  assign _T_3361 = _T_3357 | _T_3358; // @[OneHot.scala 28:28:@3790.6]
  assign _T_3362 = _T_3361[15:8]; // @[OneHot.scala 26:18:@3791.6]
  assign _T_3363 = _T_3361[7:0]; // @[OneHot.scala 27:18:@3792.6]
  assign _T_3365 = _T_3362 != 8'h0; // @[OneHot.scala 28:14:@3793.6]
  assign _T_3366 = _T_3362 | _T_3363; // @[OneHot.scala 28:28:@3794.6]
  assign _T_3367 = _T_3366[7:4]; // @[OneHot.scala 26:18:@3795.6]
  assign _T_3368 = _T_3366[3:0]; // @[OneHot.scala 27:18:@3796.6]
  assign _T_3370 = _T_3367 != 4'h0; // @[OneHot.scala 28:14:@3797.6]
  assign _T_3371 = _T_3367 | _T_3368; // @[OneHot.scala 28:28:@3798.6]
  assign _T_3372 = _T_3371[3:2]; // @[OneHot.scala 26:18:@3799.6]
  assign _T_3373 = _T_3371[1:0]; // @[OneHot.scala 27:18:@3800.6]
  assign _T_3375 = _T_3372 != 2'h0; // @[OneHot.scala 28:14:@3801.6]
  assign _T_3376 = _T_3372 | _T_3373; // @[OneHot.scala 28:28:@3802.6]
  assign _T_3377 = _T_3376[1]; // @[CircuitMath.scala 30:8:@3803.6]
  assign _T_3382 = {_T_3355,_T_3360,_T_3365,_T_3370,_T_3375,_T_3377}; // @[Cat.scala 30:58:@3808.6]
  assign _T_3385 = reset == 1'h0; // @[BTB.scala 237:13:@3810.6]
  assign _T_3386 = gb_history[0]; // @[BTB.scala 248:50:@3814.6]
  assign _T_3390 = gb_history[1]; // @[BTB.scala 248:50:@3820.6]
  assign _T_3394 = gb_history[2]; // @[BTB.scala 248:50:@3826.6]
  assign _T_3398 = gb_history[3]; // @[BTB.scala 248:50:@3832.6]
  assign _T_3402 = gb_history[4]; // @[BTB.scala 248:50:@3838.6]
  assign _T_3406 = gb_history[5]; // @[BTB.scala 248:50:@3844.6]
  assign _T_3410 = gb_history[6]; // @[BTB.scala 248:50:@3850.6]
  assign _T_3414 = gb_history[7]; // @[BTB.scala 248:50:@3856.6]
  assign _T_3418 = gb_history[8]; // @[BTB.scala 248:50:@3862.6]
  assign _T_3422 = gb_history[9]; // @[BTB.scala 249:28:@3868.6]
  assign _T_3439 = predict_1_lookup[63:32]; // @[OneHot.scala 26:18:@3885.6]
  assign _T_3440 = predict_1_lookup[31:0]; // @[OneHot.scala 27:18:@3886.6]
  assign _T_3442 = _T_3439 != 32'h0; // @[OneHot.scala 28:14:@3887.6]
  assign _T_3443 = _T_3439 | _T_3440; // @[OneHot.scala 28:28:@3888.6]
  assign _T_3444 = _T_3443[31:16]; // @[OneHot.scala 26:18:@3889.6]
  assign _T_3445 = _T_3443[15:0]; // @[OneHot.scala 27:18:@3890.6]
  assign _T_3447 = _T_3444 != 16'h0; // @[OneHot.scala 28:14:@3891.6]
  assign _T_3448 = _T_3444 | _T_3445; // @[OneHot.scala 28:28:@3892.6]
  assign _T_3449 = _T_3448[15:8]; // @[OneHot.scala 26:18:@3893.6]
  assign _T_3450 = _T_3448[7:0]; // @[OneHot.scala 27:18:@3894.6]
  assign _T_3452 = _T_3449 != 8'h0; // @[OneHot.scala 28:14:@3895.6]
  assign _T_3453 = _T_3449 | _T_3450; // @[OneHot.scala 28:28:@3896.6]
  assign _T_3454 = _T_3453[7:4]; // @[OneHot.scala 26:18:@3897.6]
  assign _T_3455 = _T_3453[3:0]; // @[OneHot.scala 27:18:@3898.6]
  assign _T_3457 = _T_3454 != 4'h0; // @[OneHot.scala 28:14:@3899.6]
  assign _T_3458 = _T_3454 | _T_3455; // @[OneHot.scala 28:28:@3900.6]
  assign _T_3459 = _T_3458[3:2]; // @[OneHot.scala 26:18:@3901.6]
  assign _T_3460 = _T_3458[1:0]; // @[OneHot.scala 27:18:@3902.6]
  assign _T_3462 = _T_3459 != 2'h0; // @[OneHot.scala 28:14:@3903.6]
  assign _T_3463 = _T_3459 | _T_3460; // @[OneHot.scala 28:28:@3904.6]
  assign _T_3464 = _T_3463[1]; // @[CircuitMath.scala 30:8:@3905.6]
  assign _T_3469 = {_T_3442,_T_3447,_T_3452,_T_3457,_T_3462,_T_3464}; // @[Cat.scala 30:58:@3910.6]
  assign io_predict_0_redirect = _T_1246 & _T_1254; // @[BTB.scala 116:28:@1967.4]
  assign io_predict_0_history = gb_history; // @[BTB.scala 118:28:@1972.4]
  assign io_predict_0_diff = _T_1241 ^ _T_1242; // @[BTB.scala 117:28:@1971.4]
  assign io_predict_0_tgt = _T_1260 ? RAS_io_peek : _T_1270; // @[BTB.scala 119:28:@1983.4]
  assign io_predict_1_redirect = _T_2323 & _T_2331; // @[BTB.scala 116:28:@2850.4]
  assign io_predict_1_history = gb_history; // @[BTB.scala 118:28:@2855.4]
  assign io_predict_1_diff = _T_2318 ^ _T_2319; // @[BTB.scala 117:28:@2854.4]
  assign io_predict_1_tgt = _T_2337 ? RAS_io_peek : _T_2347; // @[BTB.scala 119:28:@2866.4]
  assign io_split = io_predict_0_redirect & _T_186; // @[BTB.scala 101:12:@1099.4]
  assign RAS_clock = clock; // @[:@760.4]
  assign RAS_reset = reset; // @[:@761.4]
  assign RAS_io_push_valid = io_ras_push_valid; // @[BTB.scala 81:12:@764.4]
  assign RAS_io_push_bits = io_ras_push_bits; // @[BTB.scala 81:12:@763.4]
  assign RAS_io_pop = io_ras_pop; // @[BTB.scala 80:12:@762.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bht[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    arb[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  gb_history = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  btb_valid_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  btb_valid_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  btb_valid_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  btb_valid_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  btb_valid_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  btb_valid_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  btb_valid_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  btb_valid_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  btb_valid_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  btb_valid_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  btb_valid_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  btb_valid_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  btb_valid_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  btb_valid_13 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  btb_valid_14 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  btb_valid_15 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  btb_valid_16 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  btb_valid_17 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  btb_valid_18 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  btb_valid_19 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  btb_valid_20 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  btb_valid_21 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  btb_valid_22 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  btb_valid_23 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  btb_valid_24 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  btb_valid_25 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  btb_valid_26 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  btb_valid_27 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  btb_valid_28 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  btb_valid_29 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  btb_valid_30 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  btb_valid_31 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  btb_valid_32 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  btb_valid_33 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  btb_valid_34 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  btb_valid_35 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  btb_valid_36 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  btb_valid_37 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  btb_valid_38 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  btb_valid_39 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  btb_valid_40 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  btb_valid_41 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  btb_valid_42 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  btb_valid_43 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  btb_valid_44 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  btb_valid_45 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  btb_valid_46 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  btb_valid_47 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  btb_valid_48 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  btb_valid_49 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  btb_valid_50 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  btb_valid_51 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  btb_valid_52 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  btb_valid_53 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  btb_valid_54 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  btb_valid_55 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  btb_valid_56 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  btb_valid_57 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  btb_valid_58 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  btb_valid_59 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  btb_valid_60 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  btb_valid_61 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  btb_valid_62 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  btb_valid_63 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  btb_pc_0 = _RAND_67[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  btb_pc_1 = _RAND_68[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  btb_pc_2 = _RAND_69[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  btb_pc_3 = _RAND_70[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  btb_pc_4 = _RAND_71[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  btb_pc_5 = _RAND_72[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  btb_pc_6 = _RAND_73[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  btb_pc_7 = _RAND_74[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  btb_pc_8 = _RAND_75[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  btb_pc_9 = _RAND_76[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  btb_pc_10 = _RAND_77[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  btb_pc_11 = _RAND_78[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  btb_pc_12 = _RAND_79[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  btb_pc_13 = _RAND_80[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  btb_pc_14 = _RAND_81[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  btb_pc_15 = _RAND_82[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  btb_pc_16 = _RAND_83[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  btb_pc_17 = _RAND_84[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  btb_pc_18 = _RAND_85[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  btb_pc_19 = _RAND_86[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  btb_pc_20 = _RAND_87[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  btb_pc_21 = _RAND_88[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  btb_pc_22 = _RAND_89[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  btb_pc_23 = _RAND_90[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  btb_pc_24 = _RAND_91[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  btb_pc_25 = _RAND_92[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  btb_pc_26 = _RAND_93[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  btb_pc_27 = _RAND_94[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  btb_pc_28 = _RAND_95[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  btb_pc_29 = _RAND_96[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  btb_pc_30 = _RAND_97[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  btb_pc_31 = _RAND_98[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  btb_pc_32 = _RAND_99[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  btb_pc_33 = _RAND_100[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  btb_pc_34 = _RAND_101[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  btb_pc_35 = _RAND_102[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  btb_pc_36 = _RAND_103[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  btb_pc_37 = _RAND_104[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  btb_pc_38 = _RAND_105[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  btb_pc_39 = _RAND_106[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  btb_pc_40 = _RAND_107[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  btb_pc_41 = _RAND_108[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  btb_pc_42 = _RAND_109[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  btb_pc_43 = _RAND_110[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  btb_pc_44 = _RAND_111[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  btb_pc_45 = _RAND_112[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  btb_pc_46 = _RAND_113[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  btb_pc_47 = _RAND_114[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  btb_pc_48 = _RAND_115[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  btb_pc_49 = _RAND_116[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  btb_pc_50 = _RAND_117[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  btb_pc_51 = _RAND_118[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  btb_pc_52 = _RAND_119[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  btb_pc_53 = _RAND_120[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  btb_pc_54 = _RAND_121[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  btb_pc_55 = _RAND_122[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  btb_pc_56 = _RAND_123[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  btb_pc_57 = _RAND_124[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  btb_pc_58 = _RAND_125[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  btb_pc_59 = _RAND_126[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  btb_pc_60 = _RAND_127[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  btb_pc_61 = _RAND_128[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  btb_pc_62 = _RAND_129[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  btb_pc_63 = _RAND_130[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  btb_tgt_0 = _RAND_131[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  btb_tgt_1 = _RAND_132[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  btb_tgt_2 = _RAND_133[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  btb_tgt_3 = _RAND_134[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  btb_tgt_4 = _RAND_135[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  btb_tgt_5 = _RAND_136[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  btb_tgt_6 = _RAND_137[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  btb_tgt_7 = _RAND_138[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  btb_tgt_8 = _RAND_139[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  btb_tgt_9 = _RAND_140[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  btb_tgt_10 = _RAND_141[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  btb_tgt_11 = _RAND_142[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  btb_tgt_12 = _RAND_143[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  btb_tgt_13 = _RAND_144[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  btb_tgt_14 = _RAND_145[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  btb_tgt_15 = _RAND_146[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  btb_tgt_16 = _RAND_147[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  btb_tgt_17 = _RAND_148[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  btb_tgt_18 = _RAND_149[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  btb_tgt_19 = _RAND_150[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  btb_tgt_20 = _RAND_151[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  btb_tgt_21 = _RAND_152[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  btb_tgt_22 = _RAND_153[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  btb_tgt_23 = _RAND_154[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  btb_tgt_24 = _RAND_155[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  btb_tgt_25 = _RAND_156[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  btb_tgt_26 = _RAND_157[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  btb_tgt_27 = _RAND_158[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  btb_tgt_28 = _RAND_159[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  btb_tgt_29 = _RAND_160[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  btb_tgt_30 = _RAND_161[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  btb_tgt_31 = _RAND_162[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  btb_tgt_32 = _RAND_163[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  btb_tgt_33 = _RAND_164[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  btb_tgt_34 = _RAND_165[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  btb_tgt_35 = _RAND_166[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  btb_tgt_36 = _RAND_167[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  btb_tgt_37 = _RAND_168[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  btb_tgt_38 = _RAND_169[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  btb_tgt_39 = _RAND_170[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  btb_tgt_40 = _RAND_171[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  btb_tgt_41 = _RAND_172[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  btb_tgt_42 = _RAND_173[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  btb_tgt_43 = _RAND_174[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  btb_tgt_44 = _RAND_175[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  btb_tgt_45 = _RAND_176[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  btb_tgt_46 = _RAND_177[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  btb_tgt_47 = _RAND_178[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  btb_tgt_48 = _RAND_179[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  btb_tgt_49 = _RAND_180[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  btb_tgt_50 = _RAND_181[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  btb_tgt_51 = _RAND_182[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  btb_tgt_52 = _RAND_183[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  btb_tgt_53 = _RAND_184[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  btb_tgt_54 = _RAND_185[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  btb_tgt_55 = _RAND_186[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  btb_tgt_56 = _RAND_187[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  btb_tgt_57 = _RAND_188[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  btb_tgt_58 = _RAND_189[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  btb_tgt_59 = _RAND_190[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  btb_tgt_60 = _RAND_191[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  btb_tgt_61 = _RAND_192[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  btb_tgt_62 = _RAND_193[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  btb_tgt_63 = _RAND_194[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  btb_bj_type_0 = _RAND_195[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  btb_bj_type_1 = _RAND_196[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  btb_bj_type_2 = _RAND_197[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  btb_bj_type_3 = _RAND_198[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  btb_bj_type_4 = _RAND_199[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  btb_bj_type_5 = _RAND_200[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  btb_bj_type_6 = _RAND_201[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  btb_bj_type_7 = _RAND_202[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  btb_bj_type_8 = _RAND_203[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  btb_bj_type_9 = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  btb_bj_type_10 = _RAND_205[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  btb_bj_type_11 = _RAND_206[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  btb_bj_type_12 = _RAND_207[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  btb_bj_type_13 = _RAND_208[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  btb_bj_type_14 = _RAND_209[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  btb_bj_type_15 = _RAND_210[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  btb_bj_type_16 = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  btb_bj_type_17 = _RAND_212[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  btb_bj_type_18 = _RAND_213[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  btb_bj_type_19 = _RAND_214[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  btb_bj_type_20 = _RAND_215[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  btb_bj_type_21 = _RAND_216[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  btb_bj_type_22 = _RAND_217[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  btb_bj_type_23 = _RAND_218[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  btb_bj_type_24 = _RAND_219[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  btb_bj_type_25 = _RAND_220[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  btb_bj_type_26 = _RAND_221[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  btb_bj_type_27 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  btb_bj_type_28 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  btb_bj_type_29 = _RAND_224[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  btb_bj_type_30 = _RAND_225[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  btb_bj_type_31 = _RAND_226[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  btb_bj_type_32 = _RAND_227[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  btb_bj_type_33 = _RAND_228[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  btb_bj_type_34 = _RAND_229[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  btb_bj_type_35 = _RAND_230[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  btb_bj_type_36 = _RAND_231[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  btb_bj_type_37 = _RAND_232[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  btb_bj_type_38 = _RAND_233[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  btb_bj_type_39 = _RAND_234[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  btb_bj_type_40 = _RAND_235[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  btb_bj_type_41 = _RAND_236[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  btb_bj_type_42 = _RAND_237[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  btb_bj_type_43 = _RAND_238[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  btb_bj_type_44 = _RAND_239[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  btb_bj_type_45 = _RAND_240[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  btb_bj_type_46 = _RAND_241[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  btb_bj_type_47 = _RAND_242[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  btb_bj_type_48 = _RAND_243[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  btb_bj_type_49 = _RAND_244[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  btb_bj_type_50 = _RAND_245[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  btb_bj_type_51 = _RAND_246[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  btb_bj_type_52 = _RAND_247[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  btb_bj_type_53 = _RAND_248[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  btb_bj_type_54 = _RAND_249[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  btb_bj_type_55 = _RAND_250[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  btb_bj_type_56 = _RAND_251[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  btb_bj_type_57 = _RAND_252[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  btb_bj_type_58 = _RAND_253[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  btb_bj_type_59 = _RAND_254[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  btb_bj_type_60 = _RAND_255[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  btb_bj_type_61 = _RAND_256[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  btb_bj_type_62 = _RAND_257[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  btb_bj_type_63 = _RAND_258[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  btb_h_count_0 = _RAND_259[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  btb_h_count_1 = _RAND_260[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  btb_h_count_2 = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  btb_h_count_3 = _RAND_262[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  btb_h_count_4 = _RAND_263[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  btb_h_count_5 = _RAND_264[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  btb_h_count_6 = _RAND_265[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  btb_h_count_7 = _RAND_266[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  btb_h_count_8 = _RAND_267[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  btb_h_count_9 = _RAND_268[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  btb_h_count_10 = _RAND_269[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  btb_h_count_11 = _RAND_270[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  btb_h_count_12 = _RAND_271[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  btb_h_count_13 = _RAND_272[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  btb_h_count_14 = _RAND_273[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  btb_h_count_15 = _RAND_274[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  btb_h_count_16 = _RAND_275[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  btb_h_count_17 = _RAND_276[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  btb_h_count_18 = _RAND_277[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  btb_h_count_19 = _RAND_278[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  btb_h_count_20 = _RAND_279[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  btb_h_count_21 = _RAND_280[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  btb_h_count_22 = _RAND_281[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  btb_h_count_23 = _RAND_282[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  btb_h_count_24 = _RAND_283[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  btb_h_count_25 = _RAND_284[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  btb_h_count_26 = _RAND_285[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  btb_h_count_27 = _RAND_286[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  btb_h_count_28 = _RAND_287[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  btb_h_count_29 = _RAND_288[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  btb_h_count_30 = _RAND_289[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  btb_h_count_31 = _RAND_290[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  btb_h_count_32 = _RAND_291[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  btb_h_count_33 = _RAND_292[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  btb_h_count_34 = _RAND_293[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  btb_h_count_35 = _RAND_294[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  btb_h_count_36 = _RAND_295[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  btb_h_count_37 = _RAND_296[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  btb_h_count_38 = _RAND_297[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  btb_h_count_39 = _RAND_298[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  btb_h_count_40 = _RAND_299[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  btb_h_count_41 = _RAND_300[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  btb_h_count_42 = _RAND_301[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  btb_h_count_43 = _RAND_302[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  btb_h_count_44 = _RAND_303[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  btb_h_count_45 = _RAND_304[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  btb_h_count_46 = _RAND_305[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  btb_h_count_47 = _RAND_306[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  btb_h_count_48 = _RAND_307[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  btb_h_count_49 = _RAND_308[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  btb_h_count_50 = _RAND_309[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  btb_h_count_51 = _RAND_310[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  btb_h_count_52 = _RAND_311[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  btb_h_count_53 = _RAND_312[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  btb_h_count_54 = _RAND_313[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  btb_h_count_55 = _RAND_314[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  btb_h_count_56 = _RAND_315[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  btb_h_count_57 = _RAND_316[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  btb_h_count_58 = _RAND_317[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  btb_h_count_59 = _RAND_318[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  btb_h_count_60 = _RAND_319[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  btb_h_count_61 = _RAND_320[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  btb_h_count_62 = _RAND_321[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  btb_h_count_63 = _RAND_322[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  shift_reg = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  fb_reg_valid = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  fb_reg_miss = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  fb_reg_redirect = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  fb_reg_btb_type = _RAND_327[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  fb_reg_pc = _RAND_328[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  fb_reg_tgt = _RAND_329[29:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  fb_reg_diff = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  fb_reg_gshxor = _RAND_331[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  fb_reg_lfsr = _RAND_332[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(bht__T_3298_en & bht__T_3298_mask) begin
      bht[bht__T_3298_addr] <= bht__T_3298_data; // @[BTB.scala 77:16:@757.4]
    end
    if(bht__T_3316_en & bht__T_3316_mask) begin
      bht[bht__T_3316_addr] <= bht__T_3316_data; // @[BTB.scala 77:16:@757.4]
    end
    if(bht__T_3327_en & bht__T_3327_mask) begin
      bht[bht__T_3327_addr] <= bht__T_3327_data; // @[BTB.scala 77:16:@757.4]
    end
    if(arb__T_3335_en & arb__T_3335_mask) begin
      arb[arb__T_3335_addr] <= arb__T_3335_data; // @[BTB.scala 78:16:@758.4]
    end
    if(arb__T_3337_en & arb__T_3337_mask) begin
      arb[arb__T_3337_addr] <= arb__T_3337_data; // @[BTB.scala 78:16:@758.4]
    end
    if (reset) begin
      gb_history <= 10'h0;
    end else begin
      if (io_fb_pc_valid) begin
        if (_T_2351) begin
          gb_history <= _T_2353;
        end else begin
          gb_history <= io_feedBack_history;
        end
      end else begin
        if (io_if_pc_valid) begin
          if (shift_wire) begin
            gb_history <= _T_2370;
          end else begin
            if (_T_2360) begin
              if (_T_2364) begin
                gb_history <= _T_2384;
              end else begin
                gb_history <= predict_0_history;
              end
            end else begin
              if (_T_2364) begin
                gb_history <= predict_1_history;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_0 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_valid_0 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h0 == feedback_idx) begin
              btb_valid_0 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_1 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_valid_1 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1 == feedback_idx) begin
              btb_valid_1 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_2 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_valid_2 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2 == feedback_idx) begin
              btb_valid_2 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_3 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_valid_3 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3 == feedback_idx) begin
              btb_valid_3 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_4 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_valid_4 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h4 == feedback_idx) begin
              btb_valid_4 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_5 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_valid_5 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h5 == feedback_idx) begin
              btb_valid_5 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_6 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_valid_6 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h6 == feedback_idx) begin
              btb_valid_6 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_7 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_valid_7 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h7 == feedback_idx) begin
              btb_valid_7 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_8 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_valid_8 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h8 == feedback_idx) begin
              btb_valid_8 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_9 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_valid_9 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h9 == feedback_idx) begin
              btb_valid_9 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_10 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_valid_10 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'ha == feedback_idx) begin
              btb_valid_10 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_11 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_valid_11 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'hb == feedback_idx) begin
              btb_valid_11 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_12 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_valid_12 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'hc == feedback_idx) begin
              btb_valid_12 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_13 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_valid_13 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'hd == feedback_idx) begin
              btb_valid_13 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_14 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_valid_14 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'he == feedback_idx) begin
              btb_valid_14 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_15 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_valid_15 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'hf == feedback_idx) begin
              btb_valid_15 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_16 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_valid_16 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h10 == feedback_idx) begin
              btb_valid_16 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_17 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_valid_17 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h11 == feedback_idx) begin
              btb_valid_17 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_18 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_valid_18 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h12 == feedback_idx) begin
              btb_valid_18 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_19 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_valid_19 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h13 == feedback_idx) begin
              btb_valid_19 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_20 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_valid_20 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h14 == feedback_idx) begin
              btb_valid_20 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_21 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_valid_21 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h15 == feedback_idx) begin
              btb_valid_21 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_22 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_valid_22 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h16 == feedback_idx) begin
              btb_valid_22 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_23 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_valid_23 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h17 == feedback_idx) begin
              btb_valid_23 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_24 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_valid_24 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h18 == feedback_idx) begin
              btb_valid_24 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_25 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_valid_25 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h19 == feedback_idx) begin
              btb_valid_25 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_26 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_valid_26 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1a == feedback_idx) begin
              btb_valid_26 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_27 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_valid_27 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1b == feedback_idx) begin
              btb_valid_27 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_28 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_valid_28 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1c == feedback_idx) begin
              btb_valid_28 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_29 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_valid_29 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1d == feedback_idx) begin
              btb_valid_29 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_30 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_valid_30 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1e == feedback_idx) begin
              btb_valid_30 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_31 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_valid_31 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h1f == feedback_idx) begin
              btb_valid_31 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_32 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_valid_32 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h20 == feedback_idx) begin
              btb_valid_32 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_33 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_valid_33 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h21 == feedback_idx) begin
              btb_valid_33 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_34 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_valid_34 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h22 == feedback_idx) begin
              btb_valid_34 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_35 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_valid_35 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h23 == feedback_idx) begin
              btb_valid_35 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_36 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_valid_36 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h24 == feedback_idx) begin
              btb_valid_36 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_37 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_valid_37 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h25 == feedback_idx) begin
              btb_valid_37 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_38 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_valid_38 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h26 == feedback_idx) begin
              btb_valid_38 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_39 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_valid_39 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h27 == feedback_idx) begin
              btb_valid_39 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_40 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_valid_40 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h28 == feedback_idx) begin
              btb_valid_40 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_41 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_valid_41 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h29 == feedback_idx) begin
              btb_valid_41 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_42 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_valid_42 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2a == feedback_idx) begin
              btb_valid_42 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_43 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_valid_43 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2b == feedback_idx) begin
              btb_valid_43 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_44 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_valid_44 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2c == feedback_idx) begin
              btb_valid_44 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_45 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_valid_45 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2d == feedback_idx) begin
              btb_valid_45 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_46 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_valid_46 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2e == feedback_idx) begin
              btb_valid_46 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_47 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_valid_47 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h2f == feedback_idx) begin
              btb_valid_47 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_48 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_valid_48 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h30 == feedback_idx) begin
              btb_valid_48 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_49 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_valid_49 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h31 == feedback_idx) begin
              btb_valid_49 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_50 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_valid_50 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h32 == feedback_idx) begin
              btb_valid_50 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_51 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_valid_51 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h33 == feedback_idx) begin
              btb_valid_51 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_52 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_valid_52 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h34 == feedback_idx) begin
              btb_valid_52 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_53 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_valid_53 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h35 == feedback_idx) begin
              btb_valid_53 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_54 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_valid_54 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h36 == feedback_idx) begin
              btb_valid_54 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_55 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_valid_55 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h37 == feedback_idx) begin
              btb_valid_55 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_56 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_valid_56 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h38 == feedback_idx) begin
              btb_valid_56 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_57 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_valid_57 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h39 == feedback_idx) begin
              btb_valid_57 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_58 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_valid_58 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3a == feedback_idx) begin
              btb_valid_58 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_59 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_valid_59 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3b == feedback_idx) begin
              btb_valid_59 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_60 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_valid_60 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3c == feedback_idx) begin
              btb_valid_60 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_61 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_valid_61 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3d == feedback_idx) begin
              btb_valid_61 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_62 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_valid_62 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3e == feedback_idx) begin
              btb_valid_62 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_63 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_valid_63 <= 1'h1;
          end
        end else begin
          if (_T_2925) begin
            if (6'h3f == feedback_idx) begin
              btb_valid_63 <= _T_3285;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_pc_0 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_pc_0 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_1 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_pc_1 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_2 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_pc_2 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_3 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_pc_3 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_4 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_pc_4 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_5 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_pc_5 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_6 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_pc_6 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_7 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_pc_7 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_8 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_pc_8 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_9 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_pc_9 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_10 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_pc_10 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_11 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_pc_11 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_12 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_pc_12 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_13 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_pc_13 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_14 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_pc_14 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_15 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_pc_15 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_16 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_pc_16 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_17 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_pc_17 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_18 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_pc_18 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_19 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_pc_19 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_20 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_pc_20 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_21 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_pc_21 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_22 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_pc_22 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_23 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_pc_23 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_24 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_pc_24 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_25 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_pc_25 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_26 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_pc_26 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_27 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_pc_27 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_28 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_pc_28 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_29 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_pc_29 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_30 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_pc_30 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_31 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_pc_31 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_32 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_pc_32 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_33 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_pc_33 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_34 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_pc_34 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_35 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_pc_35 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_36 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_pc_36 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_37 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_pc_37 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_38 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_pc_38 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_39 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_pc_39 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_40 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_pc_40 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_41 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_pc_41 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_42 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_pc_42 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_43 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_pc_43 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_44 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_pc_44 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_45 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_pc_45 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_46 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_pc_46 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_47 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_pc_47 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_48 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_pc_48 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_49 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_pc_49 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_50 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_pc_50 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_51 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_pc_51 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_52 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_pc_52 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_53 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_pc_53 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_54 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_pc_54 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_55 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_pc_55 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_56 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_pc_56 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_57 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_pc_57 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_58 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_pc_58 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_59 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_pc_59 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_60 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_pc_60 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_61 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_pc_61 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_62 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_pc_62 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_63 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_pc_63 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_0 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_tgt_0 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_1 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_tgt_1 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_2 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_tgt_2 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_3 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_tgt_3 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_4 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_tgt_4 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_5 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_tgt_5 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_6 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_tgt_6 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_7 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_tgt_7 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_8 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_tgt_8 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_9 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_tgt_9 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_10 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_tgt_10 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_11 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_tgt_11 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_12 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_tgt_12 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_13 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_tgt_13 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_14 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_tgt_14 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_15 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_tgt_15 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_16 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_tgt_16 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_17 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_tgt_17 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_18 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_tgt_18 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_19 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_tgt_19 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_20 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_tgt_20 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_21 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_tgt_21 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_22 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_tgt_22 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_23 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_tgt_23 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_24 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_tgt_24 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_25 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_tgt_25 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_26 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_tgt_26 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_27 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_tgt_27 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_28 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_tgt_28 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_29 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_tgt_29 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_30 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_tgt_30 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_31 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_tgt_31 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_32 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_tgt_32 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_33 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_tgt_33 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_34 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_tgt_34 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_35 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_tgt_35 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_36 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_tgt_36 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_37 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_tgt_37 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_38 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_tgt_38 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_39 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_tgt_39 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_40 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_tgt_40 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_41 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_tgt_41 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_42 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_tgt_42 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_43 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_tgt_43 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_44 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_tgt_44 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_45 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_tgt_45 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_46 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_tgt_46 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_47 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_tgt_47 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_48 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_tgt_48 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_49 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_tgt_49 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_50 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_tgt_50 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_51 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_tgt_51 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_52 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_tgt_52 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_53 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_tgt_53 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_54 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_tgt_54 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_55 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_tgt_55 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_56 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_tgt_56 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_57 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_tgt_57 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_58 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_tgt_58 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_59 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_tgt_59 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_60 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_tgt_60 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_61 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_tgt_61 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_62 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_tgt_62 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_63 <= 30'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_tgt_63 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_bj_type_0 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_bj_type_1 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_bj_type_2 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_bj_type_3 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_bj_type_4 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_bj_type_5 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_bj_type_6 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_bj_type_7 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_bj_type_8 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_bj_type_9 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_bj_type_10 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_bj_type_11 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_bj_type_12 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_bj_type_13 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_bj_type_14 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_bj_type_15 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_bj_type_16 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_bj_type_17 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_bj_type_18 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_bj_type_19 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_bj_type_20 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_bj_type_21 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_bj_type_22 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_bj_type_23 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_bj_type_24 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_bj_type_25 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_bj_type_26 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_bj_type_27 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_bj_type_28 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_bj_type_29 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_bj_type_30 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_bj_type_31 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_bj_type_32 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_bj_type_33 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_bj_type_34 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_bj_type_35 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_bj_type_36 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_bj_type_37 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_bj_type_38 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_bj_type_39 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_bj_type_40 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_bj_type_41 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_bj_type_42 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_bj_type_43 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_bj_type_44 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_bj_type_45 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_bj_type_46 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_bj_type_47 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_bj_type_48 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_bj_type_49 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_bj_type_50 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_bj_type_51 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_bj_type_52 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_bj_type_53 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_bj_type_54 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_bj_type_55 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_bj_type_56 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_bj_type_57 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_bj_type_58 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_bj_type_59 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_bj_type_60 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_bj_type_61 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_bj_type_62 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_bj_type_63 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= _T_3297;
              end
            end else begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= _T_3297;
              end
            end else begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= _T_3297;
              end
            end else begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= _T_3297;
              end
            end else begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= _T_3297;
              end
            end else begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= _T_3297;
              end
            end else begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= _T_3297;
              end
            end else begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= _T_3297;
              end
            end else begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= _T_3297;
              end
            end else begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= _T_3297;
              end
            end else begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= _T_3297;
              end
            end else begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= _T_3297;
              end
            end else begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= _T_3297;
              end
            end else begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= _T_3297;
              end
            end else begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= _T_3297;
              end
            end else begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= _T_3297;
              end
            end else begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= _T_3297;
              end
            end else begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= _T_3297;
              end
            end else begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= _T_3297;
              end
            end else begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= _T_3297;
              end
            end else begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= _T_3297;
              end
            end else begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= _T_3297;
              end
            end else begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= _T_3297;
              end
            end else begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= _T_3297;
              end
            end else begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= _T_3297;
              end
            end else begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= _T_3297;
              end
            end else begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= _T_3297;
              end
            end else begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= _T_3297;
              end
            end else begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= _T_3297;
              end
            end else begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= _T_3297;
              end
            end else begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= _T_3297;
              end
            end else begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= _T_3297;
              end
            end else begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= _T_3297;
              end
            end else begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= _T_3297;
              end
            end else begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= _T_3297;
              end
            end else begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= _T_3297;
              end
            end else begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= _T_3297;
              end
            end else begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= _T_3297;
              end
            end else begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= _T_3297;
              end
            end else begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= _T_3297;
              end
            end else begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= _T_3297;
              end
            end else begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= _T_3297;
              end
            end else begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= _T_3297;
              end
            end else begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= _T_3297;
              end
            end else begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= _T_3297;
              end
            end else begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= _T_3297;
              end
            end else begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= _T_3297;
              end
            end else begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= _T_3297;
              end
            end else begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= _T_3297;
              end
            end else begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= _T_3297;
              end
            end else begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= _T_3297;
              end
            end else begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= _T_3297;
              end
            end else begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= _T_3297;
              end
            end else begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= _T_3297;
              end
            end else begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= _T_3297;
              end
            end else begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= _T_3297;
              end
            end else begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= _T_3297;
              end
            end else begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= _T_3297;
              end
            end else begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= _T_3297;
              end
            end else begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= _T_3297;
              end
            end else begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= _T_3297;
              end
            end else begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= _T_3297;
              end
            end else begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= _T_3297;
              end
            end else begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_3285) begin
          if (_T_2925) begin
            if (fb_reg_redirect) begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= _T_3297;
              end
            end else begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= _T_3315;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (!(io_fb_pc_valid)) begin
      if (io_if_pc_valid) begin
        shift_reg <= _T_2367;
      end
    end
    if (reset) begin
      fb_reg_valid <= 1'h0;
    end else begin
      fb_reg_valid <= io_feedBack_valid;
    end
    if (reset) begin
      fb_reg_miss <= 1'h0;
    end else begin
      fb_reg_miss <= io_fb_pc_valid;
    end
    if (reset) begin
      fb_reg_redirect <= 1'h0;
    end else begin
      fb_reg_redirect <= io_feedBack_redirect;
    end
    if (reset) begin
      fb_reg_btb_type <= 2'h0;
    end else begin
      fb_reg_btb_type <= io_fb_type;
    end
    if (reset) begin
      fb_reg_pc <= 30'h0;
    end else begin
      fb_reg_pc <= _T_2393;
    end
    if (reset) begin
      fb_reg_tgt <= 30'h0;
    end else begin
      fb_reg_tgt <= _T_2394;
    end
    if (reset) begin
      fb_reg_diff <= 1'h0;
    end else begin
      fb_reg_diff <= io_feedBack_diff;
    end
    if (reset) begin
      fb_reg_gshxor <= 10'h0;
    end else begin
      fb_reg_gshxor <= _T_2397;
    end
    if (reset) begin
      fb_reg_lfsr <= 6'h1;
    end else begin
      fb_reg_lfsr <= _T_2402;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002,"BTB: Cyc= %d valid %x pc %x redirect %x index %d select %d gshare %d hcount %d bhtIdx %d <",io_cyc,io_if_pc_valid,_T_3342,_T_1255,_T_3382,predict_0_select,predict_0_gshare,predict_0_h_count,predict_0_gshxor); // @[BTB.scala 237:13:@3812.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3386); // @[BTB.scala 248:34:@3818.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3390); // @[BTB.scala 248:34:@3824.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3394); // @[BTB.scala 248:34:@3830.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3398); // @[BTB.scala 248:34:@3836.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3402); // @[BTB.scala 248:34:@3842.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3406); // @[BTB.scala 248:34:@3848.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3410); // @[BTB.scala 248:34:@3854.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3414); // @[BTB.scala 248:34:@3860.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3418); // @[BTB.scala 248:34:@3866.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1246 & _T_3385) begin
          $fwrite(32'h80000002,"%d\n",_T_3422); // @[BTB.scala 249:13:@3872.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002,"BTB: Cyc= %d valid %x pc %x redirect %x index %d select %d gshare %d hcount %d bhtIdx %d <",io_cyc,io_if_pc_valid,predict_0_cont_tgt,_T_2332,_T_3469,predict_1_select,predict_1_gshare,predict_1_h_count,predict_1_gshxor); // @[BTB.scala 237:13:@3914.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3386); // @[BTB.scala 248:34:@3920.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3390); // @[BTB.scala 248:34:@3926.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3394); // @[BTB.scala 248:34:@3932.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3398); // @[BTB.scala 248:34:@3938.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3402); // @[BTB.scala 248:34:@3944.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3406); // @[BTB.scala 248:34:@3950.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3410); // @[BTB.scala 248:34:@3956.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3414); // @[BTB.scala 248:34:@3962.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002," %d",_T_3418); // @[BTB.scala 248:34:@3968.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_2323 & _T_3385) begin
          $fwrite(32'h80000002,"%d\n",_T_3422); // @[BTB.scala 249:13:@3974.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module FetchInst( // @[:@3978.2]
  input         clock, // @[:@3979.4]
  input         reset, // @[:@3980.4]
  input         io_mem_addr_ready, // @[:@3981.4]
  output        io_mem_addr_valid, // @[:@3981.4]
  output [31:0] io_mem_addr_bits, // @[:@3981.4]
  input         io_mem_inst_0_valid, // @[:@3981.4]
  input  [31:0] io_mem_inst_0_bits, // @[:@3981.4]
  input         io_mem_inst_1_valid, // @[:@3981.4]
  input  [31:0] io_mem_inst_1_bits, // @[:@3981.4]
  input         io_if_btb_0_redirect, // @[:@3981.4]
  input  [9:0]  io_if_btb_0_history, // @[:@3981.4]
  input         io_if_btb_0_diff, // @[:@3981.4]
  input  [31:0] io_if_btb_0_tgt, // @[:@3981.4]
  input         io_if_btb_1_redirect, // @[:@3981.4]
  input  [9:0]  io_if_btb_1_history, // @[:@3981.4]
  input         io_if_btb_1_diff, // @[:@3981.4]
  input  [31:0] io_if_btb_1_tgt, // @[:@3981.4]
  output        io_dec_btb_0_redirect, // @[:@3981.4]
  output [9:0]  io_dec_btb_0_history, // @[:@3981.4]
  output        io_dec_btb_0_diff, // @[:@3981.4]
  output [31:0] io_dec_btb_0_tgt, // @[:@3981.4]
  output        io_dec_btb_1_redirect, // @[:@3981.4]
  output [9:0]  io_dec_btb_1_history, // @[:@3981.4]
  output        io_dec_btb_1_diff, // @[:@3981.4]
  output [31:0] io_dec_btb_1_tgt, // @[:@3981.4]
  input  [31:0] io_pc, // @[:@3981.4]
  input         io_pc_split, // @[:@3981.4]
  output        io_pc_forward, // @[:@3981.4]
  input         io_forward_0, // @[:@3981.4]
  input         io_forward_1, // @[:@3981.4]
  input         io_if_kill, // @[:@3981.4]
  input         io_dec_kill, // @[:@3981.4]
  output        io_inst_0_valid, // @[:@3981.4]
  output [31:0] io_inst_0_bits, // @[:@3981.4]
  output        io_inst_1_valid, // @[:@3981.4]
  output [31:0] io_inst_1_bits, // @[:@3981.4]
  output [31:0] io_dec_pc_0, // @[:@3981.4]
  output [31:0] io_dec_pc_1, // @[:@3981.4]
  input         io_inst_split // @[:@3981.4]
);
  reg  inst_odd; // @[FetchInst.scala 39:27:@3987.4]
  reg [31:0] _RAND_0;
  reg  inst_kill; // @[FetchInst.scala 40:27:@3988.4]
  reg [31:0] _RAND_1;
  reg  inst_split; // @[FetchInst.scala 41:27:@3989.4]
  reg [31:0] _RAND_2;
  wire  _T_169; // @[FetchInst.scala 43:44:@3991.4]
  wire  inst_valid_0; // @[FetchInst.scala 43:41:@3992.4]
  reg [1:0] state; // @[FetchInst.scala 47:22:@3995.4]
  reg [31:0] _RAND_3;
  wire  inst_valid_orR; // @[FetchInst.scala 48:49:@3996.4]
  wire  _T_172; // @[FetchInst.scala 49:40:@3997.4]
  wire  _T_173; // @[FetchInst.scala 49:77:@3998.4]
  wire  _T_176; // @[FetchInst.scala 49:98:@4000.4]
  wire  _T_177; // @[FetchInst.scala 49:59:@4001.4]
  wire  if_forward; // @[FetchInst.scala 49:53:@4002.4]
  wire  _T_178; // @[Conditional.scala 37:30:@4003.4]
  wire [1:0] _GEN_0; // @[FetchInst.scala 52:25:@4005.6]
  wire  _T_179; // @[Conditional.scala 37:30:@4010.6]
  wire [1:0] _T_180; // @[FetchInst.scala 57:23:@4014.12]
  wire [1:0] _GEN_1; // @[FetchInst.scala 58:34:@4018.12]
  wire [1:0] _GEN_2; // @[FetchInst.scala 56:26:@4013.10]
  wire [1:0] _GEN_3; // @[FetchInst.scala 55:27:@4012.8]
  wire  _T_181; // @[Conditional.scala 37:30:@4027.8]
  wire [1:0] _GEN_4; // @[FetchInst.scala 65:32:@4034.12]
  wire [1:0] _GEN_5; // @[FetchInst.scala 63:27:@4029.10]
  wire [1:0] _GEN_6; // @[Conditional.scala 39:67:@4028.8]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@4011.6]
  wire [1:0] _GEN_8; // @[Conditional.scala 40:58:@4004.4]
  wire  _T_184; // @[FetchInst.scala 71:35:@4046.8]
  wire  _T_185; // @[FetchInst.scala 71:26:@4047.8]
  wire  _GEN_9; // @[FetchInst.scala 71:50:@4048.8]
  wire  _GEN_10; // @[FetchInst.scala 70:30:@4042.6]
  wire  _T_191; // @[FetchInst.scala 76:21:@4053.4]
  wire  _T_192; // @[FetchInst.scala 77:21:@4054.4]
  wire  _T_193; // @[FetchInst.scala 76:35:@4055.4]
  wire  _T_194; // @[FetchInst.scala 78:12:@4056.4]
  wire  _T_195; // @[FetchInst.scala 78:27:@4057.4]
  wire  pc_valid; // @[FetchInst.scala 77:36:@4058.4]
  wire  _GEN_11; // @[FetchInst.scala 69:19:@4038.4]
  reg  pc_odd_reg; // @[FetchInst.scala 73:27:@4051.4]
  reg [31:0] _RAND_4;
  reg  state_WtForward; // @[FetchInst.scala 74:32:@4052.4]
  reg [31:0] _RAND_5;
  wire  _T_199; // @[FetchInst.scala 81:30:@4061.4]
  wire  _T_200; // @[FetchInst.scala 81:27:@4062.4]
  wire  _T_203; // @[FetchInst.scala 81:45:@4065.4]
  wire  _T_206; // @[FetchInst.scala 83:33:@4068.4]
  wire  _T_207; // @[FetchInst.scala 83:17:@4069.4]
  wire  _T_208; // @[FetchInst.scala 84:38:@4070.4]
  wire  _T_209; // @[FetchInst.scala 84:20:@4071.4]
  wire  _T_210; // @[FetchInst.scala 83:62:@4072.4]
  wire  _T_211; // @[FetchInst.scala 84:55:@4073.4]
  wire  _T_212; // @[FetchInst.scala 82:45:@4074.4]
  wire  _T_213; // @[FetchInst.scala 80:45:@4075.4]
  reg  maintain; // @[FetchInst.scala 86:25:@4078.4]
  reg [31:0] _RAND_6;
  wire  _T_218; // @[FetchInst.scala 87:42:@4079.4]
  wire  _T_219; // @[FetchInst.scala 87:39:@4080.4]
  wire  _T_223; // @[FetchInst.scala 88:39:@4084.4]
  wire  _T_225; // @[FetchInst.scala 88:79:@4086.4]
  wire  _T_226; // @[FetchInst.scala 88:54:@4087.4]
  wire  _T_228; // @[FetchInst.scala 88:96:@4088.4]
  wire  _T_232; // @[FetchInst.scala 90:41:@4092.4]
  wire  _T_235; // @[FetchInst.scala 90:59:@4094.4]
  wire  pc_odd_wire; // @[FetchInst.scala 90:74:@4096.4]
  wire  _GEN_12; // @[FetchInst.scala 92:27:@4101.6]
  wire  _GEN_13; // @[FetchInst.scala 91:21:@4097.4]
  wire  pc_odd_1; // @[FetchInst.scala 96:27:@4109.4]
  wire  pc_odd_0; // @[FetchInst.scala 95:26:@4107.4]
  wire  _T_252; // @[FetchInst.scala 100:21:@4113.4]
  wire  _GEN_14; // @[FetchInst.scala 101:43:@4120.6]
  wire  _GEN_15; // @[FetchInst.scala 100:39:@4114.4]
  wire  _T_258; // @[FetchInst.scala 103:21:@4123.4]
  wire  _T_261; // @[FetchInst.scala 104:35:@4129.6]
  wire  _GEN_16; // @[FetchInst.scala 104:53:@4130.6]
  wire  _GEN_17; // @[FetchInst.scala 103:39:@4124.4]
  reg [31:0] reg_pc_0; // @[FetchInst.scala 108:21:@4133.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_pc_1; // @[FetchInst.scala 108:21:@4133.4]
  reg [31:0] _RAND_8;
  reg  reg_pred_0_redirect; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_9;
  reg [9:0] reg_pred_0_history; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_10;
  reg  reg_pred_0_diff; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_11;
  reg [31:0] reg_pred_0_tgt; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_12;
  reg  reg_pred_1_redirect; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_13;
  reg [9:0] reg_pred_1_history; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_14;
  reg  reg_pred_1_diff; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_15;
  reg [31:0] reg_pred_1_tgt; // @[FetchInst.scala 109:21:@4134.4]
  reg [31:0] _RAND_16;
  wire  _T_278; // @[FetchInst.scala 112:19:@4137.6]
  wire  _T_279; // @[FetchInst.scala 112:30:@4138.6]
  wire [28:0] _T_282; // @[FetchInst.scala 114:49:@4142.8]
  wire [31:0] _T_286; // @[Cat.scala 30:58:@4144.8]
  wire [31:0] _GEN_18; // @[FetchInst.scala 114:25:@4141.6]
  wire [31:0] _GEN_19; // @[FetchInst.scala 114:25:@4141.6]
  wire  _GEN_20; // @[FetchInst.scala 114:25:@4141.6]
  wire [9:0] _GEN_21; // @[FetchInst.scala 114:25:@4141.6]
  wire  _GEN_22; // @[FetchInst.scala 114:25:@4141.6]
  wire  _T_288; // @[FetchInst.scala 114:13:@4151.6]
  wire [31:0] _T_293; // @[Cat.scala 30:58:@4155.8]
  wire [31:0] _GEN_23; // @[FetchInst.scala 114:25:@4152.6]
  wire [31:0] _GEN_24; // @[FetchInst.scala 114:25:@4152.6]
  wire  _GEN_25; // @[FetchInst.scala 114:25:@4152.6]
  wire [9:0] _GEN_26; // @[FetchInst.scala 114:25:@4152.6]
  wire  _GEN_27; // @[FetchInst.scala 114:25:@4152.6]
  wire  _GEN_28; // @[FetchInst.scala 110:19:@4135.4]
  wire  _GEN_29; // @[FetchInst.scala 110:19:@4135.4]
  reg [31:0] _T_375; // @[FetchInst.scala 9:29:@4170.4]
  reg [31:0] _RAND_17;
  wire [31:0] _GEN_40; // @[FetchInst.scala 10:15:@4171.4]
  reg [31:0] _T_378; // @[FetchInst.scala 9:29:@4182.4]
  reg [31:0] _RAND_18;
  wire [31:0] _GEN_41; // @[FetchInst.scala 10:15:@4183.4]
  assign _T_169 = inst_odd == 1'h0; // @[FetchInst.scala 43:44:@3991.4]
  assign inst_valid_0 = io_mem_inst_0_valid & _T_169; // @[FetchInst.scala 43:41:@3992.4]
  assign inst_valid_orR = inst_valid_0 | io_mem_inst_1_valid; // @[FetchInst.scala 48:49:@3996.4]
  assign _T_172 = io_forward_1 | inst_kill; // @[FetchInst.scala 49:40:@3997.4]
  assign _T_173 = io_pc[2]; // @[FetchInst.scala 49:77:@3998.4]
  assign _T_176 = io_mem_inst_1_valid == 1'h0; // @[FetchInst.scala 49:98:@4000.4]
  assign _T_177 = inst_split ? _T_173 : _T_176; // @[FetchInst.scala 49:59:@4001.4]
  assign if_forward = _T_172 | _T_177; // @[FetchInst.scala 49:53:@4002.4]
  assign _T_178 = 2'h0 == state; // @[Conditional.scala 37:30:@4003.4]
  assign _GEN_0 = io_mem_addr_ready ? 2'h1 : state; // @[FetchInst.scala 52:25:@4005.6]
  assign _T_179 = 2'h1 == state; // @[Conditional.scala 37:30:@4010.6]
  assign _T_180 = io_mem_addr_ready ? 2'h1 : 2'h0; // @[FetchInst.scala 57:23:@4014.12]
  assign _GEN_1 = io_dec_kill ? 2'h0 : 2'h2; // @[FetchInst.scala 58:34:@4018.12]
  assign _GEN_2 = if_forward ? _T_180 : _GEN_1; // @[FetchInst.scala 56:26:@4013.10]
  assign _GEN_3 = inst_valid_orR ? _GEN_2 : state; // @[FetchInst.scala 55:27:@4012.8]
  assign _T_181 = 2'h2 == state; // @[Conditional.scala 37:30:@4027.8]
  assign _GEN_4 = io_dec_kill ? 2'h0 : state; // @[FetchInst.scala 65:32:@4034.12]
  assign _GEN_5 = io_forward_1 ? _T_180 : _GEN_4; // @[FetchInst.scala 63:27:@4029.10]
  assign _GEN_6 = _T_181 ? _GEN_5 : state; // @[Conditional.scala 39:67:@4028.8]
  assign _GEN_7 = _T_179 ? _GEN_3 : _GEN_6; // @[Conditional.scala 39:67:@4011.6]
  assign _GEN_8 = _T_178 ? _GEN_0 : _GEN_7; // @[Conditional.scala 40:58:@4004.4]
  assign _T_184 = state == 2'h1; // @[FetchInst.scala 71:35:@4046.8]
  assign _T_185 = io_dec_kill & _T_184; // @[FetchInst.scala 71:26:@4047.8]
  assign _GEN_9 = _T_185 ? 1'h1 : inst_kill; // @[FetchInst.scala 71:50:@4048.8]
  assign _GEN_10 = inst_valid_orR ? 1'h0 : _GEN_9; // @[FetchInst.scala 70:30:@4042.6]
  assign _T_191 = state == 2'h0; // @[FetchInst.scala 76:21:@4053.4]
  assign _T_192 = inst_valid_orR & if_forward; // @[FetchInst.scala 77:21:@4054.4]
  assign _T_193 = _T_191 | _T_192; // @[FetchInst.scala 76:35:@4055.4]
  assign _T_194 = state == 2'h2; // @[FetchInst.scala 78:12:@4056.4]
  assign _T_195 = _T_194 & io_forward_1; // @[FetchInst.scala 78:27:@4057.4]
  assign pc_valid = _T_193 | _T_195; // @[FetchInst.scala 77:36:@4058.4]
  assign _GEN_11 = pc_valid ? io_if_kill : _GEN_10; // @[FetchInst.scala 69:19:@4038.4]
  assign _T_199 = pc_odd_reg == 1'h0; // @[FetchInst.scala 81:30:@4061.4]
  assign _T_200 = _T_191 & _T_199; // @[FetchInst.scala 81:27:@4062.4]
  assign _T_203 = _T_200 | _T_195; // @[FetchInst.scala 81:45:@4065.4]
  assign _T_206 = inst_split & _T_173; // @[FetchInst.scala 83:33:@4068.4]
  assign _T_207 = inst_kill | _T_206; // @[FetchInst.scala 83:17:@4069.4]
  assign _T_208 = io_mem_inst_1_valid | inst_split; // @[FetchInst.scala 84:38:@4070.4]
  assign _T_209 = io_forward_1 & _T_208; // @[FetchInst.scala 84:20:@4071.4]
  assign _T_210 = _T_207 | _T_209; // @[FetchInst.scala 83:62:@4072.4]
  assign _T_211 = _T_210 & inst_valid_orR; // @[FetchInst.scala 84:55:@4073.4]
  assign _T_212 = _T_203 | _T_211; // @[FetchInst.scala 82:45:@4074.4]
  assign _T_213 = io_mem_addr_ready & _T_212; // @[FetchInst.scala 80:45:@4075.4]
  assign _T_218 = inst_kill == 1'h0; // @[FetchInst.scala 87:42:@4079.4]
  assign _T_219 = inst_valid_0 & _T_218; // @[FetchInst.scala 87:39:@4080.4]
  assign _T_223 = io_mem_inst_1_valid & _T_218; // @[FetchInst.scala 88:39:@4084.4]
  assign _T_225 = _T_194 & maintain; // @[FetchInst.scala 88:79:@4086.4]
  assign _T_226 = _T_223 | _T_225; // @[FetchInst.scala 88:54:@4087.4]
  assign _T_228 = inst_split == 1'h0; // @[FetchInst.scala 88:96:@4088.4]
  assign _T_232 = inst_valid_0 & _T_176; // @[FetchInst.scala 90:41:@4092.4]
  assign _T_235 = _T_232 & _T_228; // @[FetchInst.scala 90:59:@4094.4]
  assign pc_odd_wire = _T_235 & _T_218; // @[FetchInst.scala 90:74:@4096.4]
  assign _GEN_12 = pc_odd_wire ? 1'h1 : pc_odd_reg; // @[FetchInst.scala 92:27:@4101.6]
  assign _GEN_13 = io_mem_addr_ready ? 1'h0 : _GEN_12; // @[FetchInst.scala 91:21:@4097.4]
  assign pc_odd_1 = pc_odd_reg | pc_odd_wire; // @[FetchInst.scala 96:27:@4109.4]
  assign pc_odd_0 = pc_odd_1 | _T_173; // @[FetchInst.scala 95:26:@4107.4]
  assign _T_252 = io_dec_kill | io_forward_0; // @[FetchInst.scala 100:21:@4113.4]
  assign _GEN_14 = _T_219 ? 1'h1 : state_WtForward; // @[FetchInst.scala 101:43:@4120.6]
  assign _GEN_15 = _T_252 ? 1'h0 : _GEN_14; // @[FetchInst.scala 100:39:@4114.4]
  assign _T_258 = io_dec_kill | io_forward_1; // @[FetchInst.scala 103:21:@4123.4]
  assign _T_261 = _T_194 & io_inst_split; // @[FetchInst.scala 104:35:@4129.6]
  assign _GEN_16 = _T_261 ? 1'h0 : maintain; // @[FetchInst.scala 104:53:@4130.6]
  assign _GEN_17 = _T_258 ? 1'h1 : _GEN_16; // @[FetchInst.scala 103:39:@4124.4]
  assign _T_278 = pc_odd_0 == 1'h0; // @[FetchInst.scala 112:19:@4137.6]
  assign _T_279 = _T_278 & io_pc_split; // @[FetchInst.scala 112:30:@4138.6]
  assign _T_282 = io_pc[31:3]; // @[FetchInst.scala 114:49:@4142.8]
  assign _T_286 = {_T_282,1'h0,2'h0}; // @[Cat.scala 30:58:@4144.8]
  assign _GEN_18 = _T_278 ? _T_286 : reg_pc_0; // @[FetchInst.scala 114:25:@4141.6]
  assign _GEN_19 = _T_278 ? io_if_btb_0_tgt : reg_pred_0_tgt; // @[FetchInst.scala 114:25:@4141.6]
  assign _GEN_20 = _T_278 ? io_if_btb_0_diff : reg_pred_0_diff; // @[FetchInst.scala 114:25:@4141.6]
  assign _GEN_21 = _T_278 ? io_if_btb_0_history : reg_pred_0_history; // @[FetchInst.scala 114:25:@4141.6]
  assign _GEN_22 = _T_278 ? io_if_btb_0_redirect : reg_pred_0_redirect; // @[FetchInst.scala 114:25:@4141.6]
  assign _T_288 = pc_odd_1 == 1'h0; // @[FetchInst.scala 114:13:@4151.6]
  assign _T_293 = {_T_282,1'h1,2'h0}; // @[Cat.scala 30:58:@4155.8]
  assign _GEN_23 = _T_288 ? _T_293 : reg_pc_1; // @[FetchInst.scala 114:25:@4152.6]
  assign _GEN_24 = _T_288 ? io_if_btb_1_tgt : reg_pred_1_tgt; // @[FetchInst.scala 114:25:@4152.6]
  assign _GEN_25 = _T_288 ? io_if_btb_1_diff : reg_pred_1_diff; // @[FetchInst.scala 114:25:@4152.6]
  assign _GEN_26 = _T_288 ? io_if_btb_1_history : reg_pred_1_history; // @[FetchInst.scala 114:25:@4152.6]
  assign _GEN_27 = _T_288 ? io_if_btb_1_redirect : reg_pred_1_redirect; // @[FetchInst.scala 114:25:@4152.6]
  assign _GEN_28 = pc_valid ? pc_odd_0 : inst_odd; // @[FetchInst.scala 110:19:@4135.4]
  assign _GEN_29 = pc_valid ? _T_279 : inst_split; // @[FetchInst.scala 110:19:@4135.4]
  assign _GEN_40 = inst_valid_0 ? io_mem_inst_0_bits : _T_375; // @[FetchInst.scala 10:15:@4171.4]
  assign _GEN_41 = io_mem_inst_1_valid ? io_mem_inst_1_bits : _T_378; // @[FetchInst.scala 10:15:@4183.4]
  assign io_mem_addr_valid = _T_193 | _T_195; // @[FetchInst.scala 38:21:@3986.4]
  assign io_mem_addr_bits = pc_odd_1 ? io_dec_pc_1 : io_pc; // @[FetchInst.scala 37:20:@3985.4]
  assign io_dec_btb_0_redirect = reg_pred_0_redirect; // @[FetchInst.scala 120:21:@4168.4]
  assign io_dec_btb_0_history = reg_pred_0_history; // @[FetchInst.scala 120:21:@4167.4]
  assign io_dec_btb_0_diff = reg_pred_0_diff; // @[FetchInst.scala 120:21:@4166.4]
  assign io_dec_btb_0_tgt = reg_pred_0_tgt; // @[FetchInst.scala 120:21:@4165.4]
  assign io_dec_btb_1_redirect = reg_pred_1_redirect; // @[FetchInst.scala 120:21:@4180.4]
  assign io_dec_btb_1_history = reg_pred_1_history; // @[FetchInst.scala 120:21:@4179.4]
  assign io_dec_btb_1_diff = reg_pred_1_diff; // @[FetchInst.scala 120:21:@4178.4]
  assign io_dec_btb_1_tgt = reg_pred_1_tgt; // @[FetchInst.scala 120:21:@4177.4]
  assign io_pc_forward = io_if_kill | _T_213; // @[FetchInst.scala 80:17:@4077.4]
  assign io_inst_0_valid = _T_219 | state_WtForward; // @[FetchInst.scala 87:20:@4082.4]
  assign io_inst_0_bits = inst_valid_0 ? io_mem_inst_0_bits : _T_375; // @[FetchInst.scala 122:21:@4175.4]
  assign io_inst_1_valid = _T_226 & _T_228; // @[FetchInst.scala 88:20:@4090.4]
  assign io_inst_1_bits = io_mem_inst_1_valid ? io_mem_inst_1_bits : _T_378; // @[FetchInst.scala 122:21:@4187.4]
  assign io_dec_pc_0 = reg_pc_0; // @[FetchInst.scala 121:21:@4169.4]
  assign io_dec_pc_1 = reg_pc_1; // @[FetchInst.scala 121:21:@4181.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  inst_odd = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inst_kill = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inst_split = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  state = _RAND_3[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  pc_odd_reg = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  state_WtForward = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  maintain = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_pc_0 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_pc_1 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_pred_0_redirect = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_pred_0_history = _RAND_10[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_pred_0_diff = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  reg_pred_0_tgt = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  reg_pred_1_redirect = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  reg_pred_1_history = _RAND_14[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  reg_pred_1_diff = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  reg_pred_1_tgt = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  _T_375 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  _T_378 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      inst_odd <= 1'h0;
    end else begin
      if (pc_valid) begin
        inst_odd <= pc_odd_0;
      end
    end
    if (reset) begin
      inst_kill <= 1'h0;
    end else begin
      if (pc_valid) begin
        inst_kill <= io_if_kill;
      end else begin
        if (inst_valid_orR) begin
          inst_kill <= 1'h0;
        end else begin
          if (_T_185) begin
            inst_kill <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      inst_split <= 1'h0;
    end else begin
      if (pc_valid) begin
        inst_split <= _T_279;
      end
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_178) begin
        if (io_mem_addr_ready) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_179) begin
          if (inst_valid_orR) begin
            if (if_forward) begin
              if (io_mem_addr_ready) begin
                state <= 2'h1;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (io_dec_kill) begin
                state <= 2'h0;
              end else begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_181) begin
            if (io_forward_1) begin
              if (io_mem_addr_ready) begin
                state <= 2'h1;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (io_dec_kill) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      pc_odd_reg <= 1'h0;
    end else begin
      if (io_mem_addr_ready) begin
        pc_odd_reg <= 1'h0;
      end else begin
        if (pc_odd_wire) begin
          pc_odd_reg <= 1'h1;
        end
      end
    end
    if (reset) begin
      state_WtForward <= 1'h0;
    end else begin
      if (_T_252) begin
        state_WtForward <= 1'h0;
      end else begin
        if (_T_219) begin
          state_WtForward <= 1'h1;
        end
      end
    end
    if (reset) begin
      maintain <= 1'h1;
    end else begin
      if (_T_258) begin
        maintain <= 1'h1;
      end else begin
        if (_T_261) begin
          maintain <= 1'h0;
        end
      end
    end
    if (pc_valid) begin
      if (_T_278) begin
        reg_pc_0 <= _T_286;
      end
    end
    if (pc_valid) begin
      if (_T_288) begin
        reg_pc_1 <= _T_293;
      end
    end
    if (pc_valid) begin
      if (_T_278) begin
        reg_pred_0_redirect <= io_if_btb_0_redirect;
      end
    end
    if (pc_valid) begin
      if (_T_278) begin
        reg_pred_0_history <= io_if_btb_0_history;
      end
    end
    if (pc_valid) begin
      if (_T_278) begin
        reg_pred_0_diff <= io_if_btb_0_diff;
      end
    end
    if (pc_valid) begin
      if (_T_278) begin
        reg_pred_0_tgt <= io_if_btb_0_tgt;
      end
    end
    if (pc_valid) begin
      if (_T_288) begin
        reg_pred_1_redirect <= io_if_btb_1_redirect;
      end
    end
    if (pc_valid) begin
      if (_T_288) begin
        reg_pred_1_history <= io_if_btb_1_history;
      end
    end
    if (pc_valid) begin
      if (_T_288) begin
        reg_pred_1_diff <= io_if_btb_1_diff;
      end
    end
    if (pc_valid) begin
      if (_T_288) begin
        reg_pred_1_tgt <= io_if_btb_1_tgt;
      end
    end
    if (reset) begin
      _T_375 <= 32'h4033;
    end else begin
      if (inst_valid_0) begin
        _T_375 <= io_mem_inst_0_bits;
      end
    end
    if (reset) begin
      _T_378 <= 32'h4033;
    end else begin
      if (io_mem_inst_1_valid) begin
        _T_378 <= io_mem_inst_1_bits;
      end
    end
  end
endmodule
module MicroDecoder( // @[:@4189.2]
  input  [31:0] io_inst, // @[:@4192.4]
  output        io_is_bj, // @[:@4192.4]
  output        io_branch, // @[:@4192.4]
  output        io_call, // @[:@4192.4]
  output        io_retn // @[:@4192.4]
);
  wire [4:0] func; // @[MicroDecoder.scala 24:22:@4194.4]
  wire  jal; // @[MicroDecoder.scala 27:20:@4197.4]
  wire  jalr; // @[MicroDecoder.scala 28:20:@4198.4]
  wire  brnch; // @[MicroDecoder.scala 29:20:@4199.4]
  wire  _T_29; // @[MicroDecoder.scala 38:19:@4208.4]
  wire [4:0] rs1_addr; // @[MicroDecoder.scala 53:25:@4211.4]
  wire [4:0] wbaddr; // @[MicroDecoder.scala 54:25:@4212.4]
  wire  _T_32; // @[MicroDecoder.scala 39:37:@4213.4]
  wire  _T_34; // @[MicroDecoder.scala 39:53:@4214.4]
  wire  _T_35; // @[MicroDecoder.scala 39:45:@4215.4]
  wire  _T_36; // @[MicroDecoder.scala 55:23:@4216.4]
  wire  _T_38; // @[MicroDecoder.scala 39:37:@4217.4]
  wire  _T_40; // @[MicroDecoder.scala 39:53:@4218.4]
  wire  _T_41; // @[MicroDecoder.scala 39:45:@4219.4]
  wire  _T_42; // @[MicroDecoder.scala 55:39:@4220.4]
  wire  _T_43; // @[MicroDecoder.scala 55:67:@4221.4]
  wire  pop_push; // @[MicroDecoder.scala 55:57:@4222.4]
  wire  _T_49; // @[MicroDecoder.scala 71:20:@4226.4]
  wire  _T_62; // @[MicroDecoder.scala 72:31:@4234.4]
  wire  _T_63; // @[MicroDecoder.scala 72:28:@4235.4]
  wire  _T_64; // @[MicroDecoder.scala 71:39:@4236.4]
  wire  _T_77; // @[MicroDecoder.scala 73:58:@4245.4]
  wire  _T_78; // @[MicroDecoder.scala 73:48:@4246.4]
  wire  _T_79; // @[MicroDecoder.scala 72:48:@4247.4]
  wire  _T_87; // @[MicroDecoder.scala 75:23:@4253.4]
  wire  _T_88; // @[MicroDecoder.scala 75:20:@4254.4]
  wire  _T_94; // @[MicroDecoder.scala 75:37:@4258.4]
  assign func = io_inst[6:2]; // @[MicroDecoder.scala 24:22:@4194.4]
  assign jal = func == 5'h1b; // @[MicroDecoder.scala 27:20:@4197.4]
  assign jalr = func == 5'h19; // @[MicroDecoder.scala 28:20:@4198.4]
  assign brnch = func == 5'h18; // @[MicroDecoder.scala 29:20:@4199.4]
  assign _T_29 = jal | jalr; // @[MicroDecoder.scala 38:19:@4208.4]
  assign rs1_addr = io_inst[19:15]; // @[MicroDecoder.scala 53:25:@4211.4]
  assign wbaddr = io_inst[11:7]; // @[MicroDecoder.scala 54:25:@4212.4]
  assign _T_32 = wbaddr == 5'h1; // @[MicroDecoder.scala 39:37:@4213.4]
  assign _T_34 = wbaddr == 5'h5; // @[MicroDecoder.scala 39:53:@4214.4]
  assign _T_35 = _T_32 | _T_34; // @[MicroDecoder.scala 39:45:@4215.4]
  assign _T_36 = jalr & _T_35; // @[MicroDecoder.scala 55:23:@4216.4]
  assign _T_38 = rs1_addr == 5'h1; // @[MicroDecoder.scala 39:37:@4217.4]
  assign _T_40 = rs1_addr == 5'h5; // @[MicroDecoder.scala 39:53:@4218.4]
  assign _T_41 = _T_38 | _T_40; // @[MicroDecoder.scala 39:45:@4219.4]
  assign _T_42 = _T_36 & _T_41; // @[MicroDecoder.scala 55:39:@4220.4]
  assign _T_43 = wbaddr != rs1_addr; // @[MicroDecoder.scala 55:67:@4221.4]
  assign pop_push = _T_42 & _T_43; // @[MicroDecoder.scala 55:57:@4222.4]
  assign _T_49 = jal & _T_35; // @[MicroDecoder.scala 71:20:@4226.4]
  assign _T_62 = _T_41 == 1'h0; // @[MicroDecoder.scala 72:31:@4234.4]
  assign _T_63 = _T_36 & _T_62; // @[MicroDecoder.scala 72:28:@4235.4]
  assign _T_64 = _T_49 | _T_63; // @[MicroDecoder.scala 71:39:@4236.4]
  assign _T_77 = wbaddr == rs1_addr; // @[MicroDecoder.scala 73:58:@4245.4]
  assign _T_78 = _T_42 & _T_77; // @[MicroDecoder.scala 73:48:@4246.4]
  assign _T_79 = _T_64 | _T_78; // @[MicroDecoder.scala 72:48:@4247.4]
  assign _T_87 = _T_35 == 1'h0; // @[MicroDecoder.scala 75:23:@4253.4]
  assign _T_88 = jalr & _T_87; // @[MicroDecoder.scala 75:20:@4254.4]
  assign _T_94 = _T_88 & _T_41; // @[MicroDecoder.scala 75:37:@4258.4]
  assign io_is_bj = _T_29 | brnch; // @[MicroDecoder.scala 38:12:@4210.4]
  assign io_branch = func == 5'h18; // @[MicroDecoder.scala 37:13:@4207.4]
  assign io_call = _T_79 | pop_push; // @[MicroDecoder.scala 71:11:@4249.4]
  assign io_retn = _T_94 | pop_push; // @[MicroDecoder.scala 75:11:@4260.4]
endmodule
module FrontEnd( // @[:@4335.2]
  input         clock, // @[:@4336.4]
  input         reset, // @[:@4337.4]
  input  [31:0] io_cyc, // @[:@4338.4]
  input         io_mem_addr_ready, // @[:@4338.4]
  output        io_mem_addr_valid, // @[:@4338.4]
  output [31:0] io_mem_addr_bits, // @[:@4338.4]
  input         io_mem_inst_0_valid, // @[:@4338.4]
  input  [31:0] io_mem_inst_0_bits, // @[:@4338.4]
  input         io_mem_inst_1_valid, // @[:@4338.4]
  input  [31:0] io_mem_inst_1_bits, // @[:@4338.4]
  input         io_back_xcpt_valid, // @[:@4338.4]
  input  [31:0] io_back_xcpt_bits, // @[:@4338.4]
  input         io_back_kill, // @[:@4338.4]
  input         io_back_forward_0, // @[:@4338.4]
  input         io_back_forward_1, // @[:@4338.4]
  output        io_back_inst_0_valid, // @[:@4338.4]
  output [31:0] io_back_inst_0_bits, // @[:@4338.4]
  output        io_back_inst_1_valid, // @[:@4338.4]
  output [31:0] io_back_inst_1_bits, // @[:@4338.4]
  output [31:0] io_back_pc_0, // @[:@4338.4]
  output [31:0] io_back_pc_1, // @[:@4338.4]
  output        io_back_split, // @[:@4338.4]
  output        io_back_pred_redirect, // @[:@4338.4]
  output [9:0]  io_back_pred_history, // @[:@4338.4]
  output        io_back_pred_diff, // @[:@4338.4]
  output [31:0] io_back_pred_tgt, // @[:@4338.4]
  output        io_back_branch, // @[:@4338.4]
  output        io_back_call, // @[:@4338.4]
  output        io_back_retn, // @[:@4338.4]
  output        io_back_bj_sel_0, // @[:@4338.4]
  output        io_back_bj_sel_1, // @[:@4338.4]
  input         io_back_ras_pop, // @[:@4338.4]
  input         io_back_ras_push_valid, // @[:@4338.4]
  input  [31:0] io_back_ras_push_bits, // @[:@4338.4]
  input  [31:0] io_back_fb_pc, // @[:@4338.4]
  input  [1:0]  io_back_fb_type, // @[:@4338.4]
  input         io_back_feedBack_redirect, // @[:@4338.4]
  input  [9:0]  io_back_feedBack_history, // @[:@4338.4]
  input         io_back_feedBack_diff, // @[:@4338.4]
  input  [31:0] io_back_feedBack_tgt, // @[:@4338.4]
  input         io_back_feedBack_valid // @[:@4338.4]
);
  wire  BTB_clock; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_reset; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_if_pc_valid; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_if_pc_bits; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_predict_0_redirect; // @[FrontEnd.scala 12:24:@4340.4]
  wire [9:0] BTB_io_predict_0_history; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_predict_0_diff; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_predict_0_tgt; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_predict_1_redirect; // @[FrontEnd.scala 12:24:@4340.4]
  wire [9:0] BTB_io_predict_1_history; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_predict_1_diff; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_predict_1_tgt; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_split; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_branch; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_ras_pop; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_ras_push_valid; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_ras_push_bits; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_fb_pc_valid; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_fb_pc_bits; // @[FrontEnd.scala 12:24:@4340.4]
  wire [1:0] BTB_io_fb_type; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_feedBack_redirect; // @[FrontEnd.scala 12:24:@4340.4]
  wire [9:0] BTB_io_feedBack_history; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_feedBack_diff; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_feedBack_tgt; // @[FrontEnd.scala 12:24:@4340.4]
  wire  BTB_io_feedBack_valid; // @[FrontEnd.scala 12:24:@4340.4]
  wire [31:0] BTB_io_cyc; // @[FrontEnd.scala 12:24:@4340.4]
  wire  FetchInst_clock; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_reset; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_mem_addr_ready; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_mem_addr_valid; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_mem_addr_bits; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_mem_inst_0_valid; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_mem_inst_0_bits; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_mem_inst_1_valid; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_mem_inst_1_bits; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_if_btb_0_redirect; // @[FrontEnd.scala 13:24:@4343.4]
  wire [9:0] FetchInst_io_if_btb_0_history; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_if_btb_0_diff; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_if_btb_0_tgt; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_if_btb_1_redirect; // @[FrontEnd.scala 13:24:@4343.4]
  wire [9:0] FetchInst_io_if_btb_1_history; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_if_btb_1_diff; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_if_btb_1_tgt; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_dec_btb_0_redirect; // @[FrontEnd.scala 13:24:@4343.4]
  wire [9:0] FetchInst_io_dec_btb_0_history; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_dec_btb_0_diff; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_dec_btb_0_tgt; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_dec_btb_1_redirect; // @[FrontEnd.scala 13:24:@4343.4]
  wire [9:0] FetchInst_io_dec_btb_1_history; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_dec_btb_1_diff; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_dec_btb_1_tgt; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_pc; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_pc_split; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_pc_forward; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_forward_0; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_forward_1; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_if_kill; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_dec_kill; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_inst_0_valid; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_inst_0_bits; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_inst_1_valid; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_inst_1_bits; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_dec_pc_0; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] FetchInst_io_dec_pc_1; // @[FrontEnd.scala 13:24:@4343.4]
  wire  FetchInst_io_inst_split; // @[FrontEnd.scala 13:24:@4343.4]
  wire [31:0] MicroDecoder_io_inst; // @[FrontEnd.scala 14:38:@4346.4]
  wire  MicroDecoder_io_is_bj; // @[FrontEnd.scala 14:38:@4346.4]
  wire  MicroDecoder_io_branch; // @[FrontEnd.scala 14:38:@4346.4]
  wire  MicroDecoder_io_call; // @[FrontEnd.scala 14:38:@4346.4]
  wire  MicroDecoder_io_retn; // @[FrontEnd.scala 14:38:@4346.4]
  wire [31:0] MicroDecoder_1_io_inst; // @[FrontEnd.scala 14:38:@4349.4]
  wire  MicroDecoder_1_io_is_bj; // @[FrontEnd.scala 14:38:@4349.4]
  wire  MicroDecoder_1_io_branch; // @[FrontEnd.scala 14:38:@4349.4]
  wire  MicroDecoder_1_io_call; // @[FrontEnd.scala 14:38:@4349.4]
  wire  MicroDecoder_1_io_retn; // @[FrontEnd.scala 14:38:@4349.4]
  wire  dec_isbj_0; // @[FrontEnd.scala 15:60:@4352.4]
  wire  dec_isbj_1; // @[FrontEnd.scala 15:60:@4353.4]
  wire  _T_163; // @[FrontEnd.scala 16:62:@4354.4]
  wire  _T_164; // @[FrontEnd.scala 16:62:@4355.4]
  reg [31:0] if_reg_pc; // @[FrontEnd.scala 21:27:@4360.4]
  reg [31:0] _RAND_0;
  wire [32:0] _T_174; // @[FrontEnd.scala 26:50:@4361.4]
  wire [31:0] _T_175; // @[FrontEnd.scala 26:50:@4362.4]
  wire [31:0] _T_176; // @[FrontEnd.scala 27:12:@4363.4]
  wire  _T_199; // @[FrontEnd.scala 47:56:@4422.4]
  wire  _T_200; // @[FrontEnd.scala 47:53:@4423.4]
  wire  _T_201; // @[FrontEnd.scala 47:75:@4424.4]
  reg  _T_204; // @[BackEnd.scala 62:27:@4425.4]
  reg [31:0] _RAND_1;
  wire  dec_btb_error_1; // @[BackEnd.scala 65:8:@4433.4]
  wire [31:0] _T_177; // @[FrontEnd.scala 26:12:@4364.4]
  wire  _T_189; // @[FrontEnd.scala 47:56:@4408.4]
  wire  _T_190; // @[FrontEnd.scala 47:53:@4409.4]
  wire  _T_191; // @[FrontEnd.scala 47:75:@4410.4]
  reg  _T_194; // @[BackEnd.scala 62:27:@4411.4]
  reg [31:0] _RAND_2;
  wire  dec_btb_error_0; // @[BackEnd.scala 65:8:@4419.4]
  wire [31:0] _T_178; // @[FrontEnd.scala 25:12:@4365.4]
  wire [31:0] _T_179; // @[FrontEnd.scala 24:12:@4366.4]
  wire [31:0] if_next_pc; // @[FrontEnd.scala 23:12:@4367.4]
  wire [31:0] _GEN_0; // @[FrontEnd.scala 30:28:@4368.4]
  wire  _T_180; // @[FrontEnd.scala 36:35:@4388.4]
  wire  _T_181; // @[FrontEnd.scala 36:82:@4389.4]
  wire  _T_184; // @[FrontEnd.scala 39:64:@4395.4]
  wire  _T_186; // @[FrontEnd.scala 39:46:@4396.4]
  wire  _GEN_1; // @[BackEnd.scala 64:20:@4416.6]
  wire  _GEN_2; // @[BackEnd.scala 63:20:@4412.4]
  wire  _GEN_3; // @[BackEnd.scala 64:20:@4430.6]
  wire  _GEN_4; // @[BackEnd.scala 63:20:@4426.4]
  BTB BTB ( // @[FrontEnd.scala 12:24:@4340.4]
    .clock(BTB_clock),
    .reset(BTB_reset),
    .io_if_pc_valid(BTB_io_if_pc_valid),
    .io_if_pc_bits(BTB_io_if_pc_bits),
    .io_predict_0_redirect(BTB_io_predict_0_redirect),
    .io_predict_0_history(BTB_io_predict_0_history),
    .io_predict_0_diff(BTB_io_predict_0_diff),
    .io_predict_0_tgt(BTB_io_predict_0_tgt),
    .io_predict_1_redirect(BTB_io_predict_1_redirect),
    .io_predict_1_history(BTB_io_predict_1_history),
    .io_predict_1_diff(BTB_io_predict_1_diff),
    .io_predict_1_tgt(BTB_io_predict_1_tgt),
    .io_split(BTB_io_split),
    .io_branch(BTB_io_branch),
    .io_ras_pop(BTB_io_ras_pop),
    .io_ras_push_valid(BTB_io_ras_push_valid),
    .io_ras_push_bits(BTB_io_ras_push_bits),
    .io_fb_pc_valid(BTB_io_fb_pc_valid),
    .io_fb_pc_bits(BTB_io_fb_pc_bits),
    .io_fb_type(BTB_io_fb_type),
    .io_feedBack_redirect(BTB_io_feedBack_redirect),
    .io_feedBack_history(BTB_io_feedBack_history),
    .io_feedBack_diff(BTB_io_feedBack_diff),
    .io_feedBack_tgt(BTB_io_feedBack_tgt),
    .io_feedBack_valid(BTB_io_feedBack_valid),
    .io_cyc(BTB_io_cyc)
  );
  FetchInst FetchInst ( // @[FrontEnd.scala 13:24:@4343.4]
    .clock(FetchInst_clock),
    .reset(FetchInst_reset),
    .io_mem_addr_ready(FetchInst_io_mem_addr_ready),
    .io_mem_addr_valid(FetchInst_io_mem_addr_valid),
    .io_mem_addr_bits(FetchInst_io_mem_addr_bits),
    .io_mem_inst_0_valid(FetchInst_io_mem_inst_0_valid),
    .io_mem_inst_0_bits(FetchInst_io_mem_inst_0_bits),
    .io_mem_inst_1_valid(FetchInst_io_mem_inst_1_valid),
    .io_mem_inst_1_bits(FetchInst_io_mem_inst_1_bits),
    .io_if_btb_0_redirect(FetchInst_io_if_btb_0_redirect),
    .io_if_btb_0_history(FetchInst_io_if_btb_0_history),
    .io_if_btb_0_diff(FetchInst_io_if_btb_0_diff),
    .io_if_btb_0_tgt(FetchInst_io_if_btb_0_tgt),
    .io_if_btb_1_redirect(FetchInst_io_if_btb_1_redirect),
    .io_if_btb_1_history(FetchInst_io_if_btb_1_history),
    .io_if_btb_1_diff(FetchInst_io_if_btb_1_diff),
    .io_if_btb_1_tgt(FetchInst_io_if_btb_1_tgt),
    .io_dec_btb_0_redirect(FetchInst_io_dec_btb_0_redirect),
    .io_dec_btb_0_history(FetchInst_io_dec_btb_0_history),
    .io_dec_btb_0_diff(FetchInst_io_dec_btb_0_diff),
    .io_dec_btb_0_tgt(FetchInst_io_dec_btb_0_tgt),
    .io_dec_btb_1_redirect(FetchInst_io_dec_btb_1_redirect),
    .io_dec_btb_1_history(FetchInst_io_dec_btb_1_history),
    .io_dec_btb_1_diff(FetchInst_io_dec_btb_1_diff),
    .io_dec_btb_1_tgt(FetchInst_io_dec_btb_1_tgt),
    .io_pc(FetchInst_io_pc),
    .io_pc_split(FetchInst_io_pc_split),
    .io_pc_forward(FetchInst_io_pc_forward),
    .io_forward_0(FetchInst_io_forward_0),
    .io_forward_1(FetchInst_io_forward_1),
    .io_if_kill(FetchInst_io_if_kill),
    .io_dec_kill(FetchInst_io_dec_kill),
    .io_inst_0_valid(FetchInst_io_inst_0_valid),
    .io_inst_0_bits(FetchInst_io_inst_0_bits),
    .io_inst_1_valid(FetchInst_io_inst_1_valid),
    .io_inst_1_bits(FetchInst_io_inst_1_bits),
    .io_dec_pc_0(FetchInst_io_dec_pc_0),
    .io_dec_pc_1(FetchInst_io_dec_pc_1),
    .io_inst_split(FetchInst_io_inst_split)
  );
  MicroDecoder MicroDecoder ( // @[FrontEnd.scala 14:38:@4346.4]
    .io_inst(MicroDecoder_io_inst),
    .io_is_bj(MicroDecoder_io_is_bj),
    .io_branch(MicroDecoder_io_branch),
    .io_call(MicroDecoder_io_call),
    .io_retn(MicroDecoder_io_retn)
  );
  MicroDecoder MicroDecoder_1 ( // @[FrontEnd.scala 14:38:@4349.4]
    .io_inst(MicroDecoder_1_io_inst),
    .io_is_bj(MicroDecoder_1_io_is_bj),
    .io_branch(MicroDecoder_1_io_branch),
    .io_call(MicroDecoder_1_io_call),
    .io_retn(MicroDecoder_1_io_retn)
  );
  assign dec_isbj_0 = FetchInst_io_inst_0_valid & MicroDecoder_io_is_bj; // @[FrontEnd.scala 15:60:@4352.4]
  assign dec_isbj_1 = FetchInst_io_inst_1_valid & MicroDecoder_1_io_is_bj; // @[FrontEnd.scala 15:60:@4353.4]
  assign _T_163 = FetchInst_io_inst_0_valid & MicroDecoder_io_branch; // @[FrontEnd.scala 16:62:@4354.4]
  assign _T_164 = FetchInst_io_inst_1_valid & MicroDecoder_1_io_branch; // @[FrontEnd.scala 16:62:@4355.4]
  assign _T_174 = FetchInst_io_dec_pc_1 + 32'h4; // @[FrontEnd.scala 26:50:@4361.4]
  assign _T_175 = FetchInst_io_dec_pc_1 + 32'h4; // @[FrontEnd.scala 26:50:@4362.4]
  assign _T_176 = BTB_io_split ? BTB_io_predict_0_tgt : BTB_io_predict_1_tgt; // @[FrontEnd.scala 27:12:@4363.4]
  assign _T_199 = MicroDecoder_1_io_is_bj == 1'h0; // @[FrontEnd.scala 47:56:@4422.4]
  assign _T_200 = FetchInst_io_inst_1_valid & _T_199; // @[FrontEnd.scala 47:53:@4423.4]
  assign _T_201 = _T_200 & FetchInst_io_dec_btb_1_redirect; // @[FrontEnd.scala 47:75:@4424.4]
  assign dec_btb_error_1 = _T_201 & _T_204; // @[BackEnd.scala 65:8:@4433.4]
  assign _T_177 = dec_btb_error_1 ? _T_175 : _T_176; // @[FrontEnd.scala 26:12:@4364.4]
  assign _T_189 = MicroDecoder_io_is_bj == 1'h0; // @[FrontEnd.scala 47:56:@4408.4]
  assign _T_190 = FetchInst_io_inst_0_valid & _T_189; // @[FrontEnd.scala 47:53:@4409.4]
  assign _T_191 = _T_190 & FetchInst_io_dec_btb_0_redirect; // @[FrontEnd.scala 47:75:@4410.4]
  assign dec_btb_error_0 = _T_191 & _T_194; // @[BackEnd.scala 65:8:@4419.4]
  assign _T_178 = dec_btb_error_0 ? FetchInst_io_dec_pc_1 : _T_177; // @[FrontEnd.scala 25:12:@4365.4]
  assign _T_179 = io_back_kill ? io_back_feedBack_tgt : _T_178; // @[FrontEnd.scala 24:12:@4366.4]
  assign if_next_pc = io_back_xcpt_valid ? io_back_xcpt_bits : _T_179; // @[FrontEnd.scala 23:12:@4367.4]
  assign _GEN_0 = FetchInst_io_pc_forward ? if_next_pc : if_reg_pc; // @[FrontEnd.scala 30:28:@4368.4]
  assign _T_180 = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 36:35:@4388.4]
  assign _T_181 = dec_btb_error_0 | dec_btb_error_1; // @[FrontEnd.scala 36:82:@4389.4]
  assign _T_184 = dec_isbj_0 & dec_isbj_1; // @[FrontEnd.scala 39:64:@4395.4]
  assign _T_186 = _T_184 == 1'h0; // @[FrontEnd.scala 39:46:@4396.4]
  assign _GEN_1 = _T_191 ? 1'h0 : _T_194; // @[BackEnd.scala 64:20:@4416.6]
  assign _GEN_2 = io_back_forward_0 ? 1'h1 : _GEN_1; // @[BackEnd.scala 63:20:@4412.4]
  assign _GEN_3 = _T_201 ? 1'h0 : _T_204; // @[BackEnd.scala 64:20:@4430.6]
  assign _GEN_4 = io_back_forward_1 ? 1'h1 : _GEN_3; // @[BackEnd.scala 63:20:@4426.4]
  assign io_mem_addr_valid = FetchInst_io_mem_addr_valid; // @[FrontEnd.scala 32:19:@4376.4]
  assign io_mem_addr_bits = FetchInst_io_mem_addr_bits; // @[FrontEnd.scala 32:19:@4375.4]
  assign io_back_inst_0_valid = FetchInst_io_inst_0_valid; // @[FrontEnd.scala 42:17:@4403.4]
  assign io_back_inst_0_bits = FetchInst_io_inst_0_bits; // @[FrontEnd.scala 42:17:@4402.4]
  assign io_back_inst_1_valid = FetchInst_io_inst_1_valid; // @[FrontEnd.scala 42:17:@4405.4]
  assign io_back_inst_1_bits = FetchInst_io_inst_1_bits; // @[FrontEnd.scala 42:17:@4404.4]
  assign io_back_pc_0 = FetchInst_io_dec_pc_0; // @[FrontEnd.scala 41:17:@4400.4]
  assign io_back_pc_1 = FetchInst_io_dec_pc_1; // @[FrontEnd.scala 41:17:@4401.4]
  assign io_back_split = _T_191 & _T_194; // @[FrontEnd.scala 43:17:@4406.4]
  assign io_back_pred_redirect = dec_isbj_0 ? FetchInst_io_dec_btb_0_redirect : FetchInst_io_dec_btb_1_redirect; // @[FrontEnd.scala 54:18:@4447.4]
  assign io_back_pred_history = dec_isbj_0 ? FetchInst_io_dec_btb_0_history : FetchInst_io_dec_btb_1_history; // @[FrontEnd.scala 54:18:@4446.4]
  assign io_back_pred_diff = dec_isbj_0 ? FetchInst_io_dec_btb_0_diff : FetchInst_io_dec_btb_1_diff; // @[FrontEnd.scala 54:18:@4445.4]
  assign io_back_pred_tgt = dec_isbj_0 ? FetchInst_io_dec_btb_0_tgt : FetchInst_io_dec_btb_1_tgt; // @[FrontEnd.scala 54:18:@4444.4]
  assign io_back_branch = dec_isbj_0 ? MicroDecoder_io_branch : MicroDecoder_1_io_branch; // @[FrontEnd.scala 51:18:@4438.4]
  assign io_back_call = dec_isbj_0 ? MicroDecoder_io_call : MicroDecoder_1_io_call; // @[FrontEnd.scala 52:18:@4440.4]
  assign io_back_retn = dec_isbj_0 ? MicroDecoder_io_retn : MicroDecoder_1_io_retn; // @[FrontEnd.scala 53:18:@4442.4]
  assign io_back_bj_sel_0 = MicroDecoder_io_is_bj; // @[FrontEnd.scala 50:18:@4435.4]
  assign io_back_bj_sel_1 = MicroDecoder_1_io_is_bj; // @[FrontEnd.scala 50:18:@4436.4]
  assign BTB_clock = clock; // @[:@4341.4]
  assign BTB_reset = reset; // @[:@4342.4]
  assign BTB_io_if_pc_valid = FetchInst_io_pc_forward; // @[FrontEnd.scala 56:19:@4448.4]
  assign BTB_io_if_pc_bits = if_reg_pc; // @[FrontEnd.scala 57:19:@4449.4]
  assign BTB_io_branch = _T_163 | _T_164; // @[FrontEnd.scala 61:16:@4452.4]
  assign BTB_io_ras_pop = io_back_ras_pop; // @[FrontEnd.scala 66:16:@4461.4]
  assign BTB_io_ras_push_valid = io_back_ras_push_valid; // @[FrontEnd.scala 65:16:@4460.4]
  assign BTB_io_ras_push_bits = io_back_ras_push_bits; // @[FrontEnd.scala 65:16:@4459.4]
  assign BTB_io_fb_pc_valid = io_back_kill; // @[FrontEnd.scala 58:19:@4450.4]
  assign BTB_io_fb_pc_bits = io_back_fb_pc; // @[FrontEnd.scala 59:19:@4451.4]
  assign BTB_io_fb_type = io_back_fb_type; // @[FrontEnd.scala 63:16:@4453.4]
  assign BTB_io_feedBack_redirect = io_back_feedBack_redirect; // @[FrontEnd.scala 64:16:@4458.4]
  assign BTB_io_feedBack_history = io_back_feedBack_history; // @[FrontEnd.scala 64:16:@4457.4]
  assign BTB_io_feedBack_diff = io_back_feedBack_diff; // @[FrontEnd.scala 64:16:@4456.4]
  assign BTB_io_feedBack_tgt = io_back_feedBack_tgt; // @[FrontEnd.scala 64:16:@4455.4]
  assign BTB_io_feedBack_valid = io_back_feedBack_valid; // @[FrontEnd.scala 64:16:@4454.4]
  assign BTB_io_cyc = io_cyc; // @[FrontEnd.scala 17:14:@4357.4]
  assign FetchInst_clock = clock; // @[:@4344.4]
  assign FetchInst_reset = reset; // @[:@4345.4]
  assign FetchInst_io_mem_addr_ready = io_mem_addr_ready; // @[FrontEnd.scala 32:19:@4377.4]
  assign FetchInst_io_mem_inst_0_valid = io_mem_inst_0_valid; // @[FrontEnd.scala 32:19:@4372.4]
  assign FetchInst_io_mem_inst_0_bits = io_mem_inst_0_bits; // @[FrontEnd.scala 32:19:@4371.4]
  assign FetchInst_io_mem_inst_1_valid = io_mem_inst_1_valid; // @[FrontEnd.scala 32:19:@4374.4]
  assign FetchInst_io_mem_inst_1_bits = io_mem_inst_1_bits; // @[FrontEnd.scala 32:19:@4373.4]
  assign FetchInst_io_if_btb_0_redirect = BTB_io_predict_0_redirect; // @[FrontEnd.scala 35:19:@4383.4]
  assign FetchInst_io_if_btb_0_history = BTB_io_predict_0_history; // @[FrontEnd.scala 35:19:@4382.4]
  assign FetchInst_io_if_btb_0_diff = BTB_io_predict_0_diff; // @[FrontEnd.scala 35:19:@4381.4]
  assign FetchInst_io_if_btb_0_tgt = BTB_io_predict_0_tgt; // @[FrontEnd.scala 35:19:@4380.4]
  assign FetchInst_io_if_btb_1_redirect = BTB_io_predict_1_redirect; // @[FrontEnd.scala 35:19:@4387.4]
  assign FetchInst_io_if_btb_1_history = BTB_io_predict_1_history; // @[FrontEnd.scala 35:19:@4386.4]
  assign FetchInst_io_if_btb_1_diff = BTB_io_predict_1_diff; // @[FrontEnd.scala 35:19:@4385.4]
  assign FetchInst_io_if_btb_1_tgt = BTB_io_predict_1_tgt; // @[FrontEnd.scala 35:19:@4384.4]
  assign FetchInst_io_pc = if_reg_pc; // @[FrontEnd.scala 33:19:@4378.4]
  assign FetchInst_io_pc_split = BTB_io_split; // @[FrontEnd.scala 34:19:@4379.4]
  assign FetchInst_io_forward_0 = io_back_forward_0; // @[FrontEnd.scala 38:21:@4394.4]
  assign FetchInst_io_forward_1 = io_back_forward_1 & _T_186; // @[FrontEnd.scala 39:21:@4398.4]
  assign FetchInst_io_if_kill = _T_180 | _T_181; // @[FrontEnd.scala 36:19:@4391.4]
  assign FetchInst_io_dec_kill = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 37:19:@4393.4]
  assign FetchInst_io_inst_split = _T_191 & _T_194; // @[FrontEnd.scala 40:21:@4399.4]
  assign MicroDecoder_io_inst = FetchInst_io_inst_0_bits; // @[FrontEnd.scala 46:23:@4407.4]
  assign MicroDecoder_1_io_inst = FetchInst_io_inst_1_bits; // @[FrontEnd.scala 46:23:@4421.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_reg_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  _T_204 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  _T_194 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      if_reg_pc <= 32'h80000000;
    end else begin
      if (FetchInst_io_pc_forward) begin
        if (io_back_xcpt_valid) begin
          if_reg_pc <= io_back_xcpt_bits;
        end else begin
          if (io_back_kill) begin
            if_reg_pc <= io_back_feedBack_tgt;
          end else begin
            if (dec_btb_error_0) begin
              if_reg_pc <= FetchInst_io_dec_pc_1;
            end else begin
              if (dec_btb_error_1) begin
                if_reg_pc <= _T_175;
              end else begin
                if (BTB_io_split) begin
                  if_reg_pc <= BTB_io_predict_0_tgt;
                end else begin
                  if_reg_pc <= BTB_io_predict_1_tgt;
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      _T_204 <= 1'h1;
    end else begin
      if (io_back_forward_1) begin
        _T_204 <= 1'h1;
      end else begin
        if (_T_201) begin
          _T_204 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_194 <= 1'h1;
    end else begin
      if (io_back_forward_0) begin
        _T_194 <= 1'h1;
      end else begin
        if (_T_191) begin
          _T_194 <= 1'h0;
        end
      end
    end
  end
endmodule
module CSRFile( // @[:@4463.2]
  input         clock, // @[:@4464.4]
  input         reset, // @[:@4465.4]
  input  [2:0]  io_rw_cmd, // @[:@4466.4]
  input  [11:0] io_rw_addr, // @[:@4466.4]
  output [31:0] io_rw_rdata, // @[:@4466.4]
  input  [31:0] io_rw_wdata, // @[:@4466.4]
  output        io_eret, // @[:@4466.4]
  output [1:0]  io_status_prv, // @[:@4466.4]
  output [13:0] io_status_unimp5, // @[:@4466.4]
  output        io_status_mprv, // @[:@4466.4]
  output [1:0]  io_status_unimp4, // @[:@4466.4]
  output [1:0]  io_status_mpp, // @[:@4466.4]
  output [2:0]  io_status_unimp3, // @[:@4466.4]
  output        io_status_mpie, // @[:@4466.4]
  output [2:0]  io_status_unimp2, // @[:@4466.4]
  output        io_status_mie, // @[:@4466.4]
  output [2:0]  io_status_unimp1, // @[:@4466.4]
  input         io_xcpt, // @[:@4466.4]
  input  [31:0] io_cause, // @[:@4466.4]
  input  [31:0] io_tval, // @[:@4466.4]
  output [31:0] io_evec, // @[:@4466.4]
  input         io_illegal, // @[:@4466.4]
  input  [1:0]  io_retire, // @[:@4466.4]
  input  [31:0] io_pc, // @[:@4466.4]
  output [31:0] io_time // @[:@4466.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 112:28:@4593.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 112:28:@4593.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 112:28:@4593.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[CSR.scala 113:21:@4594.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[CSR.scala 114:23:@4595.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[CSR.scala 115:22:@4596.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[CSR.scala 116:25:@4597.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[CSR.scala 118:24:@4599.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[CSR.scala 120:24:@4617.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[CSR.scala 120:24:@4617.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[CSR.scala 121:24:@4635.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[CSR.scala 121:24:@4635.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_240; // @[Util.scala 112:41:@4638.4]
  reg [31:0] _RAND_12;
  wire [6:0] _T_241; // @[Util.scala 113:33:@4639.4]
  reg [57:0] _T_244; // @[Util.scala 117:31:@4641.4]
  reg [63:0] _RAND_13;
  wire  _T_245; // @[Util.scala 118:20:@4642.4]
  wire [58:0] _T_247; // @[Util.scala 118:43:@4644.6]
  wire [57:0] _T_248; // @[Util.scala 118:43:@4645.6]
  wire [57:0] _GEN_0; // @[Util.scala 118:34:@4643.4]
  wire [63:0] _T_249; // @[Cat.scala 30:58:@4648.4]
  reg [5:0] _T_252; // @[Util.scala 112:41:@4649.4]
  reg [31:0] _RAND_14;
  wire [5:0] _GEN_147; // @[Util.scala 113:33:@4650.4]
  wire [6:0] _T_253; // @[Util.scala 113:33:@4650.4]
  reg [57:0] _T_256; // @[Util.scala 117:31:@4652.4]
  reg [63:0] _RAND_15;
  wire  _T_257; // @[Util.scala 118:20:@4653.4]
  wire [58:0] _T_259; // @[Util.scala 118:43:@4655.6]
  wire [57:0] _T_260; // @[Util.scala 118:43:@4656.6]
  wire [57:0] _GEN_1; // @[Util.scala 118:34:@4654.4]
  wire [63:0] _T_261; // @[Cat.scala 30:58:@4659.4]
  reg [39:0] _T_264; // @[Util.scala 112:74:@4661.4]
  reg [63:0] _RAND_16;
  wire [40:0] _T_265; // @[Util.scala 113:33:@4662.4]
  reg [39:0] _T_267; // @[Util.scala 112:74:@4664.4]
  reg [63:0] _RAND_17;
  wire [40:0] _T_268; // @[Util.scala 113:33:@4665.4]
  reg [39:0] _T_270; // @[Util.scala 112:74:@4667.4]
  reg [63:0] _RAND_18;
  wire [40:0] _T_271; // @[Util.scala 113:33:@4668.4]
  reg [39:0] _T_273; // @[Util.scala 112:74:@4670.4]
  reg [63:0] _RAND_19;
  wire [40:0] _T_274; // @[Util.scala 113:33:@4671.4]
  reg [39:0] _T_276; // @[Util.scala 112:74:@4673.4]
  reg [63:0] _RAND_20;
  wire [40:0] _T_277; // @[Util.scala 113:33:@4674.4]
  reg [39:0] _T_279; // @[Util.scala 112:74:@4676.4]
  reg [63:0] _RAND_21;
  wire [40:0] _T_280; // @[Util.scala 113:33:@4677.4]
  reg [39:0] _T_282; // @[Util.scala 112:74:@4679.4]
  reg [63:0] _RAND_22;
  wire [40:0] _T_283; // @[Util.scala 113:33:@4680.4]
  reg [39:0] _T_285; // @[Util.scala 112:74:@4682.4]
  reg [63:0] _RAND_23;
  wire [40:0] _T_286; // @[Util.scala 113:33:@4683.4]
  reg [39:0] _T_288; // @[Util.scala 112:74:@4685.4]
  reg [63:0] _RAND_24;
  wire [40:0] _T_289; // @[Util.scala 113:33:@4686.4]
  reg [39:0] _T_291; // @[Util.scala 112:74:@4688.4]
  reg [63:0] _RAND_25;
  wire [40:0] _T_292; // @[Util.scala 113:33:@4689.4]
  reg [39:0] _T_294; // @[Util.scala 112:74:@4691.4]
  reg [63:0] _RAND_26;
  wire [40:0] _T_295; // @[Util.scala 113:33:@4692.4]
  reg [39:0] _T_297; // @[Util.scala 112:74:@4694.4]
  reg [63:0] _RAND_27;
  wire [40:0] _T_298; // @[Util.scala 113:33:@4695.4]
  reg [39:0] _T_300; // @[Util.scala 112:74:@4697.4]
  reg [63:0] _RAND_28;
  wire [40:0] _T_301; // @[Util.scala 113:33:@4698.4]
  reg [39:0] _T_303; // @[Util.scala 112:74:@4700.4]
  reg [63:0] _RAND_29;
  wire [40:0] _T_304; // @[Util.scala 113:33:@4701.4]
  reg [39:0] _T_306; // @[Util.scala 112:74:@4703.4]
  reg [63:0] _RAND_30;
  wire [40:0] _T_307; // @[Util.scala 113:33:@4704.4]
  reg [39:0] _T_309; // @[Util.scala 112:74:@4706.4]
  reg [63:0] _RAND_31;
  wire [40:0] _T_310; // @[Util.scala 113:33:@4707.4]
  reg [39:0] _T_312; // @[Util.scala 112:74:@4709.4]
  reg [63:0] _RAND_32;
  wire [40:0] _T_313; // @[Util.scala 113:33:@4710.4]
  reg [39:0] _T_315; // @[Util.scala 112:74:@4712.4]
  reg [63:0] _RAND_33;
  wire [40:0] _T_316; // @[Util.scala 113:33:@4713.4]
  reg [39:0] _T_318; // @[Util.scala 112:74:@4715.4]
  reg [63:0] _RAND_34;
  wire [40:0] _T_319; // @[Util.scala 113:33:@4716.4]
  reg [39:0] _T_321; // @[Util.scala 112:74:@4718.4]
  reg [63:0] _RAND_35;
  wire [40:0] _T_322; // @[Util.scala 113:33:@4719.4]
  reg [39:0] _T_324; // @[Util.scala 112:74:@4721.4]
  reg [63:0] _RAND_36;
  wire [40:0] _T_325; // @[Util.scala 113:33:@4722.4]
  reg [39:0] _T_327; // @[Util.scala 112:74:@4724.4]
  reg [63:0] _RAND_37;
  wire [40:0] _T_328; // @[Util.scala 113:33:@4725.4]
  reg [39:0] _T_330; // @[Util.scala 112:74:@4727.4]
  reg [63:0] _RAND_38;
  wire [40:0] _T_331; // @[Util.scala 113:33:@4728.4]
  reg [39:0] _T_333; // @[Util.scala 112:74:@4730.4]
  reg [63:0] _RAND_39;
  wire [40:0] _T_334; // @[Util.scala 113:33:@4731.4]
  reg [39:0] _T_336; // @[Util.scala 112:74:@4733.4]
  reg [63:0] _RAND_40;
  wire [40:0] _T_337; // @[Util.scala 113:33:@4734.4]
  reg [39:0] _T_339; // @[Util.scala 112:74:@4736.4]
  reg [63:0] _RAND_41;
  wire [40:0] _T_340; // @[Util.scala 113:33:@4737.4]
  reg [39:0] _T_342; // @[Util.scala 112:74:@4739.4]
  reg [63:0] _RAND_42;
  wire [40:0] _T_343; // @[Util.scala 113:33:@4740.4]
  reg [39:0] _T_345; // @[Util.scala 112:74:@4742.4]
  reg [63:0] _RAND_43;
  wire [40:0] _T_346; // @[Util.scala 113:33:@4743.4]
  reg [39:0] _T_348; // @[Util.scala 112:74:@4745.4]
  reg [63:0] _RAND_44;
  wire [40:0] _T_349; // @[Util.scala 113:33:@4746.4]
  reg [39:0] _T_351; // @[Util.scala 112:74:@4748.4]
  reg [63:0] _RAND_45;
  wire [40:0] _T_352; // @[Util.scala 113:33:@4749.4]
  reg [39:0] _T_354; // @[Util.scala 112:74:@4751.4]
  reg [63:0] _RAND_46;
  wire [40:0] _T_355; // @[Util.scala 113:33:@4752.4]
  reg [39:0] _T_357; // @[Util.scala 112:74:@4754.4]
  reg [63:0] _RAND_47;
  wire [40:0] _T_358; // @[Util.scala 113:33:@4755.4]
  reg [31:0] reg_dscratch; // @[CSR.scala 134:25:@4844.4]
  reg [31:0] _RAND_48;
  wire  system_insn; // @[CSR.scala 137:31:@4846.4]
  wire  _T_446; // @[CSR.scala 138:27:@4847.4]
  wire  _T_448; // @[CSR.scala 138:40:@4848.4]
  wire  cpu_ren; // @[CSR.scala 138:37:@4849.4]
  wire [31:0] read_mstatus; // @[CSR.scala 140:32:@4858.4]
  wire [15:0] _T_468; // @[CSR.scala 156:25:@4864.4]
  wire [15:0] _T_474; // @[CSR.scala 157:25:@4870.4]
  wire  _T_478; // @[CSR.scala 177:73:@4871.4]
  wire  _T_480; // @[CSR.scala 177:73:@4872.4]
  wire  _T_482; // @[CSR.scala 177:73:@4873.4]
  wire  _T_488; // @[CSR.scala 177:73:@4876.4]
  wire  _T_490; // @[CSR.scala 177:73:@4877.4]
  wire  _T_492; // @[CSR.scala 177:73:@4878.4]
  wire  _T_494; // @[CSR.scala 177:73:@4879.4]
  wire  _T_496; // @[CSR.scala 177:73:@4880.4]
  wire  _T_498; // @[CSR.scala 177:73:@4881.4]
  wire  _T_500; // @[CSR.scala 177:73:@4882.4]
  wire  _T_502; // @[CSR.scala 177:73:@4883.4]
  wire  _T_504; // @[CSR.scala 177:73:@4884.4]
  wire  _T_508; // @[CSR.scala 177:73:@4886.4]
  wire  _T_510; // @[CSR.scala 177:73:@4887.4]
  wire  _T_512; // @[CSR.scala 177:73:@4888.4]
  wire  _T_514; // @[CSR.scala 177:73:@4889.4]
  wire  _T_516; // @[CSR.scala 177:73:@4890.4]
  wire  _T_518; // @[CSR.scala 177:73:@4891.4]
  wire  _T_520; // @[CSR.scala 177:73:@4892.4]
  wire  _T_522; // @[CSR.scala 177:73:@4893.4]
  wire  _T_524; // @[CSR.scala 177:73:@4894.4]
  wire  _T_526; // @[CSR.scala 177:73:@4895.4]
  wire  _T_528; // @[CSR.scala 177:73:@4896.4]
  wire  _T_530; // @[CSR.scala 177:73:@4897.4]
  wire  _T_532; // @[CSR.scala 177:73:@4898.4]
  wire  _T_534; // @[CSR.scala 177:73:@4899.4]
  wire  _T_536; // @[CSR.scala 177:73:@4900.4]
  wire  _T_538; // @[CSR.scala 177:73:@4901.4]
  wire  _T_540; // @[CSR.scala 177:73:@4902.4]
  wire  _T_542; // @[CSR.scala 177:73:@4903.4]
  wire  _T_544; // @[CSR.scala 177:73:@4904.4]
  wire  _T_546; // @[CSR.scala 177:73:@4905.4]
  wire  _T_548; // @[CSR.scala 177:73:@4906.4]
  wire  _T_550; // @[CSR.scala 177:73:@4907.4]
  wire  _T_552; // @[CSR.scala 177:73:@4908.4]
  wire  _T_554; // @[CSR.scala 177:73:@4909.4]
  wire  _T_556; // @[CSR.scala 177:73:@4910.4]
  wire  _T_558; // @[CSR.scala 177:73:@4911.4]
  wire  _T_560; // @[CSR.scala 177:73:@4912.4]
  wire  _T_562; // @[CSR.scala 177:73:@4913.4]
  wire  _T_564; // @[CSR.scala 177:73:@4914.4]
  wire  _T_566; // @[CSR.scala 177:73:@4915.4]
  wire  _T_568; // @[CSR.scala 177:73:@4916.4]
  wire  _T_570; // @[CSR.scala 177:73:@4917.4]
  wire  _T_572; // @[CSR.scala 177:73:@4918.4]
  wire  _T_574; // @[CSR.scala 177:73:@4919.4]
  wire  _T_576; // @[CSR.scala 177:73:@4920.4]
  wire  _T_578; // @[CSR.scala 177:73:@4921.4]
  wire  _T_580; // @[CSR.scala 177:73:@4922.4]
  wire  _T_582; // @[CSR.scala 177:73:@4923.4]
  wire  _T_584; // @[CSR.scala 177:73:@4924.4]
  wire  _T_586; // @[CSR.scala 177:73:@4925.4]
  wire  _T_588; // @[CSR.scala 177:73:@4926.4]
  wire  _T_590; // @[CSR.scala 177:73:@4927.4]
  wire  _T_592; // @[CSR.scala 177:73:@4928.4]
  wire  _T_594; // @[CSR.scala 177:73:@4929.4]
  wire  _T_596; // @[CSR.scala 177:73:@4930.4]
  wire  _T_598; // @[CSR.scala 177:73:@4931.4]
  wire  _T_600; // @[CSR.scala 177:73:@4932.4]
  wire  _T_602; // @[CSR.scala 177:73:@4933.4]
  wire  _T_604; // @[CSR.scala 177:73:@4934.4]
  wire  _T_606; // @[CSR.scala 177:73:@4935.4]
  wire  _T_608; // @[CSR.scala 177:73:@4936.4]
  wire  _T_610; // @[CSR.scala 177:73:@4937.4]
  wire  _T_612; // @[CSR.scala 177:73:@4938.4]
  wire  _T_614; // @[CSR.scala 177:73:@4939.4]
  wire  _T_616; // @[CSR.scala 177:73:@4940.4]
  wire  _T_618; // @[CSR.scala 177:73:@4941.4]
  wire  _T_620; // @[CSR.scala 177:73:@4942.4]
  wire  _T_622; // @[CSR.scala 177:73:@4943.4]
  wire  _T_624; // @[CSR.scala 177:73:@4944.4]
  wire  _T_626; // @[CSR.scala 177:73:@4945.4]
  wire  _T_628; // @[CSR.scala 177:73:@4946.4]
  wire  _T_630; // @[CSR.scala 177:73:@4947.4]
  wire  _T_632; // @[CSR.scala 177:73:@4948.4]
  wire  _T_634; // @[CSR.scala 177:73:@4949.4]
  wire  _T_636; // @[CSR.scala 177:73:@4950.4]
  wire  _T_638; // @[CSR.scala 177:73:@4951.4]
  wire  _T_640; // @[CSR.scala 177:73:@4952.4]
  wire  _T_642; // @[CSR.scala 177:73:@4953.4]
  wire [1:0] _T_643; // @[CSR.scala 179:54:@4954.4]
  wire  priv_sufficient; // @[CSR.scala 179:41:@4955.4]
  wire [1:0] _T_644; // @[CSR.scala 180:29:@4956.4]
  wire [1:0] _T_645; // @[CSR.scala 180:37:@4957.4]
  wire  read_only; // @[CSR.scala 180:37:@4958.4]
  wire  _T_647; // @[CSR.scala 181:38:@4959.4]
  wire  _T_648; // @[CSR.scala 181:25:@4960.4]
  wire  cpu_wen; // @[CSR.scala 181:48:@4961.4]
  wire  _T_650; // @[CSR.scala 182:24:@4962.4]
  wire  wen; // @[CSR.scala 182:21:@4963.4]
  wire  _T_651; // @[Util.scala 23:47:@4964.4]
  wire  _T_652; // @[Util.scala 23:47:@4965.4]
  wire  _T_653; // @[Util.scala 23:62:@4966.4]
  wire [31:0] _T_655; // @[CSR.scala 281:9:@4967.4]
  wire [31:0] _T_656; // @[CSR.scala 281:49:@4968.4]
  wire [31:0] _T_659; // @[CSR.scala 281:64:@4970.4]
  wire [31:0] _T_660; // @[CSR.scala 281:60:@4971.4]
  wire [31:0] wdata; // @[CSR.scala 281:58:@4972.4]
  wire [2:0] _T_662; // @[CSR.scala 185:33:@4973.4]
  wire [7:0] opcode; // @[CSR.scala 185:20:@4974.4]
  wire  _T_663; // @[CSR.scala 186:40:@4975.4]
  wire  insn_call; // @[CSR.scala 186:31:@4976.4]
  wire  _T_664; // @[CSR.scala 187:41:@4977.4]
  wire  insn_break; // @[CSR.scala 187:32:@4978.4]
  wire  _T_665; // @[CSR.scala 188:39:@4979.4]
  wire  _T_666; // @[CSR.scala 188:30:@4980.4]
  wire  insn_ret; // @[CSR.scala 188:43:@4981.4]
  wire  _T_940; // @[CSR.scala 199:24:@5180.4]
  wire [1:0] _T_942; // @[Bitwise.scala 48:55:@5183.4]
  wire  _T_944; // @[CSR.scala 201:50:@5184.4]
  wire  _T_946; // @[CSR.scala 201:9:@5186.4]
  wire  _T_948; // @[CSR.scala 201:9:@5187.4]
  wire  _T_951; // @[CSR.scala 208:32:@5196.4]
  wire  _T_953; // @[CSR.scala 208:21:@5197.4]
  wire  _T_954; // @[CSR.scala 208:18:@5198.4]
  wire  _GEN_3; // @[CSR.scala 208:38:@5199.4]
  wire  _GEN_4; // @[CSR.scala 208:38:@5199.4]
  wire [1:0] new_prv; // @[CSR.scala 208:38:@5199.4]
  wire [3:0] _GEN_148; // @[CSR.scala 218:35:@5207.6]
  wire [4:0] _T_958; // @[CSR.scala 218:35:@5207.6]
  wire [3:0] _T_959; // @[CSR.scala 218:35:@5208.6]
  wire [31:0] _GEN_7; // @[CSR.scala 216:18:@5205.4]
  wire [31:0] _GEN_8; // @[CSR.scala 216:18:@5205.4]
  wire [31:0] _GEN_9; // @[CSR.scala 216:18:@5205.4]
  wire [31:0] _GEN_10; // @[CSR.scala 223:19:@5212.4]
  wire [31:0] _GEN_11; // @[CSR.scala 223:19:@5212.4]
  wire [31:0] _GEN_12; // @[CSR.scala 223:19:@5212.4]
  wire [31:0] _GEN_14; // @[CSR.scala 229:17:@5217.4]
  wire [31:0] _GEN_15; // @[CSR.scala 229:17:@5217.4]
  wire [31:0] _GEN_16; // @[CSR.scala 229:17:@5217.4]
  wire [63:0] _T_965; // @[Mux.scala 19:72:@5225.4]
  wire [63:0] _T_967; // @[Mux.scala 19:72:@5226.4]
  wire [15:0] _T_969; // @[Mux.scala 19:72:@5227.4]
  wire [30:0] _T_975; // @[Mux.scala 19:72:@5230.4]
  wire [31:0] _T_977; // @[Mux.scala 19:72:@5231.4]
  wire [8:0] _T_979; // @[Mux.scala 19:72:@5232.4]
  wire [15:0] _T_981; // @[Mux.scala 19:72:@5233.4]
  wire [15:0] _T_983; // @[Mux.scala 19:72:@5234.4]
  wire [31:0] _T_985; // @[Mux.scala 19:72:@5235.4]
  wire [31:0] _T_987; // @[Mux.scala 19:72:@5236.4]
  wire [31:0] _T_989; // @[Mux.scala 19:72:@5237.4]
  wire [31:0] _T_991; // @[Mux.scala 19:72:@5238.4]
  wire [31:0] _T_995; // @[Mux.scala 19:72:@5240.4]
  wire [31:0] _T_997; // @[Mux.scala 19:72:@5241.4]
  wire [39:0] _T_999; // @[Mux.scala 19:72:@5242.4]
  wire [39:0] _T_1001; // @[Mux.scala 19:72:@5243.4]
  wire [39:0] _T_1003; // @[Mux.scala 19:72:@5244.4]
  wire [39:0] _T_1005; // @[Mux.scala 19:72:@5245.4]
  wire [39:0] _T_1007; // @[Mux.scala 19:72:@5246.4]
  wire [39:0] _T_1009; // @[Mux.scala 19:72:@5247.4]
  wire [39:0] _T_1011; // @[Mux.scala 19:72:@5248.4]
  wire [39:0] _T_1013; // @[Mux.scala 19:72:@5249.4]
  wire [39:0] _T_1015; // @[Mux.scala 19:72:@5250.4]
  wire [39:0] _T_1017; // @[Mux.scala 19:72:@5251.4]
  wire [39:0] _T_1019; // @[Mux.scala 19:72:@5252.4]
  wire [39:0] _T_1021; // @[Mux.scala 19:72:@5253.4]
  wire [39:0] _T_1023; // @[Mux.scala 19:72:@5254.4]
  wire [39:0] _T_1025; // @[Mux.scala 19:72:@5255.4]
  wire [39:0] _T_1027; // @[Mux.scala 19:72:@5256.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:@5257.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:@5258.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:@5259.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:@5260.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:@5261.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:@5262.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:@5263.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:@5264.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:@5265.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:@5266.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:@5267.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:@5268.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:@5269.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:@5270.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:@5271.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:@5272.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:@5273.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:@5274.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:@5275.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:@5276.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:@5277.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:@5278.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:@5279.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:@5280.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:@5281.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:@5282.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:@5283.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:@5284.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:@5285.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:@5286.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:@5287.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:@5288.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:@5289.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:@5290.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:@5291.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:@5292.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:@5293.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:@5294.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:@5295.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:@5296.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:@5297.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:@5298.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:@5299.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:@5300.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:@5301.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:@5302.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:@5303.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:@5304.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:@5305.4]
  wire [63:0] _T_1130; // @[Mux.scala 19:72:@5308.4]
  wire [63:0] _GEN_149; // @[Mux.scala 19:72:@5309.4]
  wire [63:0] _T_1131; // @[Mux.scala 19:72:@5309.4]
  wire [63:0] _GEN_150; // @[Mux.scala 19:72:@5312.4]
  wire [63:0] _T_1134; // @[Mux.scala 19:72:@5312.4]
  wire [63:0] _GEN_151; // @[Mux.scala 19:72:@5313.4]
  wire [63:0] _T_1135; // @[Mux.scala 19:72:@5313.4]
  wire [63:0] _GEN_152; // @[Mux.scala 19:72:@5314.4]
  wire [63:0] _T_1136; // @[Mux.scala 19:72:@5314.4]
  wire [63:0] _GEN_153; // @[Mux.scala 19:72:@5315.4]
  wire [63:0] _T_1137; // @[Mux.scala 19:72:@5315.4]
  wire [63:0] _GEN_154; // @[Mux.scala 19:72:@5316.4]
  wire [63:0] _T_1138; // @[Mux.scala 19:72:@5316.4]
  wire [63:0] _GEN_155; // @[Mux.scala 19:72:@5317.4]
  wire [63:0] _T_1139; // @[Mux.scala 19:72:@5317.4]
  wire [63:0] _GEN_156; // @[Mux.scala 19:72:@5318.4]
  wire [63:0] _T_1140; // @[Mux.scala 19:72:@5318.4]
  wire [63:0] _GEN_157; // @[Mux.scala 19:72:@5319.4]
  wire [63:0] _T_1141; // @[Mux.scala 19:72:@5319.4]
  wire [63:0] _GEN_158; // @[Mux.scala 19:72:@5320.4]
  wire [63:0] _T_1142; // @[Mux.scala 19:72:@5320.4]
  wire [63:0] _GEN_159; // @[Mux.scala 19:72:@5322.4]
  wire [63:0] _T_1144; // @[Mux.scala 19:72:@5322.4]
  wire [63:0] _GEN_160; // @[Mux.scala 19:72:@5323.4]
  wire [63:0] _T_1145; // @[Mux.scala 19:72:@5323.4]
  wire [63:0] _GEN_161; // @[Mux.scala 19:72:@5324.4]
  wire [63:0] _T_1146; // @[Mux.scala 19:72:@5324.4]
  wire [63:0] _GEN_162; // @[Mux.scala 19:72:@5325.4]
  wire [63:0] _T_1147; // @[Mux.scala 19:72:@5325.4]
  wire [63:0] _GEN_163; // @[Mux.scala 19:72:@5326.4]
  wire [63:0] _T_1148; // @[Mux.scala 19:72:@5326.4]
  wire [63:0] _GEN_164; // @[Mux.scala 19:72:@5327.4]
  wire [63:0] _T_1149; // @[Mux.scala 19:72:@5327.4]
  wire [63:0] _GEN_165; // @[Mux.scala 19:72:@5328.4]
  wire [63:0] _T_1150; // @[Mux.scala 19:72:@5328.4]
  wire [63:0] _GEN_166; // @[Mux.scala 19:72:@5329.4]
  wire [63:0] _T_1151; // @[Mux.scala 19:72:@5329.4]
  wire [63:0] _GEN_167; // @[Mux.scala 19:72:@5330.4]
  wire [63:0] _T_1152; // @[Mux.scala 19:72:@5330.4]
  wire [63:0] _GEN_168; // @[Mux.scala 19:72:@5331.4]
  wire [63:0] _T_1153; // @[Mux.scala 19:72:@5331.4]
  wire [63:0] _GEN_169; // @[Mux.scala 19:72:@5332.4]
  wire [63:0] _T_1154; // @[Mux.scala 19:72:@5332.4]
  wire [63:0] _GEN_170; // @[Mux.scala 19:72:@5333.4]
  wire [63:0] _T_1155; // @[Mux.scala 19:72:@5333.4]
  wire [63:0] _GEN_171; // @[Mux.scala 19:72:@5334.4]
  wire [63:0] _T_1156; // @[Mux.scala 19:72:@5334.4]
  wire [63:0] _GEN_172; // @[Mux.scala 19:72:@5335.4]
  wire [63:0] _T_1157; // @[Mux.scala 19:72:@5335.4]
  wire [63:0] _GEN_173; // @[Mux.scala 19:72:@5336.4]
  wire [63:0] _T_1158; // @[Mux.scala 19:72:@5336.4]
  wire [63:0] _GEN_174; // @[Mux.scala 19:72:@5337.4]
  wire [63:0] _T_1159; // @[Mux.scala 19:72:@5337.4]
  wire [63:0] _GEN_175; // @[Mux.scala 19:72:@5338.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:@5338.4]
  wire [63:0] _GEN_176; // @[Mux.scala 19:72:@5339.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:@5339.4]
  wire [63:0] _GEN_177; // @[Mux.scala 19:72:@5340.4]
  wire [63:0] _T_1162; // @[Mux.scala 19:72:@5340.4]
  wire [63:0] _GEN_178; // @[Mux.scala 19:72:@5341.4]
  wire [63:0] _T_1163; // @[Mux.scala 19:72:@5341.4]
  wire [63:0] _GEN_179; // @[Mux.scala 19:72:@5342.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:@5342.4]
  wire [63:0] _GEN_180; // @[Mux.scala 19:72:@5343.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:@5343.4]
  wire [63:0] _GEN_181; // @[Mux.scala 19:72:@5344.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:@5344.4]
  wire [63:0] _GEN_182; // @[Mux.scala 19:72:@5345.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:@5345.4]
  wire [63:0] _GEN_183; // @[Mux.scala 19:72:@5346.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:@5346.4]
  wire [63:0] _GEN_184; // @[Mux.scala 19:72:@5347.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:@5347.4]
  wire [63:0] _GEN_185; // @[Mux.scala 19:72:@5348.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:@5348.4]
  wire [63:0] _GEN_186; // @[Mux.scala 19:72:@5349.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:@5349.4]
  wire [63:0] _GEN_187; // @[Mux.scala 19:72:@5350.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:@5350.4]
  wire [63:0] _GEN_188; // @[Mux.scala 19:72:@5351.4]
  wire [63:0] _T_1173; // @[Mux.scala 19:72:@5351.4]
  wire [63:0] _GEN_189; // @[Mux.scala 19:72:@5352.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:@5352.4]
  wire [63:0] _GEN_190; // @[Mux.scala 19:72:@5353.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:@5353.4]
  wire [63:0] _GEN_191; // @[Mux.scala 19:72:@5354.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:@5354.4]
  wire [63:0] _GEN_192; // @[Mux.scala 19:72:@5355.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:@5355.4]
  wire [63:0] _GEN_193; // @[Mux.scala 19:72:@5356.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:@5356.4]
  wire [63:0] _GEN_194; // @[Mux.scala 19:72:@5357.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:@5357.4]
  wire [63:0] _GEN_195; // @[Mux.scala 19:72:@5358.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:@5358.4]
  wire [63:0] _GEN_196; // @[Mux.scala 19:72:@5359.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:@5359.4]
  wire [63:0] _GEN_197; // @[Mux.scala 19:72:@5360.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:@5360.4]
  wire [63:0] _GEN_198; // @[Mux.scala 19:72:@5361.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:@5361.4]
  wire [63:0] _GEN_199; // @[Mux.scala 19:72:@5362.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:@5362.4]
  wire [63:0] _GEN_200; // @[Mux.scala 19:72:@5363.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:@5363.4]
  wire [63:0] _GEN_201; // @[Mux.scala 19:72:@5364.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:@5364.4]
  wire [63:0] _GEN_202; // @[Mux.scala 19:72:@5365.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:@5365.4]
  wire [63:0] _GEN_203; // @[Mux.scala 19:72:@5366.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:@5366.4]
  wire [63:0] _GEN_204; // @[Mux.scala 19:72:@5367.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:@5367.4]
  wire [63:0] _GEN_205; // @[Mux.scala 19:72:@5368.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:@5368.4]
  wire [63:0] _GEN_206; // @[Mux.scala 19:72:@5369.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:@5369.4]
  wire [63:0] _GEN_207; // @[Mux.scala 19:72:@5370.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:@5370.4]
  wire [63:0] _GEN_208; // @[Mux.scala 19:72:@5371.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:@5371.4]
  wire [63:0] _GEN_209; // @[Mux.scala 19:72:@5372.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:@5372.4]
  wire [63:0] _GEN_210; // @[Mux.scala 19:72:@5373.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:@5373.4]
  wire [63:0] _GEN_211; // @[Mux.scala 19:72:@5374.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:@5374.4]
  wire [63:0] _GEN_212; // @[Mux.scala 19:72:@5375.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:@5375.4]
  wire [63:0] _GEN_213; // @[Mux.scala 19:72:@5376.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:@5376.4]
  wire [63:0] _GEN_214; // @[Mux.scala 19:72:@5377.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:@5377.4]
  wire [63:0] _GEN_215; // @[Mux.scala 19:72:@5378.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:@5378.4]
  wire [63:0] _GEN_216; // @[Mux.scala 19:72:@5379.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:@5379.4]
  wire [63:0] _GEN_217; // @[Mux.scala 19:72:@5380.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:@5380.4]
  wire [63:0] _GEN_218; // @[Mux.scala 19:72:@5381.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:@5381.4]
  wire [63:0] _GEN_219; // @[Mux.scala 19:72:@5382.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:@5382.4]
  wire [63:0] _GEN_220; // @[Mux.scala 19:72:@5383.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:@5383.4]
  wire [63:0] _GEN_221; // @[Mux.scala 19:72:@5384.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:@5384.4]
  wire [63:0] _GEN_222; // @[Mux.scala 19:72:@5385.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:@5385.4]
  wire [63:0] _GEN_223; // @[Mux.scala 19:72:@5386.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:@5386.4]
  wire [63:0] _GEN_224; // @[Mux.scala 19:72:@5387.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:@5387.4]
  wire  _T_1220; // @[CSR.scala 245:39:@5400.8]
  wire  _T_1222; // @[CSR.scala 245:39:@5404.8]
  wire  _GEN_17; // @[CSR.scala 244:39:@5394.6]
  wire  _GEN_18; // @[CSR.scala 244:39:@5394.6]
  wire [15:0] _T_1233; // @[:@5423.8 :@5424.8]
  wire  _T_1235; // @[CSR.scala 250:35:@5427.8]
  wire  _T_1237; // @[CSR.scala 250:35:@5431.8]
  wire  _GEN_19; // @[CSR.scala 249:35:@5421.6]
  wire  _GEN_20; // @[CSR.scala 253:35:@5441.6]
  wire  _GEN_21; // @[CSR.scala 253:35:@5441.6]
  wire [7:0] _T_1253; // @[CSR.scala 277:47:@5463.8]
  wire [31:0] _T_1254; // @[CSR.scala 277:72:@5464.8]
  wire [39:0] _T_1255; // @[Cat.scala 30:58:@5465.8]
  wire [40:0] _GEN_22; // @[CSR.scala 277:29:@5462.6]
  wire [7:0] _T_1256; // @[CSR.scala 278:45:@5469.8]
  wire [39:0] _T_1257; // @[Cat.scala 30:58:@5470.8]
  wire [40:0] _GEN_23; // @[CSR.scala 278:29:@5468.6]
  wire [31:0] _T_1259; // @[CSR.scala 277:72:@5475.8]
  wire [39:0] _T_1260; // @[Cat.scala 30:58:@5476.8]
  wire [40:0] _GEN_24; // @[CSR.scala 277:29:@5473.6]
  wire [7:0] _T_1261; // @[CSR.scala 278:45:@5480.8]
  wire [39:0] _T_1262; // @[Cat.scala 30:58:@5481.8]
  wire [40:0] _GEN_25; // @[CSR.scala 278:29:@5479.6]
  wire [31:0] _T_1264; // @[CSR.scala 277:72:@5486.8]
  wire [39:0] _T_1265; // @[Cat.scala 30:58:@5487.8]
  wire [40:0] _GEN_26; // @[CSR.scala 277:29:@5484.6]
  wire [7:0] _T_1266; // @[CSR.scala 278:45:@5491.8]
  wire [39:0] _T_1267; // @[Cat.scala 30:58:@5492.8]
  wire [40:0] _GEN_27; // @[CSR.scala 278:29:@5490.6]
  wire [31:0] _T_1269; // @[CSR.scala 277:72:@5497.8]
  wire [39:0] _T_1270; // @[Cat.scala 30:58:@5498.8]
  wire [40:0] _GEN_28; // @[CSR.scala 277:29:@5495.6]
  wire [7:0] _T_1271; // @[CSR.scala 278:45:@5502.8]
  wire [39:0] _T_1272; // @[Cat.scala 30:58:@5503.8]
  wire [40:0] _GEN_29; // @[CSR.scala 278:29:@5501.6]
  wire [31:0] _T_1274; // @[CSR.scala 277:72:@5508.8]
  wire [39:0] _T_1275; // @[Cat.scala 30:58:@5509.8]
  wire [40:0] _GEN_30; // @[CSR.scala 277:29:@5506.6]
  wire [7:0] _T_1276; // @[CSR.scala 278:45:@5513.8]
  wire [39:0] _T_1277; // @[Cat.scala 30:58:@5514.8]
  wire [40:0] _GEN_31; // @[CSR.scala 278:29:@5512.6]
  wire [31:0] _T_1279; // @[CSR.scala 277:72:@5519.8]
  wire [39:0] _T_1280; // @[Cat.scala 30:58:@5520.8]
  wire [40:0] _GEN_32; // @[CSR.scala 277:29:@5517.6]
  wire [7:0] _T_1281; // @[CSR.scala 278:45:@5524.8]
  wire [39:0] _T_1282; // @[Cat.scala 30:58:@5525.8]
  wire [40:0] _GEN_33; // @[CSR.scala 278:29:@5523.6]
  wire [31:0] _T_1284; // @[CSR.scala 277:72:@5530.8]
  wire [39:0] _T_1285; // @[Cat.scala 30:58:@5531.8]
  wire [40:0] _GEN_34; // @[CSR.scala 277:29:@5528.6]
  wire [7:0] _T_1286; // @[CSR.scala 278:45:@5535.8]
  wire [39:0] _T_1287; // @[Cat.scala 30:58:@5536.8]
  wire [40:0] _GEN_35; // @[CSR.scala 278:29:@5534.6]
  wire [31:0] _T_1289; // @[CSR.scala 277:72:@5541.8]
  wire [39:0] _T_1290; // @[Cat.scala 30:58:@5542.8]
  wire [40:0] _GEN_36; // @[CSR.scala 277:29:@5539.6]
  wire [7:0] _T_1291; // @[CSR.scala 278:45:@5546.8]
  wire [39:0] _T_1292; // @[Cat.scala 30:58:@5547.8]
  wire [40:0] _GEN_37; // @[CSR.scala 278:29:@5545.6]
  wire [31:0] _T_1294; // @[CSR.scala 277:72:@5552.8]
  wire [39:0] _T_1295; // @[Cat.scala 30:58:@5553.8]
  wire [40:0] _GEN_38; // @[CSR.scala 277:29:@5550.6]
  wire [7:0] _T_1296; // @[CSR.scala 278:45:@5557.8]
  wire [39:0] _T_1297; // @[Cat.scala 30:58:@5558.8]
  wire [40:0] _GEN_39; // @[CSR.scala 278:29:@5556.6]
  wire [31:0] _T_1299; // @[CSR.scala 277:72:@5563.8]
  wire [39:0] _T_1300; // @[Cat.scala 30:58:@5564.8]
  wire [40:0] _GEN_40; // @[CSR.scala 277:29:@5561.6]
  wire [7:0] _T_1301; // @[CSR.scala 278:45:@5568.8]
  wire [39:0] _T_1302; // @[Cat.scala 30:58:@5569.8]
  wire [40:0] _GEN_41; // @[CSR.scala 278:29:@5567.6]
  wire [31:0] _T_1304; // @[CSR.scala 277:72:@5574.8]
  wire [39:0] _T_1305; // @[Cat.scala 30:58:@5575.8]
  wire [40:0] _GEN_42; // @[CSR.scala 277:29:@5572.6]
  wire [7:0] _T_1306; // @[CSR.scala 278:45:@5579.8]
  wire [39:0] _T_1307; // @[Cat.scala 30:58:@5580.8]
  wire [40:0] _GEN_43; // @[CSR.scala 278:29:@5578.6]
  wire [31:0] _T_1309; // @[CSR.scala 277:72:@5585.8]
  wire [39:0] _T_1310; // @[Cat.scala 30:58:@5586.8]
  wire [40:0] _GEN_44; // @[CSR.scala 277:29:@5583.6]
  wire [7:0] _T_1311; // @[CSR.scala 278:45:@5590.8]
  wire [39:0] _T_1312; // @[Cat.scala 30:58:@5591.8]
  wire [40:0] _GEN_45; // @[CSR.scala 278:29:@5589.6]
  wire [31:0] _T_1314; // @[CSR.scala 277:72:@5596.8]
  wire [39:0] _T_1315; // @[Cat.scala 30:58:@5597.8]
  wire [40:0] _GEN_46; // @[CSR.scala 277:29:@5594.6]
  wire [7:0] _T_1316; // @[CSR.scala 278:45:@5601.8]
  wire [39:0] _T_1317; // @[Cat.scala 30:58:@5602.8]
  wire [40:0] _GEN_47; // @[CSR.scala 278:29:@5600.6]
  wire [31:0] _T_1319; // @[CSR.scala 277:72:@5607.8]
  wire [39:0] _T_1320; // @[Cat.scala 30:58:@5608.8]
  wire [40:0] _GEN_48; // @[CSR.scala 277:29:@5605.6]
  wire [7:0] _T_1321; // @[CSR.scala 278:45:@5612.8]
  wire [39:0] _T_1322; // @[Cat.scala 30:58:@5613.8]
  wire [40:0] _GEN_49; // @[CSR.scala 278:29:@5611.6]
  wire [31:0] _T_1324; // @[CSR.scala 277:72:@5618.8]
  wire [39:0] _T_1325; // @[Cat.scala 30:58:@5619.8]
  wire [40:0] _GEN_50; // @[CSR.scala 277:29:@5616.6]
  wire [7:0] _T_1326; // @[CSR.scala 278:45:@5623.8]
  wire [39:0] _T_1327; // @[Cat.scala 30:58:@5624.8]
  wire [40:0] _GEN_51; // @[CSR.scala 278:29:@5622.6]
  wire [31:0] _T_1329; // @[CSR.scala 277:72:@5629.8]
  wire [39:0] _T_1330; // @[Cat.scala 30:58:@5630.8]
  wire [40:0] _GEN_52; // @[CSR.scala 277:29:@5627.6]
  wire [7:0] _T_1331; // @[CSR.scala 278:45:@5634.8]
  wire [39:0] _T_1332; // @[Cat.scala 30:58:@5635.8]
  wire [40:0] _GEN_53; // @[CSR.scala 278:29:@5633.6]
  wire [31:0] _T_1334; // @[CSR.scala 277:72:@5640.8]
  wire [39:0] _T_1335; // @[Cat.scala 30:58:@5641.8]
  wire [40:0] _GEN_54; // @[CSR.scala 277:29:@5638.6]
  wire [7:0] _T_1336; // @[CSR.scala 278:45:@5645.8]
  wire [39:0] _T_1337; // @[Cat.scala 30:58:@5646.8]
  wire [40:0] _GEN_55; // @[CSR.scala 278:29:@5644.6]
  wire [31:0] _T_1339; // @[CSR.scala 277:72:@5651.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:@5652.8]
  wire [40:0] _GEN_56; // @[CSR.scala 277:29:@5649.6]
  wire [7:0] _T_1341; // @[CSR.scala 278:45:@5656.8]
  wire [39:0] _T_1342; // @[Cat.scala 30:58:@5657.8]
  wire [40:0] _GEN_57; // @[CSR.scala 278:29:@5655.6]
  wire [31:0] _T_1344; // @[CSR.scala 277:72:@5662.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:@5663.8]
  wire [40:0] _GEN_58; // @[CSR.scala 277:29:@5660.6]
  wire [7:0] _T_1346; // @[CSR.scala 278:45:@5667.8]
  wire [39:0] _T_1347; // @[Cat.scala 30:58:@5668.8]
  wire [40:0] _GEN_59; // @[CSR.scala 278:29:@5666.6]
  wire [31:0] _T_1349; // @[CSR.scala 277:72:@5673.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:@5674.8]
  wire [40:0] _GEN_60; // @[CSR.scala 277:29:@5671.6]
  wire [7:0] _T_1351; // @[CSR.scala 278:45:@5678.8]
  wire [39:0] _T_1352; // @[Cat.scala 30:58:@5679.8]
  wire [40:0] _GEN_61; // @[CSR.scala 278:29:@5677.6]
  wire [31:0] _T_1354; // @[CSR.scala 277:72:@5684.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:@5685.8]
  wire [40:0] _GEN_62; // @[CSR.scala 277:29:@5682.6]
  wire [7:0] _T_1356; // @[CSR.scala 278:45:@5689.8]
  wire [39:0] _T_1357; // @[Cat.scala 30:58:@5690.8]
  wire [40:0] _GEN_63; // @[CSR.scala 278:29:@5688.6]
  wire [31:0] _T_1359; // @[CSR.scala 277:72:@5695.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:@5696.8]
  wire [40:0] _GEN_64; // @[CSR.scala 277:29:@5693.6]
  wire [7:0] _T_1361; // @[CSR.scala 278:45:@5700.8]
  wire [39:0] _T_1362; // @[Cat.scala 30:58:@5701.8]
  wire [40:0] _GEN_65; // @[CSR.scala 278:29:@5699.6]
  wire [31:0] _T_1364; // @[CSR.scala 277:72:@5706.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:@5707.8]
  wire [40:0] _GEN_66; // @[CSR.scala 277:29:@5704.6]
  wire [7:0] _T_1366; // @[CSR.scala 278:45:@5711.8]
  wire [39:0] _T_1367; // @[Cat.scala 30:58:@5712.8]
  wire [40:0] _GEN_67; // @[CSR.scala 278:29:@5710.6]
  wire [31:0] _T_1369; // @[CSR.scala 277:72:@5717.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:@5718.8]
  wire [40:0] _GEN_68; // @[CSR.scala 277:29:@5715.6]
  wire [7:0] _T_1371; // @[CSR.scala 278:45:@5722.8]
  wire [39:0] _T_1372; // @[Cat.scala 30:58:@5723.8]
  wire [40:0] _GEN_69; // @[CSR.scala 278:29:@5721.6]
  wire [31:0] _T_1374; // @[CSR.scala 277:72:@5728.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:@5729.8]
  wire [40:0] _GEN_70; // @[CSR.scala 277:29:@5726.6]
  wire [7:0] _T_1376; // @[CSR.scala 278:45:@5733.8]
  wire [39:0] _T_1377; // @[Cat.scala 30:58:@5734.8]
  wire [40:0] _GEN_71; // @[CSR.scala 278:29:@5732.6]
  wire [31:0] _T_1379; // @[CSR.scala 277:72:@5739.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:@5740.8]
  wire [40:0] _GEN_72; // @[CSR.scala 277:29:@5737.6]
  wire [7:0] _T_1381; // @[CSR.scala 278:45:@5744.8]
  wire [39:0] _T_1382; // @[Cat.scala 30:58:@5745.8]
  wire [40:0] _GEN_73; // @[CSR.scala 278:29:@5743.6]
  wire [31:0] _T_1384; // @[CSR.scala 277:72:@5750.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:@5751.8]
  wire [40:0] _GEN_74; // @[CSR.scala 277:29:@5748.6]
  wire [7:0] _T_1386; // @[CSR.scala 278:45:@5755.8]
  wire [39:0] _T_1387; // @[Cat.scala 30:58:@5756.8]
  wire [40:0] _GEN_75; // @[CSR.scala 278:29:@5754.6]
  wire [31:0] _T_1389; // @[CSR.scala 277:72:@5761.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:@5762.8]
  wire [40:0] _GEN_76; // @[CSR.scala 277:29:@5759.6]
  wire [7:0] _T_1391; // @[CSR.scala 278:45:@5766.8]
  wire [39:0] _T_1392; // @[Cat.scala 30:58:@5767.8]
  wire [40:0] _GEN_77; // @[CSR.scala 278:29:@5765.6]
  wire [31:0] _T_1394; // @[CSR.scala 277:72:@5772.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:@5773.8]
  wire [40:0] _GEN_78; // @[CSR.scala 277:29:@5770.6]
  wire [7:0] _T_1396; // @[CSR.scala 278:45:@5777.8]
  wire [39:0] _T_1397; // @[Cat.scala 30:58:@5778.8]
  wire [40:0] _GEN_79; // @[CSR.scala 278:29:@5776.6]
  wire [31:0] _T_1399; // @[CSR.scala 277:72:@5783.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:@5784.8]
  wire [40:0] _GEN_80; // @[CSR.scala 277:29:@5781.6]
  wire [7:0] _T_1401; // @[CSR.scala 278:45:@5788.8]
  wire [39:0] _T_1402; // @[Cat.scala 30:58:@5789.8]
  wire [40:0] _GEN_81; // @[CSR.scala 278:29:@5787.6]
  wire [31:0] _T_1404; // @[CSR.scala 277:72:@5794.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:@5795.8]
  wire [40:0] _GEN_82; // @[CSR.scala 277:29:@5792.6]
  wire [7:0] _T_1406; // @[CSR.scala 278:45:@5799.8]
  wire [39:0] _T_1407; // @[Cat.scala 30:58:@5800.8]
  wire [40:0] _GEN_83; // @[CSR.scala 278:29:@5798.6]
  wire [31:0] _T_1409; // @[CSR.scala 277:72:@5805.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:@5806.8]
  wire [40:0] _GEN_84; // @[CSR.scala 277:29:@5803.6]
  wire [7:0] _T_1411; // @[CSR.scala 278:45:@5810.8]
  wire [39:0] _T_1412; // @[Cat.scala 30:58:@5811.8]
  wire [40:0] _GEN_85; // @[CSR.scala 278:29:@5809.6]
  wire [31:0] _T_1414; // @[CSR.scala 277:72:@5816.8]
  wire [63:0] _T_1415; // @[Cat.scala 30:58:@5817.8]
  wire [57:0] _T_1416; // @[Util.scala 133:28:@5819.8]
  wire [63:0] _GEN_86; // @[CSR.scala 277:29:@5814.6]
  wire [57:0] _GEN_87; // @[CSR.scala 277:29:@5814.6]
  wire [31:0] _T_1417; // @[CSR.scala 278:45:@5823.8]
  wire [63:0] _T_1418; // @[Cat.scala 30:58:@5824.8]
  wire [57:0] _T_1419; // @[Util.scala 133:28:@5826.8]
  wire [63:0] _GEN_88; // @[CSR.scala 278:29:@5822.6]
  wire [57:0] _GEN_89; // @[CSR.scala 278:29:@5822.6]
  wire [31:0] _T_1421; // @[CSR.scala 277:72:@5831.8]
  wire [63:0] _T_1422; // @[Cat.scala 30:58:@5832.8]
  wire [57:0] _T_1423; // @[Util.scala 133:28:@5834.8]
  wire [63:0] _GEN_90; // @[CSR.scala 277:29:@5829.6]
  wire [57:0] _GEN_91; // @[CSR.scala 277:29:@5829.6]
  wire [31:0] _T_1424; // @[CSR.scala 278:45:@5838.8]
  wire [63:0] _T_1425; // @[Cat.scala 30:58:@5839.8]
  wire [57:0] _T_1426; // @[Util.scala 133:28:@5841.8]
  wire [63:0] _GEN_92; // @[CSR.scala 278:29:@5837.6]
  wire [57:0] _GEN_93; // @[CSR.scala 278:29:@5837.6]
  wire [31:0] _GEN_94; // @[CSR.scala 265:40:@5844.6]
  wire [31:0] _T_1429; // @[CSR.scala 267:78:@5849.8]
  wire [34:0] _GEN_225; // @[CSR.scala 267:86:@5850.8]
  wire [34:0] _T_1431; // @[CSR.scala 267:86:@5850.8]
  wire [34:0] _GEN_95; // @[CSR.scala 267:40:@5847.6]
  wire [31:0] _GEN_96; // @[CSR.scala 268:40:@5853.6]
  wire [31:0] _T_1433; // @[CSR.scala 269:62:@5857.8]
  wire [31:0] _GEN_97; // @[CSR.scala 269:40:@5856.6]
  wire [31:0] _GEN_98; // @[CSR.scala 270:40:@5860.6]
  wire [31:0] _GEN_99; // @[CSR.scala 271:42:@5864.6]
  wire  _GEN_100; // @[CSR.scala 242:14:@5393.4]
  wire  _GEN_101; // @[CSR.scala 242:14:@5393.4]
  wire  _GEN_102; // @[CSR.scala 242:14:@5393.4]
  wire  _GEN_103; // @[CSR.scala 242:14:@5393.4]
  wire  _GEN_104; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_105; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_106; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_107; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_108; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_109; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_110; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_111; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_112; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_113; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_114; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_115; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_116; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_117; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_118; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_119; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_120; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_121; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_122; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_123; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_124; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_125; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_126; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_127; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_128; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_129; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_130; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_131; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_132; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_133; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_134; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_135; // @[CSR.scala 242:14:@5393.4]
  wire [40:0] _GEN_136; // @[CSR.scala 242:14:@5393.4]
  wire [63:0] _GEN_137; // @[CSR.scala 242:14:@5393.4]
  wire [57:0] _GEN_138; // @[CSR.scala 242:14:@5393.4]
  wire [63:0] _GEN_139; // @[CSR.scala 242:14:@5393.4]
  wire [57:0] _GEN_140; // @[CSR.scala 242:14:@5393.4]
  wire [34:0] _GEN_142; // @[CSR.scala 242:14:@5393.4]
  assign _T_241 = _T_240 + 6'h1; // @[Util.scala 113:33:@4639.4]
  assign _T_245 = _T_241[6]; // @[Util.scala 118:20:@4642.4]
  assign _T_247 = _T_244 + 58'h1; // @[Util.scala 118:43:@4644.6]
  assign _T_248 = _T_244 + 58'h1; // @[Util.scala 118:43:@4645.6]
  assign _GEN_0 = _T_245 ? _T_248 : _T_244; // @[Util.scala 118:34:@4643.4]
  assign _T_249 = {_T_244,_T_240}; // @[Cat.scala 30:58:@4648.4]
  assign _GEN_147 = {{4'd0}, io_retire}; // @[Util.scala 113:33:@4650.4]
  assign _T_253 = _T_252 + _GEN_147; // @[Util.scala 113:33:@4650.4]
  assign _T_257 = _T_253[6]; // @[Util.scala 118:20:@4653.4]
  assign _T_259 = _T_256 + 58'h1; // @[Util.scala 118:43:@4655.6]
  assign _T_260 = _T_256 + 58'h1; // @[Util.scala 118:43:@4656.6]
  assign _GEN_1 = _T_257 ? _T_260 : _T_256; // @[Util.scala 118:34:@4654.4]
  assign _T_261 = {_T_256,_T_252}; // @[Cat.scala 30:58:@4659.4]
  assign _T_265 = {{1'd0}, _T_264}; // @[Util.scala 113:33:@4662.4]
  assign _T_268 = {{1'd0}, _T_267}; // @[Util.scala 113:33:@4665.4]
  assign _T_271 = {{1'd0}, _T_270}; // @[Util.scala 113:33:@4668.4]
  assign _T_274 = {{1'd0}, _T_273}; // @[Util.scala 113:33:@4671.4]
  assign _T_277 = {{1'd0}, _T_276}; // @[Util.scala 113:33:@4674.4]
  assign _T_280 = {{1'd0}, _T_279}; // @[Util.scala 113:33:@4677.4]
  assign _T_283 = {{1'd0}, _T_282}; // @[Util.scala 113:33:@4680.4]
  assign _T_286 = {{1'd0}, _T_285}; // @[Util.scala 113:33:@4683.4]
  assign _T_289 = {{1'd0}, _T_288}; // @[Util.scala 113:33:@4686.4]
  assign _T_292 = {{1'd0}, _T_291}; // @[Util.scala 113:33:@4689.4]
  assign _T_295 = {{1'd0}, _T_294}; // @[Util.scala 113:33:@4692.4]
  assign _T_298 = {{1'd0}, _T_297}; // @[Util.scala 113:33:@4695.4]
  assign _T_301 = {{1'd0}, _T_300}; // @[Util.scala 113:33:@4698.4]
  assign _T_304 = {{1'd0}, _T_303}; // @[Util.scala 113:33:@4701.4]
  assign _T_307 = {{1'd0}, _T_306}; // @[Util.scala 113:33:@4704.4]
  assign _T_310 = {{1'd0}, _T_309}; // @[Util.scala 113:33:@4707.4]
  assign _T_313 = {{1'd0}, _T_312}; // @[Util.scala 113:33:@4710.4]
  assign _T_316 = {{1'd0}, _T_315}; // @[Util.scala 113:33:@4713.4]
  assign _T_319 = {{1'd0}, _T_318}; // @[Util.scala 113:33:@4716.4]
  assign _T_322 = {{1'd0}, _T_321}; // @[Util.scala 113:33:@4719.4]
  assign _T_325 = {{1'd0}, _T_324}; // @[Util.scala 113:33:@4722.4]
  assign _T_328 = {{1'd0}, _T_327}; // @[Util.scala 113:33:@4725.4]
  assign _T_331 = {{1'd0}, _T_330}; // @[Util.scala 113:33:@4728.4]
  assign _T_334 = {{1'd0}, _T_333}; // @[Util.scala 113:33:@4731.4]
  assign _T_337 = {{1'd0}, _T_336}; // @[Util.scala 113:33:@4734.4]
  assign _T_340 = {{1'd0}, _T_339}; // @[Util.scala 113:33:@4737.4]
  assign _T_343 = {{1'd0}, _T_342}; // @[Util.scala 113:33:@4740.4]
  assign _T_346 = {{1'd0}, _T_345}; // @[Util.scala 113:33:@4743.4]
  assign _T_349 = {{1'd0}, _T_348}; // @[Util.scala 113:33:@4746.4]
  assign _T_352 = {{1'd0}, _T_351}; // @[Util.scala 113:33:@4749.4]
  assign _T_355 = {{1'd0}, _T_354}; // @[Util.scala 113:33:@4752.4]
  assign _T_358 = {{1'd0}, _T_357}; // @[Util.scala 113:33:@4755.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 137:31:@4846.4]
  assign _T_446 = io_rw_cmd != 3'h0; // @[CSR.scala 138:27:@4847.4]
  assign _T_448 = system_insn == 1'h0; // @[CSR.scala 138:40:@4848.4]
  assign cpu_ren = _T_446 & _T_448; // @[CSR.scala 138:37:@4849.4]
  assign read_mstatus = {io_status_prv,io_status_unimp5,io_status_mprv,io_status_unimp4,io_status_mpp,io_status_unimp3,io_status_mpie,io_status_unimp2,io_status_mie,io_status_unimp1}; // @[CSR.scala 140:32:@4858.4]
  assign _T_468 = {5'h0,3'h0,reg_mip_mtip,3'h0,reg_mip_msip,3'h0}; // @[CSR.scala 156:25:@4864.4]
  assign _T_474 = {5'h0,3'h0,reg_mie_mtip,3'h0,reg_mie_msip,3'h0}; // @[CSR.scala 157:25:@4870.4]
  assign _T_478 = io_rw_addr == 12'hb00; // @[CSR.scala 177:73:@4871.4]
  assign _T_480 = io_rw_addr == 12'hb02; // @[CSR.scala 177:73:@4872.4]
  assign _T_482 = io_rw_addr == 12'hf13; // @[CSR.scala 177:73:@4873.4]
  assign _T_488 = io_rw_addr == 12'h301; // @[CSR.scala 177:73:@4876.4]
  assign _T_490 = io_rw_addr == 12'h300; // @[CSR.scala 177:73:@4877.4]
  assign _T_492 = io_rw_addr == 12'h305; // @[CSR.scala 177:73:@4878.4]
  assign _T_494 = io_rw_addr == 12'h344; // @[CSR.scala 177:73:@4879.4]
  assign _T_496 = io_rw_addr == 12'h304; // @[CSR.scala 177:73:@4880.4]
  assign _T_498 = io_rw_addr == 12'h340; // @[CSR.scala 177:73:@4881.4]
  assign _T_500 = io_rw_addr == 12'h341; // @[CSR.scala 177:73:@4882.4]
  assign _T_502 = io_rw_addr == 12'h343; // @[CSR.scala 177:73:@4883.4]
  assign _T_504 = io_rw_addr == 12'h342; // @[CSR.scala 177:73:@4884.4]
  assign _T_508 = io_rw_addr == 12'h7b2; // @[CSR.scala 177:73:@4886.4]
  assign _T_510 = io_rw_addr == 12'h302; // @[CSR.scala 177:73:@4887.4]
  assign _T_512 = io_rw_addr == 12'hb03; // @[CSR.scala 177:73:@4888.4]
  assign _T_514 = io_rw_addr == 12'hb83; // @[CSR.scala 177:73:@4889.4]
  assign _T_516 = io_rw_addr == 12'hb04; // @[CSR.scala 177:73:@4890.4]
  assign _T_518 = io_rw_addr == 12'hb84; // @[CSR.scala 177:73:@4891.4]
  assign _T_520 = io_rw_addr == 12'hb05; // @[CSR.scala 177:73:@4892.4]
  assign _T_522 = io_rw_addr == 12'hb85; // @[CSR.scala 177:73:@4893.4]
  assign _T_524 = io_rw_addr == 12'hb06; // @[CSR.scala 177:73:@4894.4]
  assign _T_526 = io_rw_addr == 12'hb86; // @[CSR.scala 177:73:@4895.4]
  assign _T_528 = io_rw_addr == 12'hb07; // @[CSR.scala 177:73:@4896.4]
  assign _T_530 = io_rw_addr == 12'hb87; // @[CSR.scala 177:73:@4897.4]
  assign _T_532 = io_rw_addr == 12'hb08; // @[CSR.scala 177:73:@4898.4]
  assign _T_534 = io_rw_addr == 12'hb88; // @[CSR.scala 177:73:@4899.4]
  assign _T_536 = io_rw_addr == 12'hb09; // @[CSR.scala 177:73:@4900.4]
  assign _T_538 = io_rw_addr == 12'hb89; // @[CSR.scala 177:73:@4901.4]
  assign _T_540 = io_rw_addr == 12'hb0a; // @[CSR.scala 177:73:@4902.4]
  assign _T_542 = io_rw_addr == 12'hb8a; // @[CSR.scala 177:73:@4903.4]
  assign _T_544 = io_rw_addr == 12'hb0b; // @[CSR.scala 177:73:@4904.4]
  assign _T_546 = io_rw_addr == 12'hb8b; // @[CSR.scala 177:73:@4905.4]
  assign _T_548 = io_rw_addr == 12'hb0c; // @[CSR.scala 177:73:@4906.4]
  assign _T_550 = io_rw_addr == 12'hb8c; // @[CSR.scala 177:73:@4907.4]
  assign _T_552 = io_rw_addr == 12'hb0d; // @[CSR.scala 177:73:@4908.4]
  assign _T_554 = io_rw_addr == 12'hb8d; // @[CSR.scala 177:73:@4909.4]
  assign _T_556 = io_rw_addr == 12'hb0e; // @[CSR.scala 177:73:@4910.4]
  assign _T_558 = io_rw_addr == 12'hb8e; // @[CSR.scala 177:73:@4911.4]
  assign _T_560 = io_rw_addr == 12'hb0f; // @[CSR.scala 177:73:@4912.4]
  assign _T_562 = io_rw_addr == 12'hb8f; // @[CSR.scala 177:73:@4913.4]
  assign _T_564 = io_rw_addr == 12'hb10; // @[CSR.scala 177:73:@4914.4]
  assign _T_566 = io_rw_addr == 12'hb90; // @[CSR.scala 177:73:@4915.4]
  assign _T_568 = io_rw_addr == 12'hb11; // @[CSR.scala 177:73:@4916.4]
  assign _T_570 = io_rw_addr == 12'hb91; // @[CSR.scala 177:73:@4917.4]
  assign _T_572 = io_rw_addr == 12'hb12; // @[CSR.scala 177:73:@4918.4]
  assign _T_574 = io_rw_addr == 12'hb92; // @[CSR.scala 177:73:@4919.4]
  assign _T_576 = io_rw_addr == 12'hb13; // @[CSR.scala 177:73:@4920.4]
  assign _T_578 = io_rw_addr == 12'hb93; // @[CSR.scala 177:73:@4921.4]
  assign _T_580 = io_rw_addr == 12'hb14; // @[CSR.scala 177:73:@4922.4]
  assign _T_582 = io_rw_addr == 12'hb94; // @[CSR.scala 177:73:@4923.4]
  assign _T_584 = io_rw_addr == 12'hb15; // @[CSR.scala 177:73:@4924.4]
  assign _T_586 = io_rw_addr == 12'hb95; // @[CSR.scala 177:73:@4925.4]
  assign _T_588 = io_rw_addr == 12'hb16; // @[CSR.scala 177:73:@4926.4]
  assign _T_590 = io_rw_addr == 12'hb96; // @[CSR.scala 177:73:@4927.4]
  assign _T_592 = io_rw_addr == 12'hb17; // @[CSR.scala 177:73:@4928.4]
  assign _T_594 = io_rw_addr == 12'hb97; // @[CSR.scala 177:73:@4929.4]
  assign _T_596 = io_rw_addr == 12'hb18; // @[CSR.scala 177:73:@4930.4]
  assign _T_598 = io_rw_addr == 12'hb98; // @[CSR.scala 177:73:@4931.4]
  assign _T_600 = io_rw_addr == 12'hb19; // @[CSR.scala 177:73:@4932.4]
  assign _T_602 = io_rw_addr == 12'hb99; // @[CSR.scala 177:73:@4933.4]
  assign _T_604 = io_rw_addr == 12'hb1a; // @[CSR.scala 177:73:@4934.4]
  assign _T_606 = io_rw_addr == 12'hb9a; // @[CSR.scala 177:73:@4935.4]
  assign _T_608 = io_rw_addr == 12'hb1b; // @[CSR.scala 177:73:@4936.4]
  assign _T_610 = io_rw_addr == 12'hb9b; // @[CSR.scala 177:73:@4937.4]
  assign _T_612 = io_rw_addr == 12'hb1c; // @[CSR.scala 177:73:@4938.4]
  assign _T_614 = io_rw_addr == 12'hb9c; // @[CSR.scala 177:73:@4939.4]
  assign _T_616 = io_rw_addr == 12'hb1d; // @[CSR.scala 177:73:@4940.4]
  assign _T_618 = io_rw_addr == 12'hb9d; // @[CSR.scala 177:73:@4941.4]
  assign _T_620 = io_rw_addr == 12'hb1e; // @[CSR.scala 177:73:@4942.4]
  assign _T_622 = io_rw_addr == 12'hb9e; // @[CSR.scala 177:73:@4943.4]
  assign _T_624 = io_rw_addr == 12'hb1f; // @[CSR.scala 177:73:@4944.4]
  assign _T_626 = io_rw_addr == 12'hb9f; // @[CSR.scala 177:73:@4945.4]
  assign _T_628 = io_rw_addr == 12'hb20; // @[CSR.scala 177:73:@4946.4]
  assign _T_630 = io_rw_addr == 12'hba0; // @[CSR.scala 177:73:@4947.4]
  assign _T_632 = io_rw_addr == 12'hb21; // @[CSR.scala 177:73:@4948.4]
  assign _T_634 = io_rw_addr == 12'hba1; // @[CSR.scala 177:73:@4949.4]
  assign _T_636 = io_rw_addr == 12'hb22; // @[CSR.scala 177:73:@4950.4]
  assign _T_638 = io_rw_addr == 12'hba2; // @[CSR.scala 177:73:@4951.4]
  assign _T_640 = io_rw_addr == 12'hb80; // @[CSR.scala 177:73:@4952.4]
  assign _T_642 = io_rw_addr == 12'hb82; // @[CSR.scala 177:73:@4953.4]
  assign _T_643 = io_rw_addr[9:8]; // @[CSR.scala 179:54:@4954.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_643; // @[CSR.scala 179:41:@4955.4]
  assign _T_644 = io_rw_addr[11:10]; // @[CSR.scala 180:29:@4956.4]
  assign _T_645 = ~ _T_644; // @[CSR.scala 180:37:@4957.4]
  assign read_only = _T_645 == 2'h0; // @[CSR.scala 180:37:@4958.4]
  assign _T_647 = io_rw_cmd != 3'h5; // @[CSR.scala 181:38:@4959.4]
  assign _T_648 = cpu_ren & _T_647; // @[CSR.scala 181:25:@4960.4]
  assign cpu_wen = _T_648 & priv_sufficient; // @[CSR.scala 181:48:@4961.4]
  assign _T_650 = read_only == 1'h0; // @[CSR.scala 182:24:@4962.4]
  assign wen = cpu_wen & _T_650; // @[CSR.scala 182:21:@4963.4]
  assign _T_651 = io_rw_cmd == 3'h2; // @[Util.scala 23:47:@4964.4]
  assign _T_652 = io_rw_cmd == 3'h3; // @[Util.scala 23:47:@4965.4]
  assign _T_653 = _T_651 | _T_652; // @[Util.scala 23:62:@4966.4]
  assign _T_655 = _T_653 ? io_rw_rdata : 32'h0; // @[CSR.scala 281:9:@4967.4]
  assign _T_656 = _T_655 | io_rw_wdata; // @[CSR.scala 281:49:@4968.4]
  assign _T_659 = _T_652 ? io_rw_wdata : 32'h0; // @[CSR.scala 281:64:@4970.4]
  assign _T_660 = ~ _T_659; // @[CSR.scala 281:60:@4971.4]
  assign wdata = _T_656 & _T_660; // @[CSR.scala 281:58:@4972.4]
  assign _T_662 = io_rw_addr[2:0]; // @[CSR.scala 185:33:@4973.4]
  assign opcode = 8'h1 << _T_662; // @[CSR.scala 185:20:@4974.4]
  assign _T_663 = opcode[0]; // @[CSR.scala 186:40:@4975.4]
  assign insn_call = system_insn & _T_663; // @[CSR.scala 186:31:@4976.4]
  assign _T_664 = opcode[1]; // @[CSR.scala 187:41:@4977.4]
  assign insn_break = system_insn & _T_664; // @[CSR.scala 187:32:@4978.4]
  assign _T_665 = opcode[2]; // @[CSR.scala 188:39:@4979.4]
  assign _T_666 = system_insn & _T_665; // @[CSR.scala 188:30:@4980.4]
  assign insn_ret = _T_666 & priv_sufficient; // @[CSR.scala 188:43:@4981.4]
  assign _T_940 = insn_call | insn_break; // @[CSR.scala 199:24:@5180.4]
  assign _T_942 = {{1'd0}, insn_ret}; // @[Bitwise.scala 48:55:@5183.4]
  assign _T_944 = _T_942 <= 2'h1; // @[CSR.scala 201:50:@5184.4]
  assign _T_946 = _T_944 | reset; // @[CSR.scala 201:9:@5186.4]
  assign _T_948 = _T_946 == 1'h0; // @[CSR.scala 201:9:@5187.4]
  assign _T_951 = io_rw_addr[10]; // @[CSR.scala 208:32:@5196.4]
  assign _T_953 = _T_951 == 1'h0; // @[CSR.scala 208:21:@5197.4]
  assign _T_954 = insn_ret & _T_953; // @[CSR.scala 208:18:@5198.4]
  assign _GEN_3 = _T_954 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 208:38:@5199.4]
  assign _GEN_4 = _T_954 ? 1'h1 : reg_mstatus_mpie; // @[CSR.scala 208:38:@5199.4]
  assign new_prv = _T_954 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 208:38:@5199.4]
  assign _GEN_148 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 218:35:@5207.6]
  assign _T_958 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@5207.6]
  assign _T_959 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@5208.6]
  assign _GEN_7 = insn_call ? 32'h80000004 : reg_mepc; // @[CSR.scala 216:18:@5205.4]
  assign _GEN_8 = insn_call ? {{28'd0}, _T_959} : reg_mcause; // @[CSR.scala 216:18:@5205.4]
  assign _GEN_9 = insn_call ? io_pc : reg_mepc; // @[CSR.scala 216:18:@5205.4]
  assign _GEN_10 = insn_break ? 32'h80000004 : _GEN_7; // @[CSR.scala 223:19:@5212.4]
  assign _GEN_11 = insn_break ? 32'h3 : _GEN_8; // @[CSR.scala 223:19:@5212.4]
  assign _GEN_12 = insn_break ? io_pc : _GEN_9; // @[CSR.scala 223:19:@5212.4]
  assign _GEN_14 = io_xcpt ? io_cause : _GEN_11; // @[CSR.scala 229:17:@5217.4]
  assign _GEN_15 = io_xcpt ? io_pc : _GEN_12; // @[CSR.scala 229:17:@5217.4]
  assign _GEN_16 = io_xcpt ? io_tval : reg_mtval; // @[CSR.scala 229:17:@5217.4]
  assign _T_965 = _T_478 ? _T_249 : 64'h0; // @[Mux.scala 19:72:@5225.4]
  assign _T_967 = _T_480 ? _T_261 : 64'h0; // @[Mux.scala 19:72:@5226.4]
  assign _T_969 = _T_482 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:@5227.4]
  assign _T_975 = _T_488 ? 31'h40000100 : 31'h0; // @[Mux.scala 19:72:@5230.4]
  assign _T_977 = _T_490 ? read_mstatus : 32'h0; // @[Mux.scala 19:72:@5231.4]
  assign _T_979 = _T_492 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:@5232.4]
  assign _T_981 = _T_494 ? _T_468 : 16'h0; // @[Mux.scala 19:72:@5233.4]
  assign _T_983 = _T_496 ? _T_474 : 16'h0; // @[Mux.scala 19:72:@5234.4]
  assign _T_985 = _T_498 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:@5235.4]
  assign _T_987 = _T_500 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:@5236.4]
  assign _T_989 = _T_502 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:@5237.4]
  assign _T_991 = _T_504 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:@5238.4]
  assign _T_995 = _T_508 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:@5240.4]
  assign _T_997 = _T_510 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:@5241.4]
  assign _T_999 = _T_512 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@5242.4]
  assign _T_1001 = _T_514 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@5243.4]
  assign _T_1003 = _T_516 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@5244.4]
  assign _T_1005 = _T_518 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@5245.4]
  assign _T_1007 = _T_520 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@5246.4]
  assign _T_1009 = _T_522 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@5247.4]
  assign _T_1011 = _T_524 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@5248.4]
  assign _T_1013 = _T_526 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@5249.4]
  assign _T_1015 = _T_528 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@5250.4]
  assign _T_1017 = _T_530 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@5251.4]
  assign _T_1019 = _T_532 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@5252.4]
  assign _T_1021 = _T_534 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@5253.4]
  assign _T_1023 = _T_536 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@5254.4]
  assign _T_1025 = _T_538 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@5255.4]
  assign _T_1027 = _T_540 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@5256.4]
  assign _T_1029 = _T_542 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@5257.4]
  assign _T_1031 = _T_544 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@5258.4]
  assign _T_1033 = _T_546 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@5259.4]
  assign _T_1035 = _T_548 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@5260.4]
  assign _T_1037 = _T_550 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@5261.4]
  assign _T_1039 = _T_552 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@5262.4]
  assign _T_1041 = _T_554 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@5263.4]
  assign _T_1043 = _T_556 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@5264.4]
  assign _T_1045 = _T_558 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@5265.4]
  assign _T_1047 = _T_560 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@5266.4]
  assign _T_1049 = _T_562 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@5267.4]
  assign _T_1051 = _T_564 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@5268.4]
  assign _T_1053 = _T_566 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@5269.4]
  assign _T_1055 = _T_568 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@5270.4]
  assign _T_1057 = _T_570 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@5271.4]
  assign _T_1059 = _T_572 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@5272.4]
  assign _T_1061 = _T_574 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@5273.4]
  assign _T_1063 = _T_576 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@5274.4]
  assign _T_1065 = _T_578 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@5275.4]
  assign _T_1067 = _T_580 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@5276.4]
  assign _T_1069 = _T_582 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@5277.4]
  assign _T_1071 = _T_584 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@5278.4]
  assign _T_1073 = _T_586 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@5279.4]
  assign _T_1075 = _T_588 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@5280.4]
  assign _T_1077 = _T_590 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@5281.4]
  assign _T_1079 = _T_592 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@5282.4]
  assign _T_1081 = _T_594 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@5283.4]
  assign _T_1083 = _T_596 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@5284.4]
  assign _T_1085 = _T_598 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@5285.4]
  assign _T_1087 = _T_600 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@5286.4]
  assign _T_1089 = _T_602 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@5287.4]
  assign _T_1091 = _T_604 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@5288.4]
  assign _T_1093 = _T_606 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@5289.4]
  assign _T_1095 = _T_608 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@5290.4]
  assign _T_1097 = _T_610 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@5291.4]
  assign _T_1099 = _T_612 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@5292.4]
  assign _T_1101 = _T_614 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@5293.4]
  assign _T_1103 = _T_616 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@5294.4]
  assign _T_1105 = _T_618 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@5295.4]
  assign _T_1107 = _T_620 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@5296.4]
  assign _T_1109 = _T_622 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@5297.4]
  assign _T_1111 = _T_624 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@5298.4]
  assign _T_1113 = _T_626 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@5299.4]
  assign _T_1115 = _T_628 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@5300.4]
  assign _T_1117 = _T_630 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@5301.4]
  assign _T_1119 = _T_632 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@5302.4]
  assign _T_1121 = _T_634 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@5303.4]
  assign _T_1123 = _T_636 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@5304.4]
  assign _T_1125 = _T_638 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@5305.4]
  assign _T_1130 = _T_965 | _T_967; // @[Mux.scala 19:72:@5308.4]
  assign _GEN_149 = {{48'd0}, _T_969}; // @[Mux.scala 19:72:@5309.4]
  assign _T_1131 = _T_1130 | _GEN_149; // @[Mux.scala 19:72:@5309.4]
  assign _GEN_150 = {{33'd0}, _T_975}; // @[Mux.scala 19:72:@5312.4]
  assign _T_1134 = _T_1131 | _GEN_150; // @[Mux.scala 19:72:@5312.4]
  assign _GEN_151 = {{32'd0}, _T_977}; // @[Mux.scala 19:72:@5313.4]
  assign _T_1135 = _T_1134 | _GEN_151; // @[Mux.scala 19:72:@5313.4]
  assign _GEN_152 = {{55'd0}, _T_979}; // @[Mux.scala 19:72:@5314.4]
  assign _T_1136 = _T_1135 | _GEN_152; // @[Mux.scala 19:72:@5314.4]
  assign _GEN_153 = {{48'd0}, _T_981}; // @[Mux.scala 19:72:@5315.4]
  assign _T_1137 = _T_1136 | _GEN_153; // @[Mux.scala 19:72:@5315.4]
  assign _GEN_154 = {{48'd0}, _T_983}; // @[Mux.scala 19:72:@5316.4]
  assign _T_1138 = _T_1137 | _GEN_154; // @[Mux.scala 19:72:@5316.4]
  assign _GEN_155 = {{32'd0}, _T_985}; // @[Mux.scala 19:72:@5317.4]
  assign _T_1139 = _T_1138 | _GEN_155; // @[Mux.scala 19:72:@5317.4]
  assign _GEN_156 = {{32'd0}, _T_987}; // @[Mux.scala 19:72:@5318.4]
  assign _T_1140 = _T_1139 | _GEN_156; // @[Mux.scala 19:72:@5318.4]
  assign _GEN_157 = {{32'd0}, _T_989}; // @[Mux.scala 19:72:@5319.4]
  assign _T_1141 = _T_1140 | _GEN_157; // @[Mux.scala 19:72:@5319.4]
  assign _GEN_158 = {{32'd0}, _T_991}; // @[Mux.scala 19:72:@5320.4]
  assign _T_1142 = _T_1141 | _GEN_158; // @[Mux.scala 19:72:@5320.4]
  assign _GEN_159 = {{32'd0}, _T_995}; // @[Mux.scala 19:72:@5322.4]
  assign _T_1144 = _T_1142 | _GEN_159; // @[Mux.scala 19:72:@5322.4]
  assign _GEN_160 = {{32'd0}, _T_997}; // @[Mux.scala 19:72:@5323.4]
  assign _T_1145 = _T_1144 | _GEN_160; // @[Mux.scala 19:72:@5323.4]
  assign _GEN_161 = {{24'd0}, _T_999}; // @[Mux.scala 19:72:@5324.4]
  assign _T_1146 = _T_1145 | _GEN_161; // @[Mux.scala 19:72:@5324.4]
  assign _GEN_162 = {{24'd0}, _T_1001}; // @[Mux.scala 19:72:@5325.4]
  assign _T_1147 = _T_1146 | _GEN_162; // @[Mux.scala 19:72:@5325.4]
  assign _GEN_163 = {{24'd0}, _T_1003}; // @[Mux.scala 19:72:@5326.4]
  assign _T_1148 = _T_1147 | _GEN_163; // @[Mux.scala 19:72:@5326.4]
  assign _GEN_164 = {{24'd0}, _T_1005}; // @[Mux.scala 19:72:@5327.4]
  assign _T_1149 = _T_1148 | _GEN_164; // @[Mux.scala 19:72:@5327.4]
  assign _GEN_165 = {{24'd0}, _T_1007}; // @[Mux.scala 19:72:@5328.4]
  assign _T_1150 = _T_1149 | _GEN_165; // @[Mux.scala 19:72:@5328.4]
  assign _GEN_166 = {{24'd0}, _T_1009}; // @[Mux.scala 19:72:@5329.4]
  assign _T_1151 = _T_1150 | _GEN_166; // @[Mux.scala 19:72:@5329.4]
  assign _GEN_167 = {{24'd0}, _T_1011}; // @[Mux.scala 19:72:@5330.4]
  assign _T_1152 = _T_1151 | _GEN_167; // @[Mux.scala 19:72:@5330.4]
  assign _GEN_168 = {{24'd0}, _T_1013}; // @[Mux.scala 19:72:@5331.4]
  assign _T_1153 = _T_1152 | _GEN_168; // @[Mux.scala 19:72:@5331.4]
  assign _GEN_169 = {{24'd0}, _T_1015}; // @[Mux.scala 19:72:@5332.4]
  assign _T_1154 = _T_1153 | _GEN_169; // @[Mux.scala 19:72:@5332.4]
  assign _GEN_170 = {{24'd0}, _T_1017}; // @[Mux.scala 19:72:@5333.4]
  assign _T_1155 = _T_1154 | _GEN_170; // @[Mux.scala 19:72:@5333.4]
  assign _GEN_171 = {{24'd0}, _T_1019}; // @[Mux.scala 19:72:@5334.4]
  assign _T_1156 = _T_1155 | _GEN_171; // @[Mux.scala 19:72:@5334.4]
  assign _GEN_172 = {{24'd0}, _T_1021}; // @[Mux.scala 19:72:@5335.4]
  assign _T_1157 = _T_1156 | _GEN_172; // @[Mux.scala 19:72:@5335.4]
  assign _GEN_173 = {{24'd0}, _T_1023}; // @[Mux.scala 19:72:@5336.4]
  assign _T_1158 = _T_1157 | _GEN_173; // @[Mux.scala 19:72:@5336.4]
  assign _GEN_174 = {{24'd0}, _T_1025}; // @[Mux.scala 19:72:@5337.4]
  assign _T_1159 = _T_1158 | _GEN_174; // @[Mux.scala 19:72:@5337.4]
  assign _GEN_175 = {{24'd0}, _T_1027}; // @[Mux.scala 19:72:@5338.4]
  assign _T_1160 = _T_1159 | _GEN_175; // @[Mux.scala 19:72:@5338.4]
  assign _GEN_176 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:@5339.4]
  assign _T_1161 = _T_1160 | _GEN_176; // @[Mux.scala 19:72:@5339.4]
  assign _GEN_177 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:@5340.4]
  assign _T_1162 = _T_1161 | _GEN_177; // @[Mux.scala 19:72:@5340.4]
  assign _GEN_178 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:@5341.4]
  assign _T_1163 = _T_1162 | _GEN_178; // @[Mux.scala 19:72:@5341.4]
  assign _GEN_179 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:@5342.4]
  assign _T_1164 = _T_1163 | _GEN_179; // @[Mux.scala 19:72:@5342.4]
  assign _GEN_180 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:@5343.4]
  assign _T_1165 = _T_1164 | _GEN_180; // @[Mux.scala 19:72:@5343.4]
  assign _GEN_181 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:@5344.4]
  assign _T_1166 = _T_1165 | _GEN_181; // @[Mux.scala 19:72:@5344.4]
  assign _GEN_182 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:@5345.4]
  assign _T_1167 = _T_1166 | _GEN_182; // @[Mux.scala 19:72:@5345.4]
  assign _GEN_183 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:@5346.4]
  assign _T_1168 = _T_1167 | _GEN_183; // @[Mux.scala 19:72:@5346.4]
  assign _GEN_184 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:@5347.4]
  assign _T_1169 = _T_1168 | _GEN_184; // @[Mux.scala 19:72:@5347.4]
  assign _GEN_185 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:@5348.4]
  assign _T_1170 = _T_1169 | _GEN_185; // @[Mux.scala 19:72:@5348.4]
  assign _GEN_186 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:@5349.4]
  assign _T_1171 = _T_1170 | _GEN_186; // @[Mux.scala 19:72:@5349.4]
  assign _GEN_187 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:@5350.4]
  assign _T_1172 = _T_1171 | _GEN_187; // @[Mux.scala 19:72:@5350.4]
  assign _GEN_188 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:@5351.4]
  assign _T_1173 = _T_1172 | _GEN_188; // @[Mux.scala 19:72:@5351.4]
  assign _GEN_189 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:@5352.4]
  assign _T_1174 = _T_1173 | _GEN_189; // @[Mux.scala 19:72:@5352.4]
  assign _GEN_190 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:@5353.4]
  assign _T_1175 = _T_1174 | _GEN_190; // @[Mux.scala 19:72:@5353.4]
  assign _GEN_191 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:@5354.4]
  assign _T_1176 = _T_1175 | _GEN_191; // @[Mux.scala 19:72:@5354.4]
  assign _GEN_192 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:@5355.4]
  assign _T_1177 = _T_1176 | _GEN_192; // @[Mux.scala 19:72:@5355.4]
  assign _GEN_193 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:@5356.4]
  assign _T_1178 = _T_1177 | _GEN_193; // @[Mux.scala 19:72:@5356.4]
  assign _GEN_194 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:@5357.4]
  assign _T_1179 = _T_1178 | _GEN_194; // @[Mux.scala 19:72:@5357.4]
  assign _GEN_195 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:@5358.4]
  assign _T_1180 = _T_1179 | _GEN_195; // @[Mux.scala 19:72:@5358.4]
  assign _GEN_196 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:@5359.4]
  assign _T_1181 = _T_1180 | _GEN_196; // @[Mux.scala 19:72:@5359.4]
  assign _GEN_197 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:@5360.4]
  assign _T_1182 = _T_1181 | _GEN_197; // @[Mux.scala 19:72:@5360.4]
  assign _GEN_198 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:@5361.4]
  assign _T_1183 = _T_1182 | _GEN_198; // @[Mux.scala 19:72:@5361.4]
  assign _GEN_199 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:@5362.4]
  assign _T_1184 = _T_1183 | _GEN_199; // @[Mux.scala 19:72:@5362.4]
  assign _GEN_200 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:@5363.4]
  assign _T_1185 = _T_1184 | _GEN_200; // @[Mux.scala 19:72:@5363.4]
  assign _GEN_201 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:@5364.4]
  assign _T_1186 = _T_1185 | _GEN_201; // @[Mux.scala 19:72:@5364.4]
  assign _GEN_202 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:@5365.4]
  assign _T_1187 = _T_1186 | _GEN_202; // @[Mux.scala 19:72:@5365.4]
  assign _GEN_203 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:@5366.4]
  assign _T_1188 = _T_1187 | _GEN_203; // @[Mux.scala 19:72:@5366.4]
  assign _GEN_204 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:@5367.4]
  assign _T_1189 = _T_1188 | _GEN_204; // @[Mux.scala 19:72:@5367.4]
  assign _GEN_205 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:@5368.4]
  assign _T_1190 = _T_1189 | _GEN_205; // @[Mux.scala 19:72:@5368.4]
  assign _GEN_206 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:@5369.4]
  assign _T_1191 = _T_1190 | _GEN_206; // @[Mux.scala 19:72:@5369.4]
  assign _GEN_207 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:@5370.4]
  assign _T_1192 = _T_1191 | _GEN_207; // @[Mux.scala 19:72:@5370.4]
  assign _GEN_208 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:@5371.4]
  assign _T_1193 = _T_1192 | _GEN_208; // @[Mux.scala 19:72:@5371.4]
  assign _GEN_209 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:@5372.4]
  assign _T_1194 = _T_1193 | _GEN_209; // @[Mux.scala 19:72:@5372.4]
  assign _GEN_210 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:@5373.4]
  assign _T_1195 = _T_1194 | _GEN_210; // @[Mux.scala 19:72:@5373.4]
  assign _GEN_211 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:@5374.4]
  assign _T_1196 = _T_1195 | _GEN_211; // @[Mux.scala 19:72:@5374.4]
  assign _GEN_212 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:@5375.4]
  assign _T_1197 = _T_1196 | _GEN_212; // @[Mux.scala 19:72:@5375.4]
  assign _GEN_213 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:@5376.4]
  assign _T_1198 = _T_1197 | _GEN_213; // @[Mux.scala 19:72:@5376.4]
  assign _GEN_214 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:@5377.4]
  assign _T_1199 = _T_1198 | _GEN_214; // @[Mux.scala 19:72:@5377.4]
  assign _GEN_215 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:@5378.4]
  assign _T_1200 = _T_1199 | _GEN_215; // @[Mux.scala 19:72:@5378.4]
  assign _GEN_216 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:@5379.4]
  assign _T_1201 = _T_1200 | _GEN_216; // @[Mux.scala 19:72:@5379.4]
  assign _GEN_217 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:@5380.4]
  assign _T_1202 = _T_1201 | _GEN_217; // @[Mux.scala 19:72:@5380.4]
  assign _GEN_218 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:@5381.4]
  assign _T_1203 = _T_1202 | _GEN_218; // @[Mux.scala 19:72:@5381.4]
  assign _GEN_219 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:@5382.4]
  assign _T_1204 = _T_1203 | _GEN_219; // @[Mux.scala 19:72:@5382.4]
  assign _GEN_220 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:@5383.4]
  assign _T_1205 = _T_1204 | _GEN_220; // @[Mux.scala 19:72:@5383.4]
  assign _GEN_221 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:@5384.4]
  assign _T_1206 = _T_1205 | _GEN_221; // @[Mux.scala 19:72:@5384.4]
  assign _GEN_222 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:@5385.4]
  assign _T_1207 = _T_1206 | _GEN_222; // @[Mux.scala 19:72:@5385.4]
  assign _GEN_223 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:@5386.4]
  assign _T_1208 = _T_1207 | _GEN_223; // @[Mux.scala 19:72:@5386.4]
  assign _GEN_224 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:@5387.4]
  assign _T_1209 = _T_1208 | _GEN_224; // @[Mux.scala 19:72:@5387.4]
  assign _T_1220 = wdata[3]; // @[CSR.scala 245:39:@5400.8]
  assign _T_1222 = wdata[7]; // @[CSR.scala 245:39:@5404.8]
  assign _GEN_17 = _T_490 ? _T_1220 : _GEN_3; // @[CSR.scala 244:39:@5394.6]
  assign _GEN_18 = _T_490 ? _T_1222 : _GEN_4; // @[CSR.scala 244:39:@5394.6]
  assign _T_1233 = wdata[15:0]; // @[:@5423.8 :@5424.8]
  assign _T_1235 = _T_1233[3]; // @[CSR.scala 250:35:@5427.8]
  assign _T_1237 = _T_1233[7]; // @[CSR.scala 250:35:@5431.8]
  assign _GEN_19 = _T_494 ? _T_1235 : reg_mip_msip; // @[CSR.scala 249:35:@5421.6]
  assign _GEN_20 = _T_496 ? _T_1235 : reg_mie_msip; // @[CSR.scala 253:35:@5441.6]
  assign _GEN_21 = _T_496 ? _T_1237 : reg_mie_mtip; // @[CSR.scala 253:35:@5441.6]
  assign _T_1253 = wdata[7:0]; // @[CSR.scala 277:47:@5463.8]
  assign _T_1254 = _T_264[31:0]; // @[CSR.scala 277:72:@5464.8]
  assign _T_1255 = {_T_1253,_T_1254}; // @[Cat.scala 30:58:@5465.8]
  assign _GEN_22 = _T_514 ? {{1'd0}, _T_1255} : _T_265; // @[CSR.scala 277:29:@5462.6]
  assign _T_1256 = _T_264[39:32]; // @[CSR.scala 278:45:@5469.8]
  assign _T_1257 = {_T_1256,wdata}; // @[Cat.scala 30:58:@5470.8]
  assign _GEN_23 = _T_512 ? {{1'd0}, _T_1257} : _GEN_22; // @[CSR.scala 278:29:@5468.6]
  assign _T_1259 = _T_267[31:0]; // @[CSR.scala 277:72:@5475.8]
  assign _T_1260 = {_T_1253,_T_1259}; // @[Cat.scala 30:58:@5476.8]
  assign _GEN_24 = _T_518 ? {{1'd0}, _T_1260} : _T_268; // @[CSR.scala 277:29:@5473.6]
  assign _T_1261 = _T_267[39:32]; // @[CSR.scala 278:45:@5480.8]
  assign _T_1262 = {_T_1261,wdata}; // @[Cat.scala 30:58:@5481.8]
  assign _GEN_25 = _T_516 ? {{1'd0}, _T_1262} : _GEN_24; // @[CSR.scala 278:29:@5479.6]
  assign _T_1264 = _T_270[31:0]; // @[CSR.scala 277:72:@5486.8]
  assign _T_1265 = {_T_1253,_T_1264}; // @[Cat.scala 30:58:@5487.8]
  assign _GEN_26 = _T_522 ? {{1'd0}, _T_1265} : _T_271; // @[CSR.scala 277:29:@5484.6]
  assign _T_1266 = _T_270[39:32]; // @[CSR.scala 278:45:@5491.8]
  assign _T_1267 = {_T_1266,wdata}; // @[Cat.scala 30:58:@5492.8]
  assign _GEN_27 = _T_520 ? {{1'd0}, _T_1267} : _GEN_26; // @[CSR.scala 278:29:@5490.6]
  assign _T_1269 = _T_273[31:0]; // @[CSR.scala 277:72:@5497.8]
  assign _T_1270 = {_T_1253,_T_1269}; // @[Cat.scala 30:58:@5498.8]
  assign _GEN_28 = _T_526 ? {{1'd0}, _T_1270} : _T_274; // @[CSR.scala 277:29:@5495.6]
  assign _T_1271 = _T_273[39:32]; // @[CSR.scala 278:45:@5502.8]
  assign _T_1272 = {_T_1271,wdata}; // @[Cat.scala 30:58:@5503.8]
  assign _GEN_29 = _T_524 ? {{1'd0}, _T_1272} : _GEN_28; // @[CSR.scala 278:29:@5501.6]
  assign _T_1274 = _T_276[31:0]; // @[CSR.scala 277:72:@5508.8]
  assign _T_1275 = {_T_1253,_T_1274}; // @[Cat.scala 30:58:@5509.8]
  assign _GEN_30 = _T_530 ? {{1'd0}, _T_1275} : _T_277; // @[CSR.scala 277:29:@5506.6]
  assign _T_1276 = _T_276[39:32]; // @[CSR.scala 278:45:@5513.8]
  assign _T_1277 = {_T_1276,wdata}; // @[Cat.scala 30:58:@5514.8]
  assign _GEN_31 = _T_528 ? {{1'd0}, _T_1277} : _GEN_30; // @[CSR.scala 278:29:@5512.6]
  assign _T_1279 = _T_279[31:0]; // @[CSR.scala 277:72:@5519.8]
  assign _T_1280 = {_T_1253,_T_1279}; // @[Cat.scala 30:58:@5520.8]
  assign _GEN_32 = _T_534 ? {{1'd0}, _T_1280} : _T_280; // @[CSR.scala 277:29:@5517.6]
  assign _T_1281 = _T_279[39:32]; // @[CSR.scala 278:45:@5524.8]
  assign _T_1282 = {_T_1281,wdata}; // @[Cat.scala 30:58:@5525.8]
  assign _GEN_33 = _T_532 ? {{1'd0}, _T_1282} : _GEN_32; // @[CSR.scala 278:29:@5523.6]
  assign _T_1284 = _T_282[31:0]; // @[CSR.scala 277:72:@5530.8]
  assign _T_1285 = {_T_1253,_T_1284}; // @[Cat.scala 30:58:@5531.8]
  assign _GEN_34 = _T_538 ? {{1'd0}, _T_1285} : _T_283; // @[CSR.scala 277:29:@5528.6]
  assign _T_1286 = _T_282[39:32]; // @[CSR.scala 278:45:@5535.8]
  assign _T_1287 = {_T_1286,wdata}; // @[Cat.scala 30:58:@5536.8]
  assign _GEN_35 = _T_536 ? {{1'd0}, _T_1287} : _GEN_34; // @[CSR.scala 278:29:@5534.6]
  assign _T_1289 = _T_285[31:0]; // @[CSR.scala 277:72:@5541.8]
  assign _T_1290 = {_T_1253,_T_1289}; // @[Cat.scala 30:58:@5542.8]
  assign _GEN_36 = _T_542 ? {{1'd0}, _T_1290} : _T_286; // @[CSR.scala 277:29:@5539.6]
  assign _T_1291 = _T_285[39:32]; // @[CSR.scala 278:45:@5546.8]
  assign _T_1292 = {_T_1291,wdata}; // @[Cat.scala 30:58:@5547.8]
  assign _GEN_37 = _T_540 ? {{1'd0}, _T_1292} : _GEN_36; // @[CSR.scala 278:29:@5545.6]
  assign _T_1294 = _T_288[31:0]; // @[CSR.scala 277:72:@5552.8]
  assign _T_1295 = {_T_1253,_T_1294}; // @[Cat.scala 30:58:@5553.8]
  assign _GEN_38 = _T_546 ? {{1'd0}, _T_1295} : _T_289; // @[CSR.scala 277:29:@5550.6]
  assign _T_1296 = _T_288[39:32]; // @[CSR.scala 278:45:@5557.8]
  assign _T_1297 = {_T_1296,wdata}; // @[Cat.scala 30:58:@5558.8]
  assign _GEN_39 = _T_544 ? {{1'd0}, _T_1297} : _GEN_38; // @[CSR.scala 278:29:@5556.6]
  assign _T_1299 = _T_291[31:0]; // @[CSR.scala 277:72:@5563.8]
  assign _T_1300 = {_T_1253,_T_1299}; // @[Cat.scala 30:58:@5564.8]
  assign _GEN_40 = _T_550 ? {{1'd0}, _T_1300} : _T_292; // @[CSR.scala 277:29:@5561.6]
  assign _T_1301 = _T_291[39:32]; // @[CSR.scala 278:45:@5568.8]
  assign _T_1302 = {_T_1301,wdata}; // @[Cat.scala 30:58:@5569.8]
  assign _GEN_41 = _T_548 ? {{1'd0}, _T_1302} : _GEN_40; // @[CSR.scala 278:29:@5567.6]
  assign _T_1304 = _T_294[31:0]; // @[CSR.scala 277:72:@5574.8]
  assign _T_1305 = {_T_1253,_T_1304}; // @[Cat.scala 30:58:@5575.8]
  assign _GEN_42 = _T_554 ? {{1'd0}, _T_1305} : _T_295; // @[CSR.scala 277:29:@5572.6]
  assign _T_1306 = _T_294[39:32]; // @[CSR.scala 278:45:@5579.8]
  assign _T_1307 = {_T_1306,wdata}; // @[Cat.scala 30:58:@5580.8]
  assign _GEN_43 = _T_552 ? {{1'd0}, _T_1307} : _GEN_42; // @[CSR.scala 278:29:@5578.6]
  assign _T_1309 = _T_297[31:0]; // @[CSR.scala 277:72:@5585.8]
  assign _T_1310 = {_T_1253,_T_1309}; // @[Cat.scala 30:58:@5586.8]
  assign _GEN_44 = _T_558 ? {{1'd0}, _T_1310} : _T_298; // @[CSR.scala 277:29:@5583.6]
  assign _T_1311 = _T_297[39:32]; // @[CSR.scala 278:45:@5590.8]
  assign _T_1312 = {_T_1311,wdata}; // @[Cat.scala 30:58:@5591.8]
  assign _GEN_45 = _T_556 ? {{1'd0}, _T_1312} : _GEN_44; // @[CSR.scala 278:29:@5589.6]
  assign _T_1314 = _T_300[31:0]; // @[CSR.scala 277:72:@5596.8]
  assign _T_1315 = {_T_1253,_T_1314}; // @[Cat.scala 30:58:@5597.8]
  assign _GEN_46 = _T_562 ? {{1'd0}, _T_1315} : _T_301; // @[CSR.scala 277:29:@5594.6]
  assign _T_1316 = _T_300[39:32]; // @[CSR.scala 278:45:@5601.8]
  assign _T_1317 = {_T_1316,wdata}; // @[Cat.scala 30:58:@5602.8]
  assign _GEN_47 = _T_560 ? {{1'd0}, _T_1317} : _GEN_46; // @[CSR.scala 278:29:@5600.6]
  assign _T_1319 = _T_303[31:0]; // @[CSR.scala 277:72:@5607.8]
  assign _T_1320 = {_T_1253,_T_1319}; // @[Cat.scala 30:58:@5608.8]
  assign _GEN_48 = _T_566 ? {{1'd0}, _T_1320} : _T_304; // @[CSR.scala 277:29:@5605.6]
  assign _T_1321 = _T_303[39:32]; // @[CSR.scala 278:45:@5612.8]
  assign _T_1322 = {_T_1321,wdata}; // @[Cat.scala 30:58:@5613.8]
  assign _GEN_49 = _T_564 ? {{1'd0}, _T_1322} : _GEN_48; // @[CSR.scala 278:29:@5611.6]
  assign _T_1324 = _T_306[31:0]; // @[CSR.scala 277:72:@5618.8]
  assign _T_1325 = {_T_1253,_T_1324}; // @[Cat.scala 30:58:@5619.8]
  assign _GEN_50 = _T_570 ? {{1'd0}, _T_1325} : _T_307; // @[CSR.scala 277:29:@5616.6]
  assign _T_1326 = _T_306[39:32]; // @[CSR.scala 278:45:@5623.8]
  assign _T_1327 = {_T_1326,wdata}; // @[Cat.scala 30:58:@5624.8]
  assign _GEN_51 = _T_568 ? {{1'd0}, _T_1327} : _GEN_50; // @[CSR.scala 278:29:@5622.6]
  assign _T_1329 = _T_309[31:0]; // @[CSR.scala 277:72:@5629.8]
  assign _T_1330 = {_T_1253,_T_1329}; // @[Cat.scala 30:58:@5630.8]
  assign _GEN_52 = _T_574 ? {{1'd0}, _T_1330} : _T_310; // @[CSR.scala 277:29:@5627.6]
  assign _T_1331 = _T_309[39:32]; // @[CSR.scala 278:45:@5634.8]
  assign _T_1332 = {_T_1331,wdata}; // @[Cat.scala 30:58:@5635.8]
  assign _GEN_53 = _T_572 ? {{1'd0}, _T_1332} : _GEN_52; // @[CSR.scala 278:29:@5633.6]
  assign _T_1334 = _T_312[31:0]; // @[CSR.scala 277:72:@5640.8]
  assign _T_1335 = {_T_1253,_T_1334}; // @[Cat.scala 30:58:@5641.8]
  assign _GEN_54 = _T_578 ? {{1'd0}, _T_1335} : _T_313; // @[CSR.scala 277:29:@5638.6]
  assign _T_1336 = _T_312[39:32]; // @[CSR.scala 278:45:@5645.8]
  assign _T_1337 = {_T_1336,wdata}; // @[Cat.scala 30:58:@5646.8]
  assign _GEN_55 = _T_576 ? {{1'd0}, _T_1337} : _GEN_54; // @[CSR.scala 278:29:@5644.6]
  assign _T_1339 = _T_315[31:0]; // @[CSR.scala 277:72:@5651.8]
  assign _T_1340 = {_T_1253,_T_1339}; // @[Cat.scala 30:58:@5652.8]
  assign _GEN_56 = _T_582 ? {{1'd0}, _T_1340} : _T_316; // @[CSR.scala 277:29:@5649.6]
  assign _T_1341 = _T_315[39:32]; // @[CSR.scala 278:45:@5656.8]
  assign _T_1342 = {_T_1341,wdata}; // @[Cat.scala 30:58:@5657.8]
  assign _GEN_57 = _T_580 ? {{1'd0}, _T_1342} : _GEN_56; // @[CSR.scala 278:29:@5655.6]
  assign _T_1344 = _T_318[31:0]; // @[CSR.scala 277:72:@5662.8]
  assign _T_1345 = {_T_1253,_T_1344}; // @[Cat.scala 30:58:@5663.8]
  assign _GEN_58 = _T_586 ? {{1'd0}, _T_1345} : _T_319; // @[CSR.scala 277:29:@5660.6]
  assign _T_1346 = _T_318[39:32]; // @[CSR.scala 278:45:@5667.8]
  assign _T_1347 = {_T_1346,wdata}; // @[Cat.scala 30:58:@5668.8]
  assign _GEN_59 = _T_584 ? {{1'd0}, _T_1347} : _GEN_58; // @[CSR.scala 278:29:@5666.6]
  assign _T_1349 = _T_321[31:0]; // @[CSR.scala 277:72:@5673.8]
  assign _T_1350 = {_T_1253,_T_1349}; // @[Cat.scala 30:58:@5674.8]
  assign _GEN_60 = _T_590 ? {{1'd0}, _T_1350} : _T_322; // @[CSR.scala 277:29:@5671.6]
  assign _T_1351 = _T_321[39:32]; // @[CSR.scala 278:45:@5678.8]
  assign _T_1352 = {_T_1351,wdata}; // @[Cat.scala 30:58:@5679.8]
  assign _GEN_61 = _T_588 ? {{1'd0}, _T_1352} : _GEN_60; // @[CSR.scala 278:29:@5677.6]
  assign _T_1354 = _T_324[31:0]; // @[CSR.scala 277:72:@5684.8]
  assign _T_1355 = {_T_1253,_T_1354}; // @[Cat.scala 30:58:@5685.8]
  assign _GEN_62 = _T_594 ? {{1'd0}, _T_1355} : _T_325; // @[CSR.scala 277:29:@5682.6]
  assign _T_1356 = _T_324[39:32]; // @[CSR.scala 278:45:@5689.8]
  assign _T_1357 = {_T_1356,wdata}; // @[Cat.scala 30:58:@5690.8]
  assign _GEN_63 = _T_592 ? {{1'd0}, _T_1357} : _GEN_62; // @[CSR.scala 278:29:@5688.6]
  assign _T_1359 = _T_327[31:0]; // @[CSR.scala 277:72:@5695.8]
  assign _T_1360 = {_T_1253,_T_1359}; // @[Cat.scala 30:58:@5696.8]
  assign _GEN_64 = _T_598 ? {{1'd0}, _T_1360} : _T_328; // @[CSR.scala 277:29:@5693.6]
  assign _T_1361 = _T_327[39:32]; // @[CSR.scala 278:45:@5700.8]
  assign _T_1362 = {_T_1361,wdata}; // @[Cat.scala 30:58:@5701.8]
  assign _GEN_65 = _T_596 ? {{1'd0}, _T_1362} : _GEN_64; // @[CSR.scala 278:29:@5699.6]
  assign _T_1364 = _T_330[31:0]; // @[CSR.scala 277:72:@5706.8]
  assign _T_1365 = {_T_1253,_T_1364}; // @[Cat.scala 30:58:@5707.8]
  assign _GEN_66 = _T_602 ? {{1'd0}, _T_1365} : _T_331; // @[CSR.scala 277:29:@5704.6]
  assign _T_1366 = _T_330[39:32]; // @[CSR.scala 278:45:@5711.8]
  assign _T_1367 = {_T_1366,wdata}; // @[Cat.scala 30:58:@5712.8]
  assign _GEN_67 = _T_600 ? {{1'd0}, _T_1367} : _GEN_66; // @[CSR.scala 278:29:@5710.6]
  assign _T_1369 = _T_333[31:0]; // @[CSR.scala 277:72:@5717.8]
  assign _T_1370 = {_T_1253,_T_1369}; // @[Cat.scala 30:58:@5718.8]
  assign _GEN_68 = _T_606 ? {{1'd0}, _T_1370} : _T_334; // @[CSR.scala 277:29:@5715.6]
  assign _T_1371 = _T_333[39:32]; // @[CSR.scala 278:45:@5722.8]
  assign _T_1372 = {_T_1371,wdata}; // @[Cat.scala 30:58:@5723.8]
  assign _GEN_69 = _T_604 ? {{1'd0}, _T_1372} : _GEN_68; // @[CSR.scala 278:29:@5721.6]
  assign _T_1374 = _T_336[31:0]; // @[CSR.scala 277:72:@5728.8]
  assign _T_1375 = {_T_1253,_T_1374}; // @[Cat.scala 30:58:@5729.8]
  assign _GEN_70 = _T_610 ? {{1'd0}, _T_1375} : _T_337; // @[CSR.scala 277:29:@5726.6]
  assign _T_1376 = _T_336[39:32]; // @[CSR.scala 278:45:@5733.8]
  assign _T_1377 = {_T_1376,wdata}; // @[Cat.scala 30:58:@5734.8]
  assign _GEN_71 = _T_608 ? {{1'd0}, _T_1377} : _GEN_70; // @[CSR.scala 278:29:@5732.6]
  assign _T_1379 = _T_339[31:0]; // @[CSR.scala 277:72:@5739.8]
  assign _T_1380 = {_T_1253,_T_1379}; // @[Cat.scala 30:58:@5740.8]
  assign _GEN_72 = _T_614 ? {{1'd0}, _T_1380} : _T_340; // @[CSR.scala 277:29:@5737.6]
  assign _T_1381 = _T_339[39:32]; // @[CSR.scala 278:45:@5744.8]
  assign _T_1382 = {_T_1381,wdata}; // @[Cat.scala 30:58:@5745.8]
  assign _GEN_73 = _T_612 ? {{1'd0}, _T_1382} : _GEN_72; // @[CSR.scala 278:29:@5743.6]
  assign _T_1384 = _T_342[31:0]; // @[CSR.scala 277:72:@5750.8]
  assign _T_1385 = {_T_1253,_T_1384}; // @[Cat.scala 30:58:@5751.8]
  assign _GEN_74 = _T_618 ? {{1'd0}, _T_1385} : _T_343; // @[CSR.scala 277:29:@5748.6]
  assign _T_1386 = _T_342[39:32]; // @[CSR.scala 278:45:@5755.8]
  assign _T_1387 = {_T_1386,wdata}; // @[Cat.scala 30:58:@5756.8]
  assign _GEN_75 = _T_616 ? {{1'd0}, _T_1387} : _GEN_74; // @[CSR.scala 278:29:@5754.6]
  assign _T_1389 = _T_345[31:0]; // @[CSR.scala 277:72:@5761.8]
  assign _T_1390 = {_T_1253,_T_1389}; // @[Cat.scala 30:58:@5762.8]
  assign _GEN_76 = _T_622 ? {{1'd0}, _T_1390} : _T_346; // @[CSR.scala 277:29:@5759.6]
  assign _T_1391 = _T_345[39:32]; // @[CSR.scala 278:45:@5766.8]
  assign _T_1392 = {_T_1391,wdata}; // @[Cat.scala 30:58:@5767.8]
  assign _GEN_77 = _T_620 ? {{1'd0}, _T_1392} : _GEN_76; // @[CSR.scala 278:29:@5765.6]
  assign _T_1394 = _T_348[31:0]; // @[CSR.scala 277:72:@5772.8]
  assign _T_1395 = {_T_1253,_T_1394}; // @[Cat.scala 30:58:@5773.8]
  assign _GEN_78 = _T_626 ? {{1'd0}, _T_1395} : _T_349; // @[CSR.scala 277:29:@5770.6]
  assign _T_1396 = _T_348[39:32]; // @[CSR.scala 278:45:@5777.8]
  assign _T_1397 = {_T_1396,wdata}; // @[Cat.scala 30:58:@5778.8]
  assign _GEN_79 = _T_624 ? {{1'd0}, _T_1397} : _GEN_78; // @[CSR.scala 278:29:@5776.6]
  assign _T_1399 = _T_351[31:0]; // @[CSR.scala 277:72:@5783.8]
  assign _T_1400 = {_T_1253,_T_1399}; // @[Cat.scala 30:58:@5784.8]
  assign _GEN_80 = _T_630 ? {{1'd0}, _T_1400} : _T_352; // @[CSR.scala 277:29:@5781.6]
  assign _T_1401 = _T_351[39:32]; // @[CSR.scala 278:45:@5788.8]
  assign _T_1402 = {_T_1401,wdata}; // @[Cat.scala 30:58:@5789.8]
  assign _GEN_81 = _T_628 ? {{1'd0}, _T_1402} : _GEN_80; // @[CSR.scala 278:29:@5787.6]
  assign _T_1404 = _T_354[31:0]; // @[CSR.scala 277:72:@5794.8]
  assign _T_1405 = {_T_1253,_T_1404}; // @[Cat.scala 30:58:@5795.8]
  assign _GEN_82 = _T_634 ? {{1'd0}, _T_1405} : _T_355; // @[CSR.scala 277:29:@5792.6]
  assign _T_1406 = _T_354[39:32]; // @[CSR.scala 278:45:@5799.8]
  assign _T_1407 = {_T_1406,wdata}; // @[Cat.scala 30:58:@5800.8]
  assign _GEN_83 = _T_632 ? {{1'd0}, _T_1407} : _GEN_82; // @[CSR.scala 278:29:@5798.6]
  assign _T_1409 = _T_357[31:0]; // @[CSR.scala 277:72:@5805.8]
  assign _T_1410 = {_T_1253,_T_1409}; // @[Cat.scala 30:58:@5806.8]
  assign _GEN_84 = _T_638 ? {{1'd0}, _T_1410} : _T_358; // @[CSR.scala 277:29:@5803.6]
  assign _T_1411 = _T_357[39:32]; // @[CSR.scala 278:45:@5810.8]
  assign _T_1412 = {_T_1411,wdata}; // @[Cat.scala 30:58:@5811.8]
  assign _GEN_85 = _T_636 ? {{1'd0}, _T_1412} : _GEN_84; // @[CSR.scala 278:29:@5809.6]
  assign _T_1414 = _T_249[31:0]; // @[CSR.scala 277:72:@5816.8]
  assign _T_1415 = {wdata,_T_1414}; // @[Cat.scala 30:58:@5817.8]
  assign _T_1416 = _T_1415[63:6]; // @[Util.scala 133:28:@5819.8]
  assign _GEN_86 = _T_640 ? _T_1415 : {{57'd0}, _T_241}; // @[CSR.scala 277:29:@5814.6]
  assign _GEN_87 = _T_640 ? _T_1416 : _GEN_0; // @[CSR.scala 277:29:@5814.6]
  assign _T_1417 = _T_249[63:32]; // @[CSR.scala 278:45:@5823.8]
  assign _T_1418 = {_T_1417,wdata}; // @[Cat.scala 30:58:@5824.8]
  assign _T_1419 = _T_1418[63:6]; // @[Util.scala 133:28:@5826.8]
  assign _GEN_88 = _T_478 ? _T_1418 : _GEN_86; // @[CSR.scala 278:29:@5822.6]
  assign _GEN_89 = _T_478 ? _T_1419 : _GEN_87; // @[CSR.scala 278:29:@5822.6]
  assign _T_1421 = _T_261[31:0]; // @[CSR.scala 277:72:@5831.8]
  assign _T_1422 = {wdata,_T_1421}; // @[Cat.scala 30:58:@5832.8]
  assign _T_1423 = _T_1422[63:6]; // @[Util.scala 133:28:@5834.8]
  assign _GEN_90 = _T_642 ? _T_1422 : {{57'd0}, _T_253}; // @[CSR.scala 277:29:@5829.6]
  assign _GEN_91 = _T_642 ? _T_1423 : _GEN_1; // @[CSR.scala 277:29:@5829.6]
  assign _T_1424 = _T_261[63:32]; // @[CSR.scala 278:45:@5838.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:@5839.8]
  assign _T_1426 = _T_1425[63:6]; // @[Util.scala 133:28:@5841.8]
  assign _GEN_92 = _T_480 ? _T_1425 : _GEN_90; // @[CSR.scala 278:29:@5837.6]
  assign _GEN_93 = _T_480 ? _T_1426 : _GEN_91; // @[CSR.scala 278:29:@5837.6]
  assign _GEN_94 = _T_508 ? wdata : reg_dscratch; // @[CSR.scala 265:40:@5844.6]
  assign _T_1429 = wdata >> 2'h2; // @[CSR.scala 267:78:@5849.8]
  assign _GEN_225 = {{3'd0}, _T_1429}; // @[CSR.scala 267:86:@5850.8]
  assign _T_1431 = _GEN_225 << 2'h2; // @[CSR.scala 267:86:@5850.8]
  assign _GEN_95 = _T_500 ? _T_1431 : {{3'd0}, _GEN_15}; // @[CSR.scala 267:40:@5847.6]
  assign _GEN_96 = _T_498 ? wdata : reg_mscratch; // @[CSR.scala 268:40:@5853.6]
  assign _T_1433 = wdata & 32'h8000001f; // @[CSR.scala 269:62:@5857.8]
  assign _GEN_97 = _T_504 ? _T_1433 : _GEN_14; // @[CSR.scala 269:40:@5856.6]
  assign _GEN_98 = _T_502 ? wdata : _GEN_16; // @[CSR.scala 270:40:@5860.6]
  assign _GEN_99 = _T_510 ? wdata : reg_medeleg; // @[CSR.scala 271:42:@5864.6]
  assign _GEN_100 = wen ? _GEN_17 : _GEN_3; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_101 = wen ? _GEN_18 : _GEN_4; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_102 = wen ? _GEN_19 : reg_mip_msip; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_103 = wen ? _GEN_20 : reg_mie_msip; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_104 = wen ? _GEN_21 : reg_mie_mtip; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_105 = wen ? _GEN_23 : _T_265; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_106 = wen ? _GEN_25 : _T_268; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_107 = wen ? _GEN_27 : _T_271; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_108 = wen ? _GEN_29 : _T_274; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_109 = wen ? _GEN_31 : _T_277; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_110 = wen ? _GEN_33 : _T_280; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_111 = wen ? _GEN_35 : _T_283; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_112 = wen ? _GEN_37 : _T_286; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_113 = wen ? _GEN_39 : _T_289; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_114 = wen ? _GEN_41 : _T_292; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_115 = wen ? _GEN_43 : _T_295; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_116 = wen ? _GEN_45 : _T_298; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_117 = wen ? _GEN_47 : _T_301; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_118 = wen ? _GEN_49 : _T_304; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_119 = wen ? _GEN_51 : _T_307; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_120 = wen ? _GEN_53 : _T_310; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_121 = wen ? _GEN_55 : _T_313; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_122 = wen ? _GEN_57 : _T_316; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_123 = wen ? _GEN_59 : _T_319; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_124 = wen ? _GEN_61 : _T_322; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_125 = wen ? _GEN_63 : _T_325; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_126 = wen ? _GEN_65 : _T_328; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_127 = wen ? _GEN_67 : _T_331; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_128 = wen ? _GEN_69 : _T_334; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_129 = wen ? _GEN_71 : _T_337; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_130 = wen ? _GEN_73 : _T_340; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_131 = wen ? _GEN_75 : _T_343; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_132 = wen ? _GEN_77 : _T_346; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_133 = wen ? _GEN_79 : _T_349; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_134 = wen ? _GEN_81 : _T_352; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_135 = wen ? _GEN_83 : _T_355; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_136 = wen ? _GEN_85 : _T_358; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_137 = wen ? _GEN_88 : {{57'd0}, _T_241}; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_138 = wen ? _GEN_89 : _GEN_0; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_139 = wen ? _GEN_92 : {{57'd0}, _T_253}; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_140 = wen ? _GEN_93 : _GEN_1; // @[CSR.scala 242:14:@5393.4]
  assign _GEN_142 = wen ? _GEN_95 : {{3'd0}, _GEN_15}; // @[CSR.scala 242:14:@5393.4]
  assign io_rw_rdata = _T_1209[31:0]; // @[CSR.scala 240:15:@5392.4]
  assign io_eret = _T_940 | insn_ret; // @[CSR.scala 199:11:@5182.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 197:13:@5179.4]
  assign io_status_unimp5 = 14'h0; // @[CSR.scala 197:13:@5178.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 197:13:@5177.4]
  assign io_status_unimp4 = 2'h0; // @[CSR.scala 197:13:@5176.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 197:13:@5175.4]
  assign io_status_unimp3 = 3'h0; // @[CSR.scala 197:13:@5174.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 197:13:@5173.4]
  assign io_status_unimp2 = 3'h0; // @[CSR.scala 197:13:@5172.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 197:13:@5171.4]
  assign io_status_unimp1 = 3'h0; // @[CSR.scala 197:13:@5170.4]
  assign io_evec = io_xcpt ? 32'h80000004 : _GEN_10; // @[CSR.scala 212:13:@5203.6 CSR.scala 217:13:@5206.6 CSR.scala 224:13:@5213.6 CSR.scala 230:13:@5218.6]
  assign io_time = _T_249[31:0]; // @[CSR.scala 236:11:@5223.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_240 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_244 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_252 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_256 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_264 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_267 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_270 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_273 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_276 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_279 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_282 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_285 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_288 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_291 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_294 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_297 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_300 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_303 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_306 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_309 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_312 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_315 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_318 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_321 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_324 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_327 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_330 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_333 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_336 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_339 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_342 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_345 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_348 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_351 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_354 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_357 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_954) begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mpie <= _T_1222;
        end else begin
          if (_T_954) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mpie <= 1'h1;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mie <= _T_1220;
        end else begin
          if (_T_954) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end
    end
    reg_mepc <= _GEN_142[31:0];
    if (wen) begin
      if (_T_504) begin
        reg_mcause <= _T_1433;
      end else begin
        if (io_xcpt) begin
          reg_mcause <= io_cause;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_959};
            end
          end
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mcause <= io_cause;
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_959};
          end
        end
      end
    end
    if (wen) begin
      if (_T_502) begin
        reg_mtval <= wdata;
      end else begin
        if (io_xcpt) begin
          reg_mtval <= io_tval;
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mtval <= io_tval;
      end
    end
    if (wen) begin
      if (_T_498) begin
        reg_mscratch <= wdata;
      end
    end
    if (wen) begin
      if (_T_510) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (reset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_494) begin
          reg_mip_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_mtip <= _T_1237;
        end
      end
    end
    if (reset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      _T_240 <= 6'h0;
    end else begin
      _T_240 <= _GEN_137[5:0];
    end
    if (reset) begin
      _T_244 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_478) begin
          _T_244 <= _T_1419;
        end else begin
          if (_T_640) begin
            _T_244 <= _T_1416;
          end else begin
            if (_T_245) begin
              _T_244 <= _T_248;
            end
          end
        end
      end else begin
        if (_T_245) begin
          _T_244 <= _T_248;
        end
      end
    end
    if (reset) begin
      _T_252 <= 6'h0;
    end else begin
      _T_252 <= _GEN_139[5:0];
    end
    if (reset) begin
      _T_256 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_480) begin
          _T_256 <= _T_1426;
        end else begin
          if (_T_642) begin
            _T_256 <= _T_1423;
          end else begin
            if (_T_257) begin
              _T_256 <= _T_260;
            end
          end
        end
      end else begin
        if (_T_257) begin
          _T_256 <= _T_260;
        end
      end
    end
    _T_264 <= _GEN_105[39:0];
    _T_267 <= _GEN_106[39:0];
    _T_270 <= _GEN_107[39:0];
    _T_273 <= _GEN_108[39:0];
    _T_276 <= _GEN_109[39:0];
    _T_279 <= _GEN_110[39:0];
    _T_282 <= _GEN_111[39:0];
    _T_285 <= _GEN_112[39:0];
    _T_288 <= _GEN_113[39:0];
    _T_291 <= _GEN_114[39:0];
    _T_294 <= _GEN_115[39:0];
    _T_297 <= _GEN_116[39:0];
    _T_300 <= _GEN_117[39:0];
    _T_303 <= _GEN_118[39:0];
    _T_306 <= _GEN_119[39:0];
    _T_309 <= _GEN_120[39:0];
    _T_312 <= _GEN_121[39:0];
    _T_315 <= _GEN_122[39:0];
    _T_318 <= _GEN_123[39:0];
    _T_321 <= _GEN_124[39:0];
    _T_324 <= _GEN_125[39:0];
    _T_327 <= _GEN_126[39:0];
    _T_330 <= _GEN_127[39:0];
    _T_333 <= _GEN_128[39:0];
    _T_336 <= _GEN_129[39:0];
    _T_339 <= _GEN_130[39:0];
    _T_342 <= _GEN_131[39:0];
    _T_345 <= _GEN_132[39:0];
    _T_348 <= _GEN_133[39:0];
    _T_351 <= _GEN_134[39:0];
    _T_354 <= _GEN_135[39:0];
    _T_357 <= _GEN_136[39:0];
    if (wen) begin
      if (_T_508) begin
        reg_dscratch <= wdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:201 assert(PopCount(insn_ret :: io.illegal :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 201:9:@5189.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[CSR.scala 201:9:@5190.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Regfile( // @[:@5870.2]
  input         clock, // @[:@5871.4]
  input  [4:0]  io_rs1_addr_0, // @[:@5873.4]
  input  [4:0]  io_rs1_addr_1, // @[:@5873.4]
  output [31:0] io_rs1_data_0, // @[:@5873.4]
  output [31:0] io_rs1_data_1, // @[:@5873.4]
  input  [4:0]  io_rs2_addr_0, // @[:@5873.4]
  input  [4:0]  io_rs2_addr_1, // @[:@5873.4]
  output [31:0] io_rs2_data_0, // @[:@5873.4]
  output [31:0] io_rs2_data_1, // @[:@5873.4]
  input  [4:0]  io_waddr_0, // @[:@5873.4]
  input  [4:0]  io_waddr_1, // @[:@5873.4]
  input  [31:0] io_wdata_0, // @[:@5873.4]
  input  [31:0] io_wdata_1, // @[:@5873.4]
  input         io_wen_0, // @[:@5873.4]
  input         io_wen_1 // @[:@5873.4]
);
  reg [31:0] regfile [0:31]; // @[Regfile.scala 23:20:@5875.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_109_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_109_addr; // @[Regfile.scala 23:20:@5875.4]
  wire [31:0] regfile__T_114_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_114_addr; // @[Regfile.scala 23:20:@5875.4]
  wire [31:0] regfile__T_119_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_119_addr; // @[Regfile.scala 23:20:@5875.4]
  wire [31:0] regfile__T_124_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_124_addr; // @[Regfile.scala 23:20:@5875.4]
  wire [31:0] regfile__T_105_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_105_addr; // @[Regfile.scala 23:20:@5875.4]
  wire  regfile__T_105_mask; // @[Regfile.scala 23:20:@5875.4]
  wire  regfile__T_105_en; // @[Regfile.scala 23:20:@5875.4]
  wire [31:0] regfile__T_106_data; // @[Regfile.scala 23:20:@5875.4]
  wire [4:0] regfile__T_106_addr; // @[Regfile.scala 23:20:@5875.4]
  wire  regfile__T_106_mask; // @[Regfile.scala 23:20:@5875.4]
  wire  regfile__T_106_en; // @[Regfile.scala 23:20:@5875.4]
  wire  _T_108; // @[Regfile.scala 28:42:@5884.4]
  wire  _T_113; // @[Regfile.scala 29:42:@5888.4]
  wire  _T_118; // @[Regfile.scala 28:42:@5892.4]
  wire  _T_123; // @[Regfile.scala 29:42:@5896.4]
  assign regfile__T_109_addr = io_rs1_addr_0;
  assign regfile__T_109_data = regfile[regfile__T_109_addr]; // @[Regfile.scala 23:20:@5875.4]
  assign regfile__T_114_addr = io_rs2_addr_0;
  assign regfile__T_114_data = regfile[regfile__T_114_addr]; // @[Regfile.scala 23:20:@5875.4]
  assign regfile__T_119_addr = io_rs1_addr_1;
  assign regfile__T_119_data = regfile[regfile__T_119_addr]; // @[Regfile.scala 23:20:@5875.4]
  assign regfile__T_124_addr = io_rs2_addr_1;
  assign regfile__T_124_data = regfile[regfile__T_124_addr]; // @[Regfile.scala 23:20:@5875.4]
  assign regfile__T_105_data = io_wdata_0;
  assign regfile__T_105_addr = io_waddr_0;
  assign regfile__T_105_mask = 1'h1;
  assign regfile__T_105_en = io_wen_0;
  assign regfile__T_106_data = io_wdata_1;
  assign regfile__T_106_addr = io_waddr_1;
  assign regfile__T_106_mask = 1'h1;
  assign regfile__T_106_en = io_wen_1;
  assign _T_108 = io_rs1_addr_0 != 5'h0; // @[Regfile.scala 28:42:@5884.4]
  assign _T_113 = io_rs2_addr_0 != 5'h0; // @[Regfile.scala 29:42:@5888.4]
  assign _T_118 = io_rs1_addr_1 != 5'h0; // @[Regfile.scala 28:42:@5892.4]
  assign _T_123 = io_rs2_addr_1 != 5'h0; // @[Regfile.scala 29:42:@5896.4]
  assign io_rs1_data_0 = _T_108 ? regfile__T_109_data : 32'h0; // @[Regfile.scala 28:20:@5887.4]
  assign io_rs1_data_1 = _T_118 ? regfile__T_119_data : 32'h0; // @[Regfile.scala 28:20:@5895.4]
  assign io_rs2_data_0 = _T_113 ? regfile__T_114_data : 32'h0; // @[Regfile.scala 29:20:@5891.4]
  assign io_rs2_data_1 = _T_123 ? regfile__T_124_data : 32'h0; // @[Regfile.scala 29:20:@5899.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(regfile__T_105_en & regfile__T_105_mask) begin
      regfile[regfile__T_105_addr] <= regfile__T_105_data; // @[Regfile.scala 23:20:@5875.4]
    end
    if(regfile__T_106_en & regfile__T_106_mask) begin
      regfile[regfile__T_106_addr] <= regfile__T_106_data; // @[Regfile.scala 23:20:@5875.4]
    end
  end
endmodule
module ALU( // @[:@5901.2]
  input  [31:0] io_op1, // @[:@5904.4]
  input  [31:0] io_op2, // @[:@5904.4]
  input  [31:0] io_pc, // @[:@5904.4]
  input  [3:0]  io_ctrl_fun, // @[:@5904.4]
  input  [3:0]  io_ctrl_br_type, // @[:@5904.4]
  input  [1:0]  io_ctrl_wb_sel, // @[:@5904.4]
  output [1:0]  io_ctrl_pc_sel, // @[:@5904.4]
  input  [31:0] io_rs2_data, // @[:@5904.4]
  output [31:0] io_result, // @[:@5904.4]
  output [31:0] io_target_brjmp, // @[:@5904.4]
  output [31:0] io_target_jpreg, // @[:@5904.4]
  output [31:0] io_target_conti // @[:@5904.4]
);
  wire [4:0] alu_shamt; // @[ALU.scala 32:32:@5906.4]
  wire [32:0] _T_25; // @[ALU.scala 33:34:@5907.4]
  wire [31:0] add_result; // @[ALU.scala 33:34:@5908.4]
  wire  _T_29; // @[ALU.scala 38:18:@5911.4]
  wire  _T_30; // @[ALU.scala 39:18:@5912.4]
  wire [32:0] _T_31; // @[ALU.scala 39:44:@5913.4]
  wire [32:0] _T_32; // @[ALU.scala 39:44:@5914.4]
  wire [31:0] _T_33; // @[ALU.scala 39:44:@5915.4]
  wire  _T_34; // @[ALU.scala 40:18:@5916.4]
  wire [31:0] _T_35; // @[ALU.scala 40:44:@5917.4]
  wire  _T_36; // @[ALU.scala 41:18:@5918.4]
  wire [31:0] _T_37; // @[ALU.scala 41:44:@5919.4]
  wire  _T_38; // @[ALU.scala 42:18:@5920.4]
  wire [31:0] _T_39; // @[ALU.scala 42:44:@5921.4]
  wire  _T_40; // @[ALU.scala 43:18:@5922.4]
  wire [31:0] _T_41; // @[ALU.scala 43:44:@5923.4]
  wire [31:0] _T_42; // @[ALU.scala 43:60:@5924.4]
  wire  _T_43; // @[ALU.scala 43:51:@5925.4]
  wire  _T_44; // @[ALU.scala 44:18:@5926.4]
  wire  _T_45; // @[ALU.scala 44:44:@5927.4]
  wire  _T_46; // @[ALU.scala 45:18:@5928.4]
  wire [62:0] _GEN_0; // @[ALU.scala 45:44:@5929.4]
  wire [62:0] _T_47; // @[ALU.scala 45:44:@5929.4]
  wire [31:0] _T_48; // @[ALU.scala 45:57:@5930.4]
  wire  _T_49; // @[ALU.scala 46:18:@5931.4]
  wire [31:0] _T_51; // @[ALU.scala 46:51:@5933.4]
  wire [31:0] _T_52; // @[ALU.scala 46:65:@5934.4]
  wire  _T_53; // @[ALU.scala 47:18:@5935.4]
  wire [31:0] _T_54; // @[ALU.scala 47:44:@5936.4]
  wire  _T_55; // @[ALU.scala 48:18:@5937.4]
  wire  _T_56; // @[ALU.scala 49:18:@5938.4]
  wire [31:0] _T_57; // @[Mux.scala 61:16:@5939.4]
  wire [31:0] _T_58; // @[Mux.scala 61:16:@5940.4]
  wire [31:0] _T_59; // @[Mux.scala 61:16:@5941.4]
  wire [31:0] _T_60; // @[Mux.scala 61:16:@5942.4]
  wire [31:0] _T_61; // @[Mux.scala 61:16:@5943.4]
  wire [31:0] _T_62; // @[Mux.scala 61:16:@5944.4]
  wire [31:0] _T_63; // @[Mux.scala 61:16:@5945.4]
  wire [31:0] _T_64; // @[Mux.scala 61:16:@5946.4]
  wire [31:0] _T_65; // @[Mux.scala 61:16:@5947.4]
  wire [31:0] _T_66; // @[Mux.scala 61:16:@5948.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@5949.4]
  wire [31:0] result; // @[Mux.scala 61:16:@5950.4]
  wire [32:0] _T_69; // @[ALU.scala 52:31:@5952.4]
  wire [30:0] _T_71; // @[ALU.scala 53:39:@5955.4]
  wire [32:0] _T_75; // @[ALU.scala 54:31:@5958.4]
  wire  _T_77; // @[ALU.scala 55:35:@5961.4]
  wire  br_eq; // @[ALU.scala 57:29:@5964.4]
  wire [31:0] _T_80; // @[ALU.scala 58:50:@5966.4]
  wire  br_lt; // @[ALU.scala 58:36:@5967.4]
  wire  br_ltu; // @[ALU.scala 59:36:@5968.4]
  wire  _T_81; // @[ALU.scala 63:25:@5969.4]
  wire  _T_82; // @[ALU.scala 64:25:@5970.4]
  wire  _T_84; // @[ALU.scala 64:41:@5971.4]
  wire [1:0] _T_85; // @[ALU.scala 64:40:@5972.4]
  wire  _T_86; // @[ALU.scala 65:25:@5973.4]
  wire [1:0] _T_87; // @[ALU.scala 65:40:@5974.4]
  wire  _T_88; // @[ALU.scala 66:25:@5975.4]
  wire  _T_90; // @[ALU.scala 66:41:@5976.4]
  wire [1:0] _T_91; // @[ALU.scala 66:40:@5977.4]
  wire  _T_92; // @[ALU.scala 67:25:@5978.4]
  wire  _T_94; // @[ALU.scala 67:41:@5979.4]
  wire [1:0] _T_95; // @[ALU.scala 67:40:@5980.4]
  wire  _T_96; // @[ALU.scala 68:25:@5981.4]
  wire [1:0] _T_97; // @[ALU.scala 68:40:@5982.4]
  wire  _T_98; // @[ALU.scala 69:25:@5983.4]
  wire [1:0] _T_99; // @[ALU.scala 69:40:@5984.4]
  wire  _T_100; // @[ALU.scala 70:25:@5985.4]
  wire  _T_101; // @[ALU.scala 71:25:@5986.4]
  wire [1:0] _T_102; // @[ALU.scala 71:8:@5987.4]
  wire [1:0] _T_103; // @[ALU.scala 70:8:@5988.4]
  wire [1:0] _T_104; // @[ALU.scala 69:8:@5989.4]
  wire [1:0] _T_105; // @[ALU.scala 68:8:@5990.4]
  wire [1:0] _T_106; // @[ALU.scala 67:8:@5991.4]
  wire [1:0] _T_107; // @[ALU.scala 66:8:@5992.4]
  wire [1:0] _T_108; // @[ALU.scala 65:8:@5993.4]
  wire [1:0] _T_109; // @[ALU.scala 64:8:@5994.4]
  assign alu_shamt = io_op2[4:0]; // @[ALU.scala 32:32:@5906.4]
  assign _T_25 = io_op1 + io_op2; // @[ALU.scala 33:34:@5907.4]
  assign add_result = io_op1 + io_op2; // @[ALU.scala 33:34:@5908.4]
  assign _T_29 = io_ctrl_fun == 4'h0; // @[ALU.scala 38:18:@5911.4]
  assign _T_30 = io_ctrl_fun == 4'h1; // @[ALU.scala 39:18:@5912.4]
  assign _T_31 = io_op1 - io_op2; // @[ALU.scala 39:44:@5913.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 39:44:@5914.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 39:44:@5915.4]
  assign _T_34 = io_ctrl_fun == 4'h5; // @[ALU.scala 40:18:@5916.4]
  assign _T_35 = io_op1 & io_op2; // @[ALU.scala 40:44:@5917.4]
  assign _T_36 = io_ctrl_fun == 4'h6; // @[ALU.scala 41:18:@5918.4]
  assign _T_37 = io_op1 | io_op2; // @[ALU.scala 41:44:@5919.4]
  assign _T_38 = io_ctrl_fun == 4'h7; // @[ALU.scala 42:18:@5920.4]
  assign _T_39 = io_op1 ^ io_op2; // @[ALU.scala 42:44:@5921.4]
  assign _T_40 = io_ctrl_fun == 4'h8; // @[ALU.scala 43:18:@5922.4]
  assign _T_41 = $signed(io_op1); // @[ALU.scala 43:44:@5923.4]
  assign _T_42 = $signed(io_op2); // @[ALU.scala 43:60:@5924.4]
  assign _T_43 = $signed(_T_41) < $signed(_T_42); // @[ALU.scala 43:51:@5925.4]
  assign _T_44 = io_ctrl_fun == 4'h9; // @[ALU.scala 44:18:@5926.4]
  assign _T_45 = io_op1 < io_op2; // @[ALU.scala 44:44:@5927.4]
  assign _T_46 = io_ctrl_fun == 4'h2; // @[ALU.scala 45:18:@5928.4]
  assign _GEN_0 = {{31'd0}, io_op1}; // @[ALU.scala 45:44:@5929.4]
  assign _T_47 = _GEN_0 << alu_shamt; // @[ALU.scala 45:44:@5929.4]
  assign _T_48 = _T_47[31:0]; // @[ALU.scala 45:57:@5930.4]
  assign _T_49 = io_ctrl_fun == 4'h4; // @[ALU.scala 46:18:@5931.4]
  assign _T_51 = $signed(_T_41) >>> alu_shamt; // @[ALU.scala 46:51:@5933.4]
  assign _T_52 = $unsigned(_T_51); // @[ALU.scala 46:65:@5934.4]
  assign _T_53 = io_ctrl_fun == 4'h3; // @[ALU.scala 47:18:@5935.4]
  assign _T_54 = io_op1 >> alu_shamt; // @[ALU.scala 47:44:@5936.4]
  assign _T_55 = io_ctrl_fun == 4'ha; // @[ALU.scala 48:18:@5937.4]
  assign _T_56 = io_ctrl_fun == 4'hb; // @[ALU.scala 49:18:@5938.4]
  assign _T_57 = _T_56 ? io_op2 : 32'h0; // @[Mux.scala 61:16:@5939.4]
  assign _T_58 = _T_55 ? io_op1 : _T_57; // @[Mux.scala 61:16:@5940.4]
  assign _T_59 = _T_53 ? _T_54 : _T_58; // @[Mux.scala 61:16:@5941.4]
  assign _T_60 = _T_49 ? _T_52 : _T_59; // @[Mux.scala 61:16:@5942.4]
  assign _T_61 = _T_46 ? _T_48 : _T_60; // @[Mux.scala 61:16:@5943.4]
  assign _T_62 = _T_44 ? {{31'd0}, _T_45} : _T_61; // @[Mux.scala 61:16:@5944.4]
  assign _T_63 = _T_40 ? {{31'd0}, _T_43} : _T_62; // @[Mux.scala 61:16:@5945.4]
  assign _T_64 = _T_38 ? _T_39 : _T_63; // @[Mux.scala 61:16:@5946.4]
  assign _T_65 = _T_36 ? _T_37 : _T_64; // @[Mux.scala 61:16:@5947.4]
  assign _T_66 = _T_34 ? _T_35 : _T_65; // @[Mux.scala 61:16:@5948.4]
  assign _T_67 = _T_30 ? _T_33 : _T_66; // @[Mux.scala 61:16:@5949.4]
  assign result = _T_29 ? add_result : _T_67; // @[Mux.scala 61:16:@5950.4]
  assign _T_69 = io_pc + io_op2; // @[ALU.scala 52:31:@5952.4]
  assign _T_71 = add_result[31:1]; // @[ALU.scala 53:39:@5955.4]
  assign _T_75 = io_pc + 32'h4; // @[ALU.scala 54:31:@5958.4]
  assign _T_77 = io_ctrl_wb_sel == 2'h2; // @[ALU.scala 55:35:@5961.4]
  assign br_eq = io_op1 == io_rs2_data; // @[ALU.scala 57:29:@5964.4]
  assign _T_80 = $signed(io_rs2_data); // @[ALU.scala 58:50:@5966.4]
  assign br_lt = $signed(_T_41) < $signed(_T_80); // @[ALU.scala 58:36:@5967.4]
  assign br_ltu = io_op1 < io_rs2_data; // @[ALU.scala 59:36:@5968.4]
  assign _T_81 = io_ctrl_br_type == 4'h0; // @[ALU.scala 63:25:@5969.4]
  assign _T_82 = io_ctrl_br_type == 4'h1; // @[ALU.scala 64:25:@5970.4]
  assign _T_84 = br_eq == 1'h0; // @[ALU.scala 64:41:@5971.4]
  assign _T_85 = _T_84 ? 2'h1 : 2'h0; // @[ALU.scala 64:40:@5972.4]
  assign _T_86 = io_ctrl_br_type == 4'h2; // @[ALU.scala 65:25:@5973.4]
  assign _T_87 = br_eq ? 2'h1 : 2'h0; // @[ALU.scala 65:40:@5974.4]
  assign _T_88 = io_ctrl_br_type == 4'h3; // @[ALU.scala 66:25:@5975.4]
  assign _T_90 = br_lt == 1'h0; // @[ALU.scala 66:41:@5976.4]
  assign _T_91 = _T_90 ? 2'h1 : 2'h0; // @[ALU.scala 66:40:@5977.4]
  assign _T_92 = io_ctrl_br_type == 4'h4; // @[ALU.scala 67:25:@5978.4]
  assign _T_94 = br_ltu == 1'h0; // @[ALU.scala 67:41:@5979.4]
  assign _T_95 = _T_94 ? 2'h1 : 2'h0; // @[ALU.scala 67:40:@5980.4]
  assign _T_96 = io_ctrl_br_type == 4'h5; // @[ALU.scala 68:25:@5981.4]
  assign _T_97 = br_lt ? 2'h1 : 2'h0; // @[ALU.scala 68:40:@5982.4]
  assign _T_98 = io_ctrl_br_type == 4'h6; // @[ALU.scala 69:25:@5983.4]
  assign _T_99 = br_ltu ? 2'h1 : 2'h0; // @[ALU.scala 69:40:@5984.4]
  assign _T_100 = io_ctrl_br_type == 4'h7; // @[ALU.scala 70:25:@5985.4]
  assign _T_101 = io_ctrl_br_type == 4'h8; // @[ALU.scala 71:25:@5986.4]
  assign _T_102 = _T_101 ? 2'h2 : 2'h0; // @[ALU.scala 71:8:@5987.4]
  assign _T_103 = _T_100 ? 2'h1 : _T_102; // @[ALU.scala 70:8:@5988.4]
  assign _T_104 = _T_98 ? _T_99 : _T_103; // @[ALU.scala 69:8:@5989.4]
  assign _T_105 = _T_96 ? _T_97 : _T_104; // @[ALU.scala 68:8:@5990.4]
  assign _T_106 = _T_92 ? _T_95 : _T_105; // @[ALU.scala 67:8:@5991.4]
  assign _T_107 = _T_88 ? _T_91 : _T_106; // @[ALU.scala 66:8:@5992.4]
  assign _T_108 = _T_86 ? _T_87 : _T_107; // @[ALU.scala 65:8:@5993.4]
  assign _T_109 = _T_82 ? _T_85 : _T_108; // @[ALU.scala 64:8:@5994.4]
  assign io_ctrl_pc_sel = _T_81 ? 2'h0 : _T_109; // @[ALU.scala 62:18:@5996.4]
  assign io_result = _T_77 ? io_target_conti : result; // @[ALU.scala 55:13:@5963.4]
  assign io_target_brjmp = io_pc + io_op2; // @[ALU.scala 52:22:@5954.4]
  assign io_target_jpreg = {_T_71,1'h0}; // @[ALU.scala 53:22:@5957.4]
  assign io_target_conti = io_pc + 32'h4; // @[ALU.scala 54:22:@5960.4]
endmodule
module InstDecoder( // @[:@6095.2]
  input  [31:0] io_inst, // @[:@6098.4]
  output [3:0]  io_cinfo_br_type, // @[:@6098.4]
  output [1:0]  io_cinfo_op1_sel, // @[:@6098.4]
  output [2:0]  io_cinfo_op2_sel, // @[:@6098.4]
  output        io_cinfo_rs1_oen, // @[:@6098.4]
  output        io_cinfo_rs2_oen, // @[:@6098.4]
  output [3:0]  io_cinfo_alu_fun, // @[:@6098.4]
  output [1:0]  io_cinfo_wb_sel, // @[:@6098.4]
  output        io_cinfo_rf_wen, // @[:@6098.4]
  output        io_cinfo_mem_en, // @[:@6098.4]
  output        io_cinfo_mem_fcn, // @[:@6098.4]
  output [2:0]  io_cinfo_mem_typ, // @[:@6098.4]
  output [2:0]  io_cinfo_csr_cmd, // @[:@6098.4]
  output        io_cinfo_illegal, // @[:@6098.4]
  output [31:0] io_dinfo_imm_i, // @[:@6098.4]
  output [31:0] io_dinfo_imm_s, // @[:@6098.4]
  output [31:0] io_dinfo_imm_sb, // @[:@6098.4]
  output [31:0] io_dinfo_imm_u, // @[:@6098.4]
  output [31:0] io_dinfo_imm_uj, // @[:@6098.4]
  output [31:0] io_dinfo_imm_z, // @[:@6098.4]
  output [4:0]  io_rs1_addr, // @[:@6098.4]
  output [4:0]  io_rs2_addr, // @[:@6098.4]
  output [4:0]  io_wbaddr // @[:@6098.4]
);
  wire [31:0] _T_19; // @[Lookup.scala 9:38:@6100.4]
  wire  _T_20; // @[Lookup.scala 9:38:@6101.4]
  wire  _T_24; // @[Lookup.scala 9:38:@6103.4]
  wire  _T_28; // @[Lookup.scala 9:38:@6105.4]
  wire  _T_32; // @[Lookup.scala 9:38:@6107.4]
  wire  _T_36; // @[Lookup.scala 9:38:@6109.4]
  wire  _T_40; // @[Lookup.scala 9:38:@6111.4]
  wire  _T_44; // @[Lookup.scala 9:38:@6113.4]
  wire  _T_48; // @[Lookup.scala 9:38:@6115.4]
  wire [31:0] _T_51; // @[Lookup.scala 9:38:@6116.4]
  wire  _T_52; // @[Lookup.scala 9:38:@6117.4]
  wire  _T_56; // @[Lookup.scala 9:38:@6119.4]
  wire  _T_60; // @[Lookup.scala 9:38:@6121.4]
  wire  _T_64; // @[Lookup.scala 9:38:@6123.4]
  wire  _T_68; // @[Lookup.scala 9:38:@6125.4]
  wire  _T_72; // @[Lookup.scala 9:38:@6127.4]
  wire  _T_76; // @[Lookup.scala 9:38:@6129.4]
  wire  _T_80; // @[Lookup.scala 9:38:@6131.4]
  wire [31:0] _T_83; // @[Lookup.scala 9:38:@6132.4]
  wire  _T_84; // @[Lookup.scala 9:38:@6133.4]
  wire  _T_88; // @[Lookup.scala 9:38:@6135.4]
  wire  _T_92; // @[Lookup.scala 9:38:@6137.4]
  wire [31:0] _T_95; // @[Lookup.scala 9:38:@6138.4]
  wire  _T_96; // @[Lookup.scala 9:38:@6139.4]
  wire  _T_100; // @[Lookup.scala 9:38:@6141.4]
  wire  _T_104; // @[Lookup.scala 9:38:@6143.4]
  wire  _T_108; // @[Lookup.scala 9:38:@6145.4]
  wire  _T_112; // @[Lookup.scala 9:38:@6147.4]
  wire  _T_116; // @[Lookup.scala 9:38:@6149.4]
  wire  _T_120; // @[Lookup.scala 9:38:@6151.4]
  wire  _T_124; // @[Lookup.scala 9:38:@6153.4]
  wire  _T_128; // @[Lookup.scala 9:38:@6155.4]
  wire  _T_132; // @[Lookup.scala 9:38:@6157.4]
  wire  _T_136; // @[Lookup.scala 9:38:@6159.4]
  wire  _T_140; // @[Lookup.scala 9:38:@6161.4]
  wire  _T_144; // @[Lookup.scala 9:38:@6163.4]
  wire  _T_148; // @[Lookup.scala 9:38:@6165.4]
  wire  _T_152; // @[Lookup.scala 9:38:@6167.4]
  wire  _T_156; // @[Lookup.scala 9:38:@6169.4]
  wire  _T_160; // @[Lookup.scala 9:38:@6171.4]
  wire  _T_164; // @[Lookup.scala 9:38:@6173.4]
  wire  _T_168; // @[Lookup.scala 9:38:@6175.4]
  wire  _T_172; // @[Lookup.scala 9:38:@6177.4]
  wire  _T_176; // @[Lookup.scala 9:38:@6179.4]
  wire  _T_180; // @[Lookup.scala 9:38:@6181.4]
  wire  _T_184; // @[Lookup.scala 9:38:@6183.4]
  wire  _T_188; // @[Lookup.scala 9:38:@6185.4]
  wire  _T_192; // @[Lookup.scala 9:38:@6187.4]
  wire  _T_196; // @[Lookup.scala 9:38:@6189.4]
  wire  _T_200; // @[Lookup.scala 9:38:@6191.4]
  wire  _T_204; // @[Lookup.scala 9:38:@6193.4]
  wire  _T_208; // @[Lookup.scala 9:38:@6195.4]
  wire  _T_212; // @[Lookup.scala 9:38:@6197.4]
  wire  _T_216; // @[Lookup.scala 9:38:@6199.4]
  wire  _T_218; // @[Lookup.scala 11:37:@6201.4]
  wire  _T_219; // @[Lookup.scala 11:37:@6202.4]
  wire  _T_220; // @[Lookup.scala 11:37:@6203.4]
  wire  _T_221; // @[Lookup.scala 11:37:@6204.4]
  wire  _T_222; // @[Lookup.scala 11:37:@6205.4]
  wire  _T_223; // @[Lookup.scala 11:37:@6206.4]
  wire  _T_224; // @[Lookup.scala 11:37:@6207.4]
  wire  _T_225; // @[Lookup.scala 11:37:@6208.4]
  wire  _T_226; // @[Lookup.scala 11:37:@6209.4]
  wire  _T_227; // @[Lookup.scala 11:37:@6210.4]
  wire  _T_228; // @[Lookup.scala 11:37:@6211.4]
  wire  _T_229; // @[Lookup.scala 11:37:@6212.4]
  wire  _T_230; // @[Lookup.scala 11:37:@6213.4]
  wire  _T_231; // @[Lookup.scala 11:37:@6214.4]
  wire  _T_232; // @[Lookup.scala 11:37:@6215.4]
  wire  _T_233; // @[Lookup.scala 11:37:@6216.4]
  wire  _T_234; // @[Lookup.scala 11:37:@6217.4]
  wire  _T_235; // @[Lookup.scala 11:37:@6218.4]
  wire  _T_236; // @[Lookup.scala 11:37:@6219.4]
  wire  _T_237; // @[Lookup.scala 11:37:@6220.4]
  wire  _T_238; // @[Lookup.scala 11:37:@6221.4]
  wire  _T_239; // @[Lookup.scala 11:37:@6222.4]
  wire  _T_240; // @[Lookup.scala 11:37:@6223.4]
  wire  _T_241; // @[Lookup.scala 11:37:@6224.4]
  wire  _T_242; // @[Lookup.scala 11:37:@6225.4]
  wire  _T_243; // @[Lookup.scala 11:37:@6226.4]
  wire  _T_244; // @[Lookup.scala 11:37:@6227.4]
  wire  _T_245; // @[Lookup.scala 11:37:@6228.4]
  wire  _T_246; // @[Lookup.scala 11:37:@6229.4]
  wire  _T_247; // @[Lookup.scala 11:37:@6230.4]
  wire  _T_248; // @[Lookup.scala 11:37:@6231.4]
  wire  _T_249; // @[Lookup.scala 11:37:@6232.4]
  wire  _T_250; // @[Lookup.scala 11:37:@6233.4]
  wire  _T_251; // @[Lookup.scala 11:37:@6234.4]
  wire  _T_252; // @[Lookup.scala 11:37:@6235.4]
  wire  _T_253; // @[Lookup.scala 11:37:@6236.4]
  wire  _T_254; // @[Lookup.scala 11:37:@6237.4]
  wire  _T_255; // @[Lookup.scala 11:37:@6238.4]
  wire  _T_256; // @[Lookup.scala 11:37:@6239.4]
  wire  _T_257; // @[Lookup.scala 11:37:@6240.4]
  wire  _T_258; // @[Lookup.scala 11:37:@6241.4]
  wire  _T_259; // @[Lookup.scala 11:37:@6242.4]
  wire  _T_260; // @[Lookup.scala 11:37:@6243.4]
  wire  _T_261; // @[Lookup.scala 11:37:@6244.4]
  wire  _T_262; // @[Lookup.scala 11:37:@6245.4]
  wire  _T_263; // @[Lookup.scala 11:37:@6246.4]
  wire  _T_264; // @[Lookup.scala 11:37:@6247.4]
  wire  _T_265; // @[Lookup.scala 11:37:@6248.4]
  wire  signals_0; // @[Lookup.scala 11:37:@6249.4]
  wire [3:0] _T_279; // @[Lookup.scala 11:37:@6263.4]
  wire [3:0] _T_280; // @[Lookup.scala 11:37:@6264.4]
  wire [3:0] _T_281; // @[Lookup.scala 11:37:@6265.4]
  wire [3:0] _T_282; // @[Lookup.scala 11:37:@6266.4]
  wire [3:0] _T_283; // @[Lookup.scala 11:37:@6267.4]
  wire [3:0] _T_284; // @[Lookup.scala 11:37:@6268.4]
  wire [3:0] _T_285; // @[Lookup.scala 11:37:@6269.4]
  wire [3:0] _T_286; // @[Lookup.scala 11:37:@6270.4]
  wire [3:0] _T_287; // @[Lookup.scala 11:37:@6271.4]
  wire [3:0] _T_288; // @[Lookup.scala 11:37:@6272.4]
  wire [3:0] _T_289; // @[Lookup.scala 11:37:@6273.4]
  wire [3:0] _T_290; // @[Lookup.scala 11:37:@6274.4]
  wire [3:0] _T_291; // @[Lookup.scala 11:37:@6275.4]
  wire [3:0] _T_292; // @[Lookup.scala 11:37:@6276.4]
  wire [3:0] _T_293; // @[Lookup.scala 11:37:@6277.4]
  wire [3:0] _T_294; // @[Lookup.scala 11:37:@6278.4]
  wire [3:0] _T_295; // @[Lookup.scala 11:37:@6279.4]
  wire [3:0] _T_296; // @[Lookup.scala 11:37:@6280.4]
  wire [3:0] _T_297; // @[Lookup.scala 11:37:@6281.4]
  wire [3:0] _T_298; // @[Lookup.scala 11:37:@6282.4]
  wire [3:0] _T_299; // @[Lookup.scala 11:37:@6283.4]
  wire [3:0] _T_300; // @[Lookup.scala 11:37:@6284.4]
  wire [3:0] _T_301; // @[Lookup.scala 11:37:@6285.4]
  wire [3:0] _T_302; // @[Lookup.scala 11:37:@6286.4]
  wire [3:0] _T_303; // @[Lookup.scala 11:37:@6287.4]
  wire [3:0] _T_304; // @[Lookup.scala 11:37:@6288.4]
  wire [3:0] _T_305; // @[Lookup.scala 11:37:@6289.4]
  wire [3:0] _T_306; // @[Lookup.scala 11:37:@6290.4]
  wire [3:0] _T_307; // @[Lookup.scala 11:37:@6291.4]
  wire [3:0] _T_308; // @[Lookup.scala 11:37:@6292.4]
  wire [3:0] _T_309; // @[Lookup.scala 11:37:@6293.4]
  wire [3:0] _T_310; // @[Lookup.scala 11:37:@6294.4]
  wire [3:0] _T_311; // @[Lookup.scala 11:37:@6295.4]
  wire [3:0] _T_312; // @[Lookup.scala 11:37:@6296.4]
  wire [3:0] _T_313; // @[Lookup.scala 11:37:@6297.4]
  wire [3:0] _T_314; // @[Lookup.scala 11:37:@6298.4]
  wire [1:0] _T_322; // @[Lookup.scala 11:37:@6307.4]
  wire [1:0] _T_323; // @[Lookup.scala 11:37:@6308.4]
  wire [1:0] _T_324; // @[Lookup.scala 11:37:@6309.4]
  wire [1:0] _T_325; // @[Lookup.scala 11:37:@6310.4]
  wire [1:0] _T_326; // @[Lookup.scala 11:37:@6311.4]
  wire [1:0] _T_327; // @[Lookup.scala 11:37:@6312.4]
  wire [1:0] _T_328; // @[Lookup.scala 11:37:@6313.4]
  wire [1:0] _T_329; // @[Lookup.scala 11:37:@6314.4]
  wire [1:0] _T_330; // @[Lookup.scala 11:37:@6315.4]
  wire [1:0] _T_331; // @[Lookup.scala 11:37:@6316.4]
  wire [1:0] _T_332; // @[Lookup.scala 11:37:@6317.4]
  wire [1:0] _T_333; // @[Lookup.scala 11:37:@6318.4]
  wire [1:0] _T_334; // @[Lookup.scala 11:37:@6319.4]
  wire [1:0] _T_335; // @[Lookup.scala 11:37:@6320.4]
  wire [1:0] _T_336; // @[Lookup.scala 11:37:@6321.4]
  wire [1:0] _T_337; // @[Lookup.scala 11:37:@6322.4]
  wire [1:0] _T_338; // @[Lookup.scala 11:37:@6323.4]
  wire [1:0] _T_339; // @[Lookup.scala 11:37:@6324.4]
  wire [1:0] _T_340; // @[Lookup.scala 11:37:@6325.4]
  wire [1:0] _T_341; // @[Lookup.scala 11:37:@6326.4]
  wire [1:0] _T_342; // @[Lookup.scala 11:37:@6327.4]
  wire [1:0] _T_343; // @[Lookup.scala 11:37:@6328.4]
  wire [1:0] _T_344; // @[Lookup.scala 11:37:@6329.4]
  wire [1:0] _T_345; // @[Lookup.scala 11:37:@6330.4]
  wire [1:0] _T_346; // @[Lookup.scala 11:37:@6331.4]
  wire [1:0] _T_347; // @[Lookup.scala 11:37:@6332.4]
  wire [1:0] _T_348; // @[Lookup.scala 11:37:@6333.4]
  wire [1:0] _T_349; // @[Lookup.scala 11:37:@6334.4]
  wire [1:0] _T_350; // @[Lookup.scala 11:37:@6335.4]
  wire [1:0] _T_351; // @[Lookup.scala 11:37:@6336.4]
  wire [1:0] _T_352; // @[Lookup.scala 11:37:@6337.4]
  wire [1:0] _T_353; // @[Lookup.scala 11:37:@6338.4]
  wire [1:0] _T_354; // @[Lookup.scala 11:37:@6339.4]
  wire [1:0] _T_355; // @[Lookup.scala 11:37:@6340.4]
  wire [1:0] _T_356; // @[Lookup.scala 11:37:@6341.4]
  wire [1:0] _T_357; // @[Lookup.scala 11:37:@6342.4]
  wire [1:0] _T_358; // @[Lookup.scala 11:37:@6343.4]
  wire [1:0] _T_359; // @[Lookup.scala 11:37:@6344.4]
  wire [1:0] _T_360; // @[Lookup.scala 11:37:@6345.4]
  wire [1:0] _T_361; // @[Lookup.scala 11:37:@6346.4]
  wire [1:0] _T_362; // @[Lookup.scala 11:37:@6347.4]
  wire [1:0] _T_363; // @[Lookup.scala 11:37:@6348.4]
  wire [2:0] _T_377; // @[Lookup.scala 11:37:@6363.4]
  wire [2:0] _T_378; // @[Lookup.scala 11:37:@6364.4]
  wire [2:0] _T_379; // @[Lookup.scala 11:37:@6365.4]
  wire [2:0] _T_380; // @[Lookup.scala 11:37:@6366.4]
  wire [2:0] _T_381; // @[Lookup.scala 11:37:@6367.4]
  wire [2:0] _T_382; // @[Lookup.scala 11:37:@6368.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@6369.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@6370.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@6371.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@6372.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@6373.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@6374.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@6375.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@6376.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@6377.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@6378.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@6379.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@6380.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@6381.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@6382.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@6383.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@6384.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@6385.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@6386.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@6387.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@6388.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@6389.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@6390.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@6391.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@6392.4]
  wire [2:0] _T_407; // @[Lookup.scala 11:37:@6393.4]
  wire [2:0] _T_408; // @[Lookup.scala 11:37:@6394.4]
  wire [2:0] _T_409; // @[Lookup.scala 11:37:@6395.4]
  wire [2:0] _T_410; // @[Lookup.scala 11:37:@6396.4]
  wire [2:0] _T_411; // @[Lookup.scala 11:37:@6397.4]
  wire [2:0] _T_412; // @[Lookup.scala 11:37:@6398.4]
  wire  _T_421; // @[Lookup.scala 11:37:@6408.4]
  wire  _T_422; // @[Lookup.scala 11:37:@6409.4]
  wire  _T_423; // @[Lookup.scala 11:37:@6410.4]
  wire  _T_424; // @[Lookup.scala 11:37:@6411.4]
  wire  _T_425; // @[Lookup.scala 11:37:@6412.4]
  wire  _T_426; // @[Lookup.scala 11:37:@6413.4]
  wire  _T_427; // @[Lookup.scala 11:37:@6414.4]
  wire  _T_428; // @[Lookup.scala 11:37:@6415.4]
  wire  _T_429; // @[Lookup.scala 11:37:@6416.4]
  wire  _T_430; // @[Lookup.scala 11:37:@6417.4]
  wire  _T_431; // @[Lookup.scala 11:37:@6418.4]
  wire  _T_432; // @[Lookup.scala 11:37:@6419.4]
  wire  _T_433; // @[Lookup.scala 11:37:@6420.4]
  wire  _T_434; // @[Lookup.scala 11:37:@6421.4]
  wire  _T_435; // @[Lookup.scala 11:37:@6422.4]
  wire  _T_436; // @[Lookup.scala 11:37:@6423.4]
  wire  _T_437; // @[Lookup.scala 11:37:@6424.4]
  wire  _T_438; // @[Lookup.scala 11:37:@6425.4]
  wire  _T_439; // @[Lookup.scala 11:37:@6426.4]
  wire  _T_440; // @[Lookup.scala 11:37:@6427.4]
  wire  _T_441; // @[Lookup.scala 11:37:@6428.4]
  wire  _T_442; // @[Lookup.scala 11:37:@6429.4]
  wire  _T_443; // @[Lookup.scala 11:37:@6430.4]
  wire  _T_444; // @[Lookup.scala 11:37:@6431.4]
  wire  _T_445; // @[Lookup.scala 11:37:@6432.4]
  wire  _T_446; // @[Lookup.scala 11:37:@6433.4]
  wire  _T_447; // @[Lookup.scala 11:37:@6434.4]
  wire  _T_448; // @[Lookup.scala 11:37:@6435.4]
  wire  _T_449; // @[Lookup.scala 11:37:@6436.4]
  wire  _T_450; // @[Lookup.scala 11:37:@6437.4]
  wire  _T_451; // @[Lookup.scala 11:37:@6438.4]
  wire  _T_452; // @[Lookup.scala 11:37:@6439.4]
  wire  _T_453; // @[Lookup.scala 11:37:@6440.4]
  wire  _T_454; // @[Lookup.scala 11:37:@6441.4]
  wire  _T_455; // @[Lookup.scala 11:37:@6442.4]
  wire  _T_456; // @[Lookup.scala 11:37:@6443.4]
  wire  _T_457; // @[Lookup.scala 11:37:@6444.4]
  wire  _T_458; // @[Lookup.scala 11:37:@6445.4]
  wire  _T_459; // @[Lookup.scala 11:37:@6446.4]
  wire  _T_460; // @[Lookup.scala 11:37:@6447.4]
  wire  _T_461; // @[Lookup.scala 11:37:@6448.4]
  wire  _T_481; // @[Lookup.scala 11:37:@6469.4]
  wire  _T_482; // @[Lookup.scala 11:37:@6470.4]
  wire  _T_483; // @[Lookup.scala 11:37:@6471.4]
  wire  _T_484; // @[Lookup.scala 11:37:@6472.4]
  wire  _T_485; // @[Lookup.scala 11:37:@6473.4]
  wire  _T_486; // @[Lookup.scala 11:37:@6474.4]
  wire  _T_487; // @[Lookup.scala 11:37:@6475.4]
  wire  _T_488; // @[Lookup.scala 11:37:@6476.4]
  wire  _T_489; // @[Lookup.scala 11:37:@6477.4]
  wire  _T_490; // @[Lookup.scala 11:37:@6478.4]
  wire  _T_491; // @[Lookup.scala 11:37:@6479.4]
  wire  _T_492; // @[Lookup.scala 11:37:@6480.4]
  wire  _T_493; // @[Lookup.scala 11:37:@6481.4]
  wire  _T_494; // @[Lookup.scala 11:37:@6482.4]
  wire  _T_495; // @[Lookup.scala 11:37:@6483.4]
  wire  _T_496; // @[Lookup.scala 11:37:@6484.4]
  wire  _T_497; // @[Lookup.scala 11:37:@6485.4]
  wire  _T_498; // @[Lookup.scala 11:37:@6486.4]
  wire  _T_499; // @[Lookup.scala 11:37:@6487.4]
  wire  _T_500; // @[Lookup.scala 11:37:@6488.4]
  wire  _T_501; // @[Lookup.scala 11:37:@6489.4]
  wire  _T_502; // @[Lookup.scala 11:37:@6490.4]
  wire  _T_503; // @[Lookup.scala 11:37:@6491.4]
  wire  _T_504; // @[Lookup.scala 11:37:@6492.4]
  wire  _T_505; // @[Lookup.scala 11:37:@6493.4]
  wire  _T_506; // @[Lookup.scala 11:37:@6494.4]
  wire  _T_507; // @[Lookup.scala 11:37:@6495.4]
  wire  _T_508; // @[Lookup.scala 11:37:@6496.4]
  wire  _T_509; // @[Lookup.scala 11:37:@6497.4]
  wire  _T_510; // @[Lookup.scala 11:37:@6498.4]
  wire [3:0] _T_518; // @[Lookup.scala 11:37:@6507.4]
  wire [3:0] _T_519; // @[Lookup.scala 11:37:@6508.4]
  wire [3:0] _T_520; // @[Lookup.scala 11:37:@6509.4]
  wire [3:0] _T_521; // @[Lookup.scala 11:37:@6510.4]
  wire [3:0] _T_522; // @[Lookup.scala 11:37:@6511.4]
  wire [3:0] _T_523; // @[Lookup.scala 11:37:@6512.4]
  wire [3:0] _T_524; // @[Lookup.scala 11:37:@6513.4]
  wire [3:0] _T_525; // @[Lookup.scala 11:37:@6514.4]
  wire [3:0] _T_526; // @[Lookup.scala 11:37:@6515.4]
  wire [3:0] _T_527; // @[Lookup.scala 11:37:@6516.4]
  wire [3:0] _T_528; // @[Lookup.scala 11:37:@6517.4]
  wire [3:0] _T_529; // @[Lookup.scala 11:37:@6518.4]
  wire [3:0] _T_530; // @[Lookup.scala 11:37:@6519.4]
  wire [3:0] _T_531; // @[Lookup.scala 11:37:@6520.4]
  wire [3:0] _T_532; // @[Lookup.scala 11:37:@6521.4]
  wire [3:0] _T_533; // @[Lookup.scala 11:37:@6522.4]
  wire [3:0] _T_534; // @[Lookup.scala 11:37:@6523.4]
  wire [3:0] _T_535; // @[Lookup.scala 11:37:@6524.4]
  wire [3:0] _T_536; // @[Lookup.scala 11:37:@6525.4]
  wire [3:0] _T_537; // @[Lookup.scala 11:37:@6526.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:@6527.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:@6528.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:@6529.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:@6530.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:@6531.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:@6532.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:@6533.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:@6534.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:@6535.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:@6536.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:@6537.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:@6538.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:@6539.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:@6540.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:@6541.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:@6542.4]
  wire [3:0] _T_554; // @[Lookup.scala 11:37:@6543.4]
  wire [3:0] _T_555; // @[Lookup.scala 11:37:@6544.4]
  wire [3:0] _T_556; // @[Lookup.scala 11:37:@6545.4]
  wire [3:0] _T_557; // @[Lookup.scala 11:37:@6546.4]
  wire [3:0] _T_558; // @[Lookup.scala 11:37:@6547.4]
  wire [3:0] _T_559; // @[Lookup.scala 11:37:@6548.4]
  wire [1:0] _T_567; // @[Lookup.scala 11:37:@6557.4]
  wire [1:0] _T_568; // @[Lookup.scala 11:37:@6558.4]
  wire [1:0] _T_569; // @[Lookup.scala 11:37:@6559.4]
  wire [1:0] _T_570; // @[Lookup.scala 11:37:@6560.4]
  wire [1:0] _T_571; // @[Lookup.scala 11:37:@6561.4]
  wire [1:0] _T_572; // @[Lookup.scala 11:37:@6562.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@6563.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@6564.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@6565.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@6566.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@6567.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@6568.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@6569.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@6570.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@6571.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@6572.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@6573.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@6574.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@6575.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@6576.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@6577.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@6578.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@6579.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@6580.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@6581.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@6582.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@6583.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@6584.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@6585.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@6586.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@6587.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@6588.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@6589.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@6590.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@6591.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@6592.4]
  wire [1:0] _T_603; // @[Lookup.scala 11:37:@6593.4]
  wire [1:0] _T_604; // @[Lookup.scala 11:37:@6594.4]
  wire [1:0] _T_605; // @[Lookup.scala 11:37:@6595.4]
  wire [1:0] _T_606; // @[Lookup.scala 11:37:@6596.4]
  wire [1:0] _T_607; // @[Lookup.scala 11:37:@6597.4]
  wire [1:0] _T_608; // @[Lookup.scala 11:37:@6598.4]
  wire  _T_622; // @[Lookup.scala 11:37:@6613.4]
  wire  _T_623; // @[Lookup.scala 11:37:@6614.4]
  wire  _T_624; // @[Lookup.scala 11:37:@6615.4]
  wire  _T_625; // @[Lookup.scala 11:37:@6616.4]
  wire  _T_626; // @[Lookup.scala 11:37:@6617.4]
  wire  _T_627; // @[Lookup.scala 11:37:@6618.4]
  wire  _T_628; // @[Lookup.scala 11:37:@6619.4]
  wire  _T_629; // @[Lookup.scala 11:37:@6620.4]
  wire  _T_630; // @[Lookup.scala 11:37:@6621.4]
  wire  _T_631; // @[Lookup.scala 11:37:@6622.4]
  wire  _T_632; // @[Lookup.scala 11:37:@6623.4]
  wire  _T_633; // @[Lookup.scala 11:37:@6624.4]
  wire  _T_634; // @[Lookup.scala 11:37:@6625.4]
  wire  _T_635; // @[Lookup.scala 11:37:@6626.4]
  wire  _T_636; // @[Lookup.scala 11:37:@6627.4]
  wire  _T_637; // @[Lookup.scala 11:37:@6628.4]
  wire  _T_638; // @[Lookup.scala 11:37:@6629.4]
  wire  _T_639; // @[Lookup.scala 11:37:@6630.4]
  wire  _T_640; // @[Lookup.scala 11:37:@6631.4]
  wire  _T_641; // @[Lookup.scala 11:37:@6632.4]
  wire  _T_642; // @[Lookup.scala 11:37:@6633.4]
  wire  _T_643; // @[Lookup.scala 11:37:@6634.4]
  wire  _T_644; // @[Lookup.scala 11:37:@6635.4]
  wire  _T_645; // @[Lookup.scala 11:37:@6636.4]
  wire  _T_646; // @[Lookup.scala 11:37:@6637.4]
  wire  _T_647; // @[Lookup.scala 11:37:@6638.4]
  wire  _T_648; // @[Lookup.scala 11:37:@6639.4]
  wire  _T_649; // @[Lookup.scala 11:37:@6640.4]
  wire  _T_650; // @[Lookup.scala 11:37:@6641.4]
  wire  _T_651; // @[Lookup.scala 11:37:@6642.4]
  wire  _T_652; // @[Lookup.scala 11:37:@6643.4]
  wire  _T_653; // @[Lookup.scala 11:37:@6644.4]
  wire  _T_654; // @[Lookup.scala 11:37:@6645.4]
  wire  _T_655; // @[Lookup.scala 11:37:@6646.4]
  wire  _T_656; // @[Lookup.scala 11:37:@6647.4]
  wire  _T_657; // @[Lookup.scala 11:37:@6648.4]
  wire  _T_659; // @[Lookup.scala 11:37:@6651.4]
  wire  _T_660; // @[Lookup.scala 11:37:@6652.4]
  wire  _T_661; // @[Lookup.scala 11:37:@6653.4]
  wire  _T_662; // @[Lookup.scala 11:37:@6654.4]
  wire  _T_663; // @[Lookup.scala 11:37:@6655.4]
  wire  _T_664; // @[Lookup.scala 11:37:@6656.4]
  wire  _T_665; // @[Lookup.scala 11:37:@6657.4]
  wire  _T_666; // @[Lookup.scala 11:37:@6658.4]
  wire  _T_667; // @[Lookup.scala 11:37:@6659.4]
  wire  _T_668; // @[Lookup.scala 11:37:@6660.4]
  wire  _T_669; // @[Lookup.scala 11:37:@6661.4]
  wire  _T_670; // @[Lookup.scala 11:37:@6662.4]
  wire  _T_671; // @[Lookup.scala 11:37:@6663.4]
  wire  _T_672; // @[Lookup.scala 11:37:@6664.4]
  wire  _T_673; // @[Lookup.scala 11:37:@6665.4]
  wire  _T_674; // @[Lookup.scala 11:37:@6666.4]
  wire  _T_675; // @[Lookup.scala 11:37:@6667.4]
  wire  _T_676; // @[Lookup.scala 11:37:@6668.4]
  wire  _T_677; // @[Lookup.scala 11:37:@6669.4]
  wire  _T_678; // @[Lookup.scala 11:37:@6670.4]
  wire  _T_679; // @[Lookup.scala 11:37:@6671.4]
  wire  _T_680; // @[Lookup.scala 11:37:@6672.4]
  wire  _T_681; // @[Lookup.scala 11:37:@6673.4]
  wire  _T_682; // @[Lookup.scala 11:37:@6674.4]
  wire  _T_683; // @[Lookup.scala 11:37:@6675.4]
  wire  _T_684; // @[Lookup.scala 11:37:@6676.4]
  wire  _T_685; // @[Lookup.scala 11:37:@6677.4]
  wire  _T_686; // @[Lookup.scala 11:37:@6678.4]
  wire  _T_687; // @[Lookup.scala 11:37:@6679.4]
  wire  _T_688; // @[Lookup.scala 11:37:@6680.4]
  wire  _T_689; // @[Lookup.scala 11:37:@6681.4]
  wire  _T_690; // @[Lookup.scala 11:37:@6682.4]
  wire  _T_691; // @[Lookup.scala 11:37:@6683.4]
  wire  _T_692; // @[Lookup.scala 11:37:@6684.4]
  wire  _T_693; // @[Lookup.scala 11:37:@6685.4]
  wire  _T_694; // @[Lookup.scala 11:37:@6686.4]
  wire  _T_695; // @[Lookup.scala 11:37:@6687.4]
  wire  _T_696; // @[Lookup.scala 11:37:@6688.4]
  wire  _T_697; // @[Lookup.scala 11:37:@6689.4]
  wire  _T_698; // @[Lookup.scala 11:37:@6690.4]
  wire  _T_699; // @[Lookup.scala 11:37:@6691.4]
  wire  _T_700; // @[Lookup.scala 11:37:@6692.4]
  wire  _T_701; // @[Lookup.scala 11:37:@6693.4]
  wire  _T_702; // @[Lookup.scala 11:37:@6694.4]
  wire  _T_703; // @[Lookup.scala 11:37:@6695.4]
  wire  _T_704; // @[Lookup.scala 11:37:@6696.4]
  wire  _T_705; // @[Lookup.scala 11:37:@6697.4]
  wire  _T_706; // @[Lookup.scala 11:37:@6698.4]
  wire  _T_750; // @[Lookup.scala 11:37:@6743.4]
  wire  _T_751; // @[Lookup.scala 11:37:@6744.4]
  wire  _T_752; // @[Lookup.scala 11:37:@6745.4]
  wire  _T_753; // @[Lookup.scala 11:37:@6746.4]
  wire  _T_754; // @[Lookup.scala 11:37:@6747.4]
  wire  _T_755; // @[Lookup.scala 11:37:@6748.4]
  wire [2:0] _T_798; // @[Lookup.scala 11:37:@6792.4]
  wire [2:0] _T_799; // @[Lookup.scala 11:37:@6793.4]
  wire [2:0] _T_800; // @[Lookup.scala 11:37:@6794.4]
  wire [2:0] _T_801; // @[Lookup.scala 11:37:@6795.4]
  wire [2:0] _T_802; // @[Lookup.scala 11:37:@6796.4]
  wire [2:0] _T_803; // @[Lookup.scala 11:37:@6797.4]
  wire [2:0] _T_804; // @[Lookup.scala 11:37:@6798.4]
  wire [2:0] _T_808; // @[Lookup.scala 11:37:@6803.4]
  wire [2:0] _T_809; // @[Lookup.scala 11:37:@6804.4]
  wire [2:0] _T_810; // @[Lookup.scala 11:37:@6805.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@6806.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@6807.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@6808.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@6809.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@6810.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@6811.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@6812.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@6813.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@6814.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@6815.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@6816.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@6817.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@6818.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@6819.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@6820.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@6821.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@6822.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@6823.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@6824.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@6825.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@6826.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@6827.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@6828.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@6829.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@6830.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@6831.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@6832.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@6833.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@6834.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@6835.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@6836.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@6837.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@6838.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@6839.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@6840.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@6841.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@6842.4]
  wire [2:0] _T_848; // @[Lookup.scala 11:37:@6843.4]
  wire [2:0] _T_849; // @[Lookup.scala 11:37:@6844.4]
  wire [2:0] _T_850; // @[Lookup.scala 11:37:@6845.4]
  wire [2:0] _T_851; // @[Lookup.scala 11:37:@6846.4]
  wire [2:0] _T_852; // @[Lookup.scala 11:37:@6847.4]
  wire [2:0] _T_853; // @[Lookup.scala 11:37:@6848.4]
  wire [4:0] _T_905; // @[InstDecoder.scala 128:25:@6915.4]
  wire [4:0] _T_907; // @[InstDecoder.scala 130:25:@6919.4]
  wire [11:0] imm_itype; // @[InstDecoder.scala 133:27:@6921.4]
  wire [6:0] _T_908; // @[InstDecoder.scala 134:31:@6922.4]
  wire [11:0] imm_stype; // @[Cat.scala 30:58:@6924.4]
  wire  _T_910; // @[InstDecoder.scala 135:31:@6925.4]
  wire  _T_911; // @[InstDecoder.scala 135:44:@6926.4]
  wire [5:0] _T_912; // @[InstDecoder.scala 135:56:@6927.4]
  wire [3:0] _T_913; // @[InstDecoder.scala 135:73:@6928.4]
  wire [11:0] imm_sbtype; // @[Cat.scala 30:58:@6931.4]
  wire [19:0] imm_utype; // @[InstDecoder.scala 136:27:@6932.4]
  wire [7:0] _T_917; // @[InstDecoder.scala 137:44:@6934.4]
  wire  _T_918; // @[InstDecoder.scala 137:60:@6935.4]
  wire [9:0] _T_919; // @[InstDecoder.scala 137:73:@6936.4]
  wire [19:0] imm_ujtype; // @[Cat.scala 30:58:@6939.4]
  wire  _T_922; // @[InstDecoder.scala 140:43:@6940.4]
  wire [19:0] _T_926; // @[Bitwise.scala 72:12:@6942.4]
  wire  _T_928; // @[InstDecoder.scala 141:43:@6945.4]
  wire [19:0] _T_932; // @[Bitwise.scala 72:12:@6947.4]
  wire  _T_934; // @[InstDecoder.scala 142:44:@6950.4]
  wire [18:0] _T_938; // @[Bitwise.scala 72:12:@6952.4]
  wire [30:0] _T_940; // @[Cat.scala 30:58:@6953.4]
  wire  _T_948; // @[InstDecoder.scala 144:44:@6959.4]
  wire [10:0] _T_952; // @[Bitwise.scala 72:12:@6961.4]
  wire [30:0] _T_954; // @[Cat.scala 30:58:@6962.4]
  assign _T_19 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@6100.4]
  assign _T_20 = 32'h2003 == _T_19; // @[Lookup.scala 9:38:@6101.4]
  assign _T_24 = 32'h3 == _T_19; // @[Lookup.scala 9:38:@6103.4]
  assign _T_28 = 32'h4003 == _T_19; // @[Lookup.scala 9:38:@6105.4]
  assign _T_32 = 32'h1003 == _T_19; // @[Lookup.scala 9:38:@6107.4]
  assign _T_36 = 32'h5003 == _T_19; // @[Lookup.scala 9:38:@6109.4]
  assign _T_40 = 32'h2023 == _T_19; // @[Lookup.scala 9:38:@6111.4]
  assign _T_44 = 32'h23 == _T_19; // @[Lookup.scala 9:38:@6113.4]
  assign _T_48 = 32'h1023 == _T_19; // @[Lookup.scala 9:38:@6115.4]
  assign _T_51 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@6116.4]
  assign _T_52 = 32'h17 == _T_51; // @[Lookup.scala 9:38:@6117.4]
  assign _T_56 = 32'h37 == _T_51; // @[Lookup.scala 9:38:@6119.4]
  assign _T_60 = 32'h13 == _T_19; // @[Lookup.scala 9:38:@6121.4]
  assign _T_64 = 32'h7013 == _T_19; // @[Lookup.scala 9:38:@6123.4]
  assign _T_68 = 32'h6013 == _T_19; // @[Lookup.scala 9:38:@6125.4]
  assign _T_72 = 32'h4013 == _T_19; // @[Lookup.scala 9:38:@6127.4]
  assign _T_76 = 32'h2013 == _T_19; // @[Lookup.scala 9:38:@6129.4]
  assign _T_80 = 32'h3013 == _T_19; // @[Lookup.scala 9:38:@6131.4]
  assign _T_83 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@6132.4]
  assign _T_84 = 32'h1013 == _T_83; // @[Lookup.scala 9:38:@6133.4]
  assign _T_88 = 32'h40005013 == _T_83; // @[Lookup.scala 9:38:@6135.4]
  assign _T_92 = 32'h5013 == _T_83; // @[Lookup.scala 9:38:@6137.4]
  assign _T_95 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@6138.4]
  assign _T_96 = 32'h1033 == _T_95; // @[Lookup.scala 9:38:@6139.4]
  assign _T_100 = 32'h33 == _T_95; // @[Lookup.scala 9:38:@6141.4]
  assign _T_104 = 32'h40000033 == _T_95; // @[Lookup.scala 9:38:@6143.4]
  assign _T_108 = 32'h2033 == _T_95; // @[Lookup.scala 9:38:@6145.4]
  assign _T_112 = 32'h3033 == _T_95; // @[Lookup.scala 9:38:@6147.4]
  assign _T_116 = 32'h7033 == _T_95; // @[Lookup.scala 9:38:@6149.4]
  assign _T_120 = 32'h6033 == _T_95; // @[Lookup.scala 9:38:@6151.4]
  assign _T_124 = 32'h4033 == _T_95; // @[Lookup.scala 9:38:@6153.4]
  assign _T_128 = 32'h40005033 == _T_95; // @[Lookup.scala 9:38:@6155.4]
  assign _T_132 = 32'h5033 == _T_95; // @[Lookup.scala 9:38:@6157.4]
  assign _T_136 = 32'h6f == _T_51; // @[Lookup.scala 9:38:@6159.4]
  assign _T_140 = 32'h67 == _T_19; // @[Lookup.scala 9:38:@6161.4]
  assign _T_144 = 32'h63 == _T_19; // @[Lookup.scala 9:38:@6163.4]
  assign _T_148 = 32'h1063 == _T_19; // @[Lookup.scala 9:38:@6165.4]
  assign _T_152 = 32'h5063 == _T_19; // @[Lookup.scala 9:38:@6167.4]
  assign _T_156 = 32'h7063 == _T_19; // @[Lookup.scala 9:38:@6169.4]
  assign _T_160 = 32'h4063 == _T_19; // @[Lookup.scala 9:38:@6171.4]
  assign _T_164 = 32'h6063 == _T_19; // @[Lookup.scala 9:38:@6173.4]
  assign _T_168 = 32'h5073 == _T_19; // @[Lookup.scala 9:38:@6175.4]
  assign _T_172 = 32'h6073 == _T_19; // @[Lookup.scala 9:38:@6177.4]
  assign _T_176 = 32'h1073 == _T_19; // @[Lookup.scala 9:38:@6179.4]
  assign _T_180 = 32'h2073 == _T_19; // @[Lookup.scala 9:38:@6181.4]
  assign _T_184 = 32'h3073 == _T_19; // @[Lookup.scala 9:38:@6183.4]
  assign _T_188 = 32'h7073 == _T_19; // @[Lookup.scala 9:38:@6185.4]
  assign _T_192 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@6187.4]
  assign _T_196 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@6189.4]
  assign _T_200 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@6191.4]
  assign _T_204 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@6193.4]
  assign _T_208 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@6195.4]
  assign _T_212 = 32'h100f == _T_19; // @[Lookup.scala 9:38:@6197.4]
  assign _T_216 = 32'hf == _T_19; // @[Lookup.scala 9:38:@6199.4]
  assign _T_218 = _T_212 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@6201.4]
  assign _T_219 = _T_208 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@6202.4]
  assign _T_220 = _T_204 ? 1'h1 : _T_219; // @[Lookup.scala 11:37:@6203.4]
  assign _T_221 = _T_200 ? 1'h1 : _T_220; // @[Lookup.scala 11:37:@6204.4]
  assign _T_222 = _T_196 ? 1'h1 : _T_221; // @[Lookup.scala 11:37:@6205.4]
  assign _T_223 = _T_192 ? 1'h1 : _T_222; // @[Lookup.scala 11:37:@6206.4]
  assign _T_224 = _T_188 ? 1'h1 : _T_223; // @[Lookup.scala 11:37:@6207.4]
  assign _T_225 = _T_184 ? 1'h1 : _T_224; // @[Lookup.scala 11:37:@6208.4]
  assign _T_226 = _T_180 ? 1'h1 : _T_225; // @[Lookup.scala 11:37:@6209.4]
  assign _T_227 = _T_176 ? 1'h1 : _T_226; // @[Lookup.scala 11:37:@6210.4]
  assign _T_228 = _T_172 ? 1'h1 : _T_227; // @[Lookup.scala 11:37:@6211.4]
  assign _T_229 = _T_168 ? 1'h1 : _T_228; // @[Lookup.scala 11:37:@6212.4]
  assign _T_230 = _T_164 ? 1'h1 : _T_229; // @[Lookup.scala 11:37:@6213.4]
  assign _T_231 = _T_160 ? 1'h1 : _T_230; // @[Lookup.scala 11:37:@6214.4]
  assign _T_232 = _T_156 ? 1'h1 : _T_231; // @[Lookup.scala 11:37:@6215.4]
  assign _T_233 = _T_152 ? 1'h1 : _T_232; // @[Lookup.scala 11:37:@6216.4]
  assign _T_234 = _T_148 ? 1'h1 : _T_233; // @[Lookup.scala 11:37:@6217.4]
  assign _T_235 = _T_144 ? 1'h1 : _T_234; // @[Lookup.scala 11:37:@6218.4]
  assign _T_236 = _T_140 ? 1'h1 : _T_235; // @[Lookup.scala 11:37:@6219.4]
  assign _T_237 = _T_136 ? 1'h1 : _T_236; // @[Lookup.scala 11:37:@6220.4]
  assign _T_238 = _T_132 ? 1'h1 : _T_237; // @[Lookup.scala 11:37:@6221.4]
  assign _T_239 = _T_128 ? 1'h1 : _T_238; // @[Lookup.scala 11:37:@6222.4]
  assign _T_240 = _T_124 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@6223.4]
  assign _T_241 = _T_120 ? 1'h1 : _T_240; // @[Lookup.scala 11:37:@6224.4]
  assign _T_242 = _T_116 ? 1'h1 : _T_241; // @[Lookup.scala 11:37:@6225.4]
  assign _T_243 = _T_112 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@6226.4]
  assign _T_244 = _T_108 ? 1'h1 : _T_243; // @[Lookup.scala 11:37:@6227.4]
  assign _T_245 = _T_104 ? 1'h1 : _T_244; // @[Lookup.scala 11:37:@6228.4]
  assign _T_246 = _T_100 ? 1'h1 : _T_245; // @[Lookup.scala 11:37:@6229.4]
  assign _T_247 = _T_96 ? 1'h1 : _T_246; // @[Lookup.scala 11:37:@6230.4]
  assign _T_248 = _T_92 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@6231.4]
  assign _T_249 = _T_88 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@6232.4]
  assign _T_250 = _T_84 ? 1'h1 : _T_249; // @[Lookup.scala 11:37:@6233.4]
  assign _T_251 = _T_80 ? 1'h1 : _T_250; // @[Lookup.scala 11:37:@6234.4]
  assign _T_252 = _T_76 ? 1'h1 : _T_251; // @[Lookup.scala 11:37:@6235.4]
  assign _T_253 = _T_72 ? 1'h1 : _T_252; // @[Lookup.scala 11:37:@6236.4]
  assign _T_254 = _T_68 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@6237.4]
  assign _T_255 = _T_64 ? 1'h1 : _T_254; // @[Lookup.scala 11:37:@6238.4]
  assign _T_256 = _T_60 ? 1'h1 : _T_255; // @[Lookup.scala 11:37:@6239.4]
  assign _T_257 = _T_56 ? 1'h1 : _T_256; // @[Lookup.scala 11:37:@6240.4]
  assign _T_258 = _T_52 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:@6241.4]
  assign _T_259 = _T_48 ? 1'h1 : _T_258; // @[Lookup.scala 11:37:@6242.4]
  assign _T_260 = _T_44 ? 1'h1 : _T_259; // @[Lookup.scala 11:37:@6243.4]
  assign _T_261 = _T_40 ? 1'h1 : _T_260; // @[Lookup.scala 11:37:@6244.4]
  assign _T_262 = _T_36 ? 1'h1 : _T_261; // @[Lookup.scala 11:37:@6245.4]
  assign _T_263 = _T_32 ? 1'h1 : _T_262; // @[Lookup.scala 11:37:@6246.4]
  assign _T_264 = _T_28 ? 1'h1 : _T_263; // @[Lookup.scala 11:37:@6247.4]
  assign _T_265 = _T_24 ? 1'h1 : _T_264; // @[Lookup.scala 11:37:@6248.4]
  assign signals_0 = _T_20 ? 1'h1 : _T_265; // @[Lookup.scala 11:37:@6249.4]
  assign _T_279 = _T_164 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@6263.4]
  assign _T_280 = _T_160 ? 4'h5 : _T_279; // @[Lookup.scala 11:37:@6264.4]
  assign _T_281 = _T_156 ? 4'h4 : _T_280; // @[Lookup.scala 11:37:@6265.4]
  assign _T_282 = _T_152 ? 4'h3 : _T_281; // @[Lookup.scala 11:37:@6266.4]
  assign _T_283 = _T_148 ? 4'h1 : _T_282; // @[Lookup.scala 11:37:@6267.4]
  assign _T_284 = _T_144 ? 4'h2 : _T_283; // @[Lookup.scala 11:37:@6268.4]
  assign _T_285 = _T_140 ? 4'h8 : _T_284; // @[Lookup.scala 11:37:@6269.4]
  assign _T_286 = _T_136 ? 4'h7 : _T_285; // @[Lookup.scala 11:37:@6270.4]
  assign _T_287 = _T_132 ? 4'h0 : _T_286; // @[Lookup.scala 11:37:@6271.4]
  assign _T_288 = _T_128 ? 4'h0 : _T_287; // @[Lookup.scala 11:37:@6272.4]
  assign _T_289 = _T_124 ? 4'h0 : _T_288; // @[Lookup.scala 11:37:@6273.4]
  assign _T_290 = _T_120 ? 4'h0 : _T_289; // @[Lookup.scala 11:37:@6274.4]
  assign _T_291 = _T_116 ? 4'h0 : _T_290; // @[Lookup.scala 11:37:@6275.4]
  assign _T_292 = _T_112 ? 4'h0 : _T_291; // @[Lookup.scala 11:37:@6276.4]
  assign _T_293 = _T_108 ? 4'h0 : _T_292; // @[Lookup.scala 11:37:@6277.4]
  assign _T_294 = _T_104 ? 4'h0 : _T_293; // @[Lookup.scala 11:37:@6278.4]
  assign _T_295 = _T_100 ? 4'h0 : _T_294; // @[Lookup.scala 11:37:@6279.4]
  assign _T_296 = _T_96 ? 4'h0 : _T_295; // @[Lookup.scala 11:37:@6280.4]
  assign _T_297 = _T_92 ? 4'h0 : _T_296; // @[Lookup.scala 11:37:@6281.4]
  assign _T_298 = _T_88 ? 4'h0 : _T_297; // @[Lookup.scala 11:37:@6282.4]
  assign _T_299 = _T_84 ? 4'h0 : _T_298; // @[Lookup.scala 11:37:@6283.4]
  assign _T_300 = _T_80 ? 4'h0 : _T_299; // @[Lookup.scala 11:37:@6284.4]
  assign _T_301 = _T_76 ? 4'h0 : _T_300; // @[Lookup.scala 11:37:@6285.4]
  assign _T_302 = _T_72 ? 4'h0 : _T_301; // @[Lookup.scala 11:37:@6286.4]
  assign _T_303 = _T_68 ? 4'h0 : _T_302; // @[Lookup.scala 11:37:@6287.4]
  assign _T_304 = _T_64 ? 4'h0 : _T_303; // @[Lookup.scala 11:37:@6288.4]
  assign _T_305 = _T_60 ? 4'h0 : _T_304; // @[Lookup.scala 11:37:@6289.4]
  assign _T_306 = _T_56 ? 4'h0 : _T_305; // @[Lookup.scala 11:37:@6290.4]
  assign _T_307 = _T_52 ? 4'h0 : _T_306; // @[Lookup.scala 11:37:@6291.4]
  assign _T_308 = _T_48 ? 4'h0 : _T_307; // @[Lookup.scala 11:37:@6292.4]
  assign _T_309 = _T_44 ? 4'h0 : _T_308; // @[Lookup.scala 11:37:@6293.4]
  assign _T_310 = _T_40 ? 4'h0 : _T_309; // @[Lookup.scala 11:37:@6294.4]
  assign _T_311 = _T_36 ? 4'h0 : _T_310; // @[Lookup.scala 11:37:@6295.4]
  assign _T_312 = _T_32 ? 4'h0 : _T_311; // @[Lookup.scala 11:37:@6296.4]
  assign _T_313 = _T_28 ? 4'h0 : _T_312; // @[Lookup.scala 11:37:@6297.4]
  assign _T_314 = _T_24 ? 4'h0 : _T_313; // @[Lookup.scala 11:37:@6298.4]
  assign _T_322 = _T_188 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@6307.4]
  assign _T_323 = _T_184 ? 2'h0 : _T_322; // @[Lookup.scala 11:37:@6308.4]
  assign _T_324 = _T_180 ? 2'h0 : _T_323; // @[Lookup.scala 11:37:@6309.4]
  assign _T_325 = _T_176 ? 2'h0 : _T_324; // @[Lookup.scala 11:37:@6310.4]
  assign _T_326 = _T_172 ? 2'h2 : _T_325; // @[Lookup.scala 11:37:@6311.4]
  assign _T_327 = _T_168 ? 2'h2 : _T_326; // @[Lookup.scala 11:37:@6312.4]
  assign _T_328 = _T_164 ? 2'h0 : _T_327; // @[Lookup.scala 11:37:@6313.4]
  assign _T_329 = _T_160 ? 2'h0 : _T_328; // @[Lookup.scala 11:37:@6314.4]
  assign _T_330 = _T_156 ? 2'h0 : _T_329; // @[Lookup.scala 11:37:@6315.4]
  assign _T_331 = _T_152 ? 2'h0 : _T_330; // @[Lookup.scala 11:37:@6316.4]
  assign _T_332 = _T_148 ? 2'h0 : _T_331; // @[Lookup.scala 11:37:@6317.4]
  assign _T_333 = _T_144 ? 2'h0 : _T_332; // @[Lookup.scala 11:37:@6318.4]
  assign _T_334 = _T_140 ? 2'h0 : _T_333; // @[Lookup.scala 11:37:@6319.4]
  assign _T_335 = _T_136 ? 2'h0 : _T_334; // @[Lookup.scala 11:37:@6320.4]
  assign _T_336 = _T_132 ? 2'h0 : _T_335; // @[Lookup.scala 11:37:@6321.4]
  assign _T_337 = _T_128 ? 2'h0 : _T_336; // @[Lookup.scala 11:37:@6322.4]
  assign _T_338 = _T_124 ? 2'h0 : _T_337; // @[Lookup.scala 11:37:@6323.4]
  assign _T_339 = _T_120 ? 2'h0 : _T_338; // @[Lookup.scala 11:37:@6324.4]
  assign _T_340 = _T_116 ? 2'h0 : _T_339; // @[Lookup.scala 11:37:@6325.4]
  assign _T_341 = _T_112 ? 2'h0 : _T_340; // @[Lookup.scala 11:37:@6326.4]
  assign _T_342 = _T_108 ? 2'h0 : _T_341; // @[Lookup.scala 11:37:@6327.4]
  assign _T_343 = _T_104 ? 2'h0 : _T_342; // @[Lookup.scala 11:37:@6328.4]
  assign _T_344 = _T_100 ? 2'h0 : _T_343; // @[Lookup.scala 11:37:@6329.4]
  assign _T_345 = _T_96 ? 2'h0 : _T_344; // @[Lookup.scala 11:37:@6330.4]
  assign _T_346 = _T_92 ? 2'h0 : _T_345; // @[Lookup.scala 11:37:@6331.4]
  assign _T_347 = _T_88 ? 2'h0 : _T_346; // @[Lookup.scala 11:37:@6332.4]
  assign _T_348 = _T_84 ? 2'h0 : _T_347; // @[Lookup.scala 11:37:@6333.4]
  assign _T_349 = _T_80 ? 2'h0 : _T_348; // @[Lookup.scala 11:37:@6334.4]
  assign _T_350 = _T_76 ? 2'h0 : _T_349; // @[Lookup.scala 11:37:@6335.4]
  assign _T_351 = _T_72 ? 2'h0 : _T_350; // @[Lookup.scala 11:37:@6336.4]
  assign _T_352 = _T_68 ? 2'h0 : _T_351; // @[Lookup.scala 11:37:@6337.4]
  assign _T_353 = _T_64 ? 2'h0 : _T_352; // @[Lookup.scala 11:37:@6338.4]
  assign _T_354 = _T_60 ? 2'h0 : _T_353; // @[Lookup.scala 11:37:@6339.4]
  assign _T_355 = _T_56 ? 2'h0 : _T_354; // @[Lookup.scala 11:37:@6340.4]
  assign _T_356 = _T_52 ? 2'h1 : _T_355; // @[Lookup.scala 11:37:@6341.4]
  assign _T_357 = _T_48 ? 2'h0 : _T_356; // @[Lookup.scala 11:37:@6342.4]
  assign _T_358 = _T_44 ? 2'h0 : _T_357; // @[Lookup.scala 11:37:@6343.4]
  assign _T_359 = _T_40 ? 2'h0 : _T_358; // @[Lookup.scala 11:37:@6344.4]
  assign _T_360 = _T_36 ? 2'h0 : _T_359; // @[Lookup.scala 11:37:@6345.4]
  assign _T_361 = _T_32 ? 2'h0 : _T_360; // @[Lookup.scala 11:37:@6346.4]
  assign _T_362 = _T_28 ? 2'h0 : _T_361; // @[Lookup.scala 11:37:@6347.4]
  assign _T_363 = _T_24 ? 2'h0 : _T_362; // @[Lookup.scala 11:37:@6348.4]
  assign _T_377 = _T_164 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37:@6363.4]
  assign _T_378 = _T_160 ? 3'h3 : _T_377; // @[Lookup.scala 11:37:@6364.4]
  assign _T_379 = _T_156 ? 3'h3 : _T_378; // @[Lookup.scala 11:37:@6365.4]
  assign _T_380 = _T_152 ? 3'h3 : _T_379; // @[Lookup.scala 11:37:@6366.4]
  assign _T_381 = _T_148 ? 3'h3 : _T_380; // @[Lookup.scala 11:37:@6367.4]
  assign _T_382 = _T_144 ? 3'h3 : _T_381; // @[Lookup.scala 11:37:@6368.4]
  assign _T_383 = _T_140 ? 3'h1 : _T_382; // @[Lookup.scala 11:37:@6369.4]
  assign _T_384 = _T_136 ? 3'h5 : _T_383; // @[Lookup.scala 11:37:@6370.4]
  assign _T_385 = _T_132 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@6371.4]
  assign _T_386 = _T_128 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@6372.4]
  assign _T_387 = _T_124 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@6373.4]
  assign _T_388 = _T_120 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@6374.4]
  assign _T_389 = _T_116 ? 3'h0 : _T_388; // @[Lookup.scala 11:37:@6375.4]
  assign _T_390 = _T_112 ? 3'h0 : _T_389; // @[Lookup.scala 11:37:@6376.4]
  assign _T_391 = _T_108 ? 3'h0 : _T_390; // @[Lookup.scala 11:37:@6377.4]
  assign _T_392 = _T_104 ? 3'h0 : _T_391; // @[Lookup.scala 11:37:@6378.4]
  assign _T_393 = _T_100 ? 3'h0 : _T_392; // @[Lookup.scala 11:37:@6379.4]
  assign _T_394 = _T_96 ? 3'h0 : _T_393; // @[Lookup.scala 11:37:@6380.4]
  assign _T_395 = _T_92 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@6381.4]
  assign _T_396 = _T_88 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@6382.4]
  assign _T_397 = _T_84 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@6383.4]
  assign _T_398 = _T_80 ? 3'h1 : _T_397; // @[Lookup.scala 11:37:@6384.4]
  assign _T_399 = _T_76 ? 3'h1 : _T_398; // @[Lookup.scala 11:37:@6385.4]
  assign _T_400 = _T_72 ? 3'h1 : _T_399; // @[Lookup.scala 11:37:@6386.4]
  assign _T_401 = _T_68 ? 3'h1 : _T_400; // @[Lookup.scala 11:37:@6387.4]
  assign _T_402 = _T_64 ? 3'h1 : _T_401; // @[Lookup.scala 11:37:@6388.4]
  assign _T_403 = _T_60 ? 3'h1 : _T_402; // @[Lookup.scala 11:37:@6389.4]
  assign _T_404 = _T_56 ? 3'h4 : _T_403; // @[Lookup.scala 11:37:@6390.4]
  assign _T_405 = _T_52 ? 3'h4 : _T_404; // @[Lookup.scala 11:37:@6391.4]
  assign _T_406 = _T_48 ? 3'h2 : _T_405; // @[Lookup.scala 11:37:@6392.4]
  assign _T_407 = _T_44 ? 3'h2 : _T_406; // @[Lookup.scala 11:37:@6393.4]
  assign _T_408 = _T_40 ? 3'h2 : _T_407; // @[Lookup.scala 11:37:@6394.4]
  assign _T_409 = _T_36 ? 3'h1 : _T_408; // @[Lookup.scala 11:37:@6395.4]
  assign _T_410 = _T_32 ? 3'h1 : _T_409; // @[Lookup.scala 11:37:@6396.4]
  assign _T_411 = _T_28 ? 3'h1 : _T_410; // @[Lookup.scala 11:37:@6397.4]
  assign _T_412 = _T_24 ? 3'h1 : _T_411; // @[Lookup.scala 11:37:@6398.4]
  assign _T_421 = _T_184 ? 1'h1 : _T_188; // @[Lookup.scala 11:37:@6408.4]
  assign _T_422 = _T_180 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@6409.4]
  assign _T_423 = _T_176 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@6410.4]
  assign _T_424 = _T_172 ? 1'h1 : _T_423; // @[Lookup.scala 11:37:@6411.4]
  assign _T_425 = _T_168 ? 1'h1 : _T_424; // @[Lookup.scala 11:37:@6412.4]
  assign _T_426 = _T_164 ? 1'h1 : _T_425; // @[Lookup.scala 11:37:@6413.4]
  assign _T_427 = _T_160 ? 1'h1 : _T_426; // @[Lookup.scala 11:37:@6414.4]
  assign _T_428 = _T_156 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@6415.4]
  assign _T_429 = _T_152 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@6416.4]
  assign _T_430 = _T_148 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@6417.4]
  assign _T_431 = _T_144 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@6418.4]
  assign _T_432 = _T_140 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@6419.4]
  assign _T_433 = _T_136 ? 1'h0 : _T_432; // @[Lookup.scala 11:37:@6420.4]
  assign _T_434 = _T_132 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@6421.4]
  assign _T_435 = _T_128 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@6422.4]
  assign _T_436 = _T_124 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@6423.4]
  assign _T_437 = _T_120 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@6424.4]
  assign _T_438 = _T_116 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@6425.4]
  assign _T_439 = _T_112 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@6426.4]
  assign _T_440 = _T_108 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@6427.4]
  assign _T_441 = _T_104 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@6428.4]
  assign _T_442 = _T_100 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@6429.4]
  assign _T_443 = _T_96 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@6430.4]
  assign _T_444 = _T_92 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@6431.4]
  assign _T_445 = _T_88 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@6432.4]
  assign _T_446 = _T_84 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@6433.4]
  assign _T_447 = _T_80 ? 1'h1 : _T_446; // @[Lookup.scala 11:37:@6434.4]
  assign _T_448 = _T_76 ? 1'h1 : _T_447; // @[Lookup.scala 11:37:@6435.4]
  assign _T_449 = _T_72 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@6436.4]
  assign _T_450 = _T_68 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@6437.4]
  assign _T_451 = _T_64 ? 1'h1 : _T_450; // @[Lookup.scala 11:37:@6438.4]
  assign _T_452 = _T_60 ? 1'h1 : _T_451; // @[Lookup.scala 11:37:@6439.4]
  assign _T_453 = _T_56 ? 1'h0 : _T_452; // @[Lookup.scala 11:37:@6440.4]
  assign _T_454 = _T_52 ? 1'h0 : _T_453; // @[Lookup.scala 11:37:@6441.4]
  assign _T_455 = _T_48 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@6442.4]
  assign _T_456 = _T_44 ? 1'h1 : _T_455; // @[Lookup.scala 11:37:@6443.4]
  assign _T_457 = _T_40 ? 1'h1 : _T_456; // @[Lookup.scala 11:37:@6444.4]
  assign _T_458 = _T_36 ? 1'h1 : _T_457; // @[Lookup.scala 11:37:@6445.4]
  assign _T_459 = _T_32 ? 1'h1 : _T_458; // @[Lookup.scala 11:37:@6446.4]
  assign _T_460 = _T_28 ? 1'h1 : _T_459; // @[Lookup.scala 11:37:@6447.4]
  assign _T_461 = _T_24 ? 1'h1 : _T_460; // @[Lookup.scala 11:37:@6448.4]
  assign _T_481 = _T_140 ? 1'h0 : _T_431; // @[Lookup.scala 11:37:@6469.4]
  assign _T_482 = _T_136 ? 1'h0 : _T_481; // @[Lookup.scala 11:37:@6470.4]
  assign _T_483 = _T_132 ? 1'h1 : _T_482; // @[Lookup.scala 11:37:@6471.4]
  assign _T_484 = _T_128 ? 1'h1 : _T_483; // @[Lookup.scala 11:37:@6472.4]
  assign _T_485 = _T_124 ? 1'h1 : _T_484; // @[Lookup.scala 11:37:@6473.4]
  assign _T_486 = _T_120 ? 1'h1 : _T_485; // @[Lookup.scala 11:37:@6474.4]
  assign _T_487 = _T_116 ? 1'h1 : _T_486; // @[Lookup.scala 11:37:@6475.4]
  assign _T_488 = _T_112 ? 1'h1 : _T_487; // @[Lookup.scala 11:37:@6476.4]
  assign _T_489 = _T_108 ? 1'h1 : _T_488; // @[Lookup.scala 11:37:@6477.4]
  assign _T_490 = _T_104 ? 1'h1 : _T_489; // @[Lookup.scala 11:37:@6478.4]
  assign _T_491 = _T_100 ? 1'h1 : _T_490; // @[Lookup.scala 11:37:@6479.4]
  assign _T_492 = _T_96 ? 1'h1 : _T_491; // @[Lookup.scala 11:37:@6480.4]
  assign _T_493 = _T_92 ? 1'h0 : _T_492; // @[Lookup.scala 11:37:@6481.4]
  assign _T_494 = _T_88 ? 1'h0 : _T_493; // @[Lookup.scala 11:37:@6482.4]
  assign _T_495 = _T_84 ? 1'h0 : _T_494; // @[Lookup.scala 11:37:@6483.4]
  assign _T_496 = _T_80 ? 1'h0 : _T_495; // @[Lookup.scala 11:37:@6484.4]
  assign _T_497 = _T_76 ? 1'h0 : _T_496; // @[Lookup.scala 11:37:@6485.4]
  assign _T_498 = _T_72 ? 1'h0 : _T_497; // @[Lookup.scala 11:37:@6486.4]
  assign _T_499 = _T_68 ? 1'h0 : _T_498; // @[Lookup.scala 11:37:@6487.4]
  assign _T_500 = _T_64 ? 1'h0 : _T_499; // @[Lookup.scala 11:37:@6488.4]
  assign _T_501 = _T_60 ? 1'h0 : _T_500; // @[Lookup.scala 11:37:@6489.4]
  assign _T_502 = _T_56 ? 1'h0 : _T_501; // @[Lookup.scala 11:37:@6490.4]
  assign _T_503 = _T_52 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@6491.4]
  assign _T_504 = _T_48 ? 1'h1 : _T_503; // @[Lookup.scala 11:37:@6492.4]
  assign _T_505 = _T_44 ? 1'h1 : _T_504; // @[Lookup.scala 11:37:@6493.4]
  assign _T_506 = _T_40 ? 1'h1 : _T_505; // @[Lookup.scala 11:37:@6494.4]
  assign _T_507 = _T_36 ? 1'h0 : _T_506; // @[Lookup.scala 11:37:@6495.4]
  assign _T_508 = _T_32 ? 1'h0 : _T_507; // @[Lookup.scala 11:37:@6496.4]
  assign _T_509 = _T_28 ? 1'h0 : _T_508; // @[Lookup.scala 11:37:@6497.4]
  assign _T_510 = _T_24 ? 1'h0 : _T_509; // @[Lookup.scala 11:37:@6498.4]
  assign _T_518 = _T_188 ? 4'ha : 4'h0; // @[Lookup.scala 11:37:@6507.4]
  assign _T_519 = _T_184 ? 4'ha : _T_518; // @[Lookup.scala 11:37:@6508.4]
  assign _T_520 = _T_180 ? 4'ha : _T_519; // @[Lookup.scala 11:37:@6509.4]
  assign _T_521 = _T_176 ? 4'ha : _T_520; // @[Lookup.scala 11:37:@6510.4]
  assign _T_522 = _T_172 ? 4'ha : _T_521; // @[Lookup.scala 11:37:@6511.4]
  assign _T_523 = _T_168 ? 4'ha : _T_522; // @[Lookup.scala 11:37:@6512.4]
  assign _T_524 = _T_164 ? 4'h0 : _T_523; // @[Lookup.scala 11:37:@6513.4]
  assign _T_525 = _T_160 ? 4'h0 : _T_524; // @[Lookup.scala 11:37:@6514.4]
  assign _T_526 = _T_156 ? 4'h0 : _T_525; // @[Lookup.scala 11:37:@6515.4]
  assign _T_527 = _T_152 ? 4'h0 : _T_526; // @[Lookup.scala 11:37:@6516.4]
  assign _T_528 = _T_148 ? 4'h0 : _T_527; // @[Lookup.scala 11:37:@6517.4]
  assign _T_529 = _T_144 ? 4'h0 : _T_528; // @[Lookup.scala 11:37:@6518.4]
  assign _T_530 = _T_140 ? 4'h0 : _T_529; // @[Lookup.scala 11:37:@6519.4]
  assign _T_531 = _T_136 ? 4'h0 : _T_530; // @[Lookup.scala 11:37:@6520.4]
  assign _T_532 = _T_132 ? 4'h3 : _T_531; // @[Lookup.scala 11:37:@6521.4]
  assign _T_533 = _T_128 ? 4'h4 : _T_532; // @[Lookup.scala 11:37:@6522.4]
  assign _T_534 = _T_124 ? 4'h7 : _T_533; // @[Lookup.scala 11:37:@6523.4]
  assign _T_535 = _T_120 ? 4'h6 : _T_534; // @[Lookup.scala 11:37:@6524.4]
  assign _T_536 = _T_116 ? 4'h5 : _T_535; // @[Lookup.scala 11:37:@6525.4]
  assign _T_537 = _T_112 ? 4'h9 : _T_536; // @[Lookup.scala 11:37:@6526.4]
  assign _T_538 = _T_108 ? 4'h8 : _T_537; // @[Lookup.scala 11:37:@6527.4]
  assign _T_539 = _T_104 ? 4'h1 : _T_538; // @[Lookup.scala 11:37:@6528.4]
  assign _T_540 = _T_100 ? 4'h0 : _T_539; // @[Lookup.scala 11:37:@6529.4]
  assign _T_541 = _T_96 ? 4'h2 : _T_540; // @[Lookup.scala 11:37:@6530.4]
  assign _T_542 = _T_92 ? 4'h3 : _T_541; // @[Lookup.scala 11:37:@6531.4]
  assign _T_543 = _T_88 ? 4'h4 : _T_542; // @[Lookup.scala 11:37:@6532.4]
  assign _T_544 = _T_84 ? 4'h2 : _T_543; // @[Lookup.scala 11:37:@6533.4]
  assign _T_545 = _T_80 ? 4'h9 : _T_544; // @[Lookup.scala 11:37:@6534.4]
  assign _T_546 = _T_76 ? 4'h8 : _T_545; // @[Lookup.scala 11:37:@6535.4]
  assign _T_547 = _T_72 ? 4'h7 : _T_546; // @[Lookup.scala 11:37:@6536.4]
  assign _T_548 = _T_68 ? 4'h6 : _T_547; // @[Lookup.scala 11:37:@6537.4]
  assign _T_549 = _T_64 ? 4'h5 : _T_548; // @[Lookup.scala 11:37:@6538.4]
  assign _T_550 = _T_60 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:@6539.4]
  assign _T_551 = _T_56 ? 4'hb : _T_550; // @[Lookup.scala 11:37:@6540.4]
  assign _T_552 = _T_52 ? 4'h0 : _T_551; // @[Lookup.scala 11:37:@6541.4]
  assign _T_553 = _T_48 ? 4'h0 : _T_552; // @[Lookup.scala 11:37:@6542.4]
  assign _T_554 = _T_44 ? 4'h0 : _T_553; // @[Lookup.scala 11:37:@6543.4]
  assign _T_555 = _T_40 ? 4'h0 : _T_554; // @[Lookup.scala 11:37:@6544.4]
  assign _T_556 = _T_36 ? 4'h0 : _T_555; // @[Lookup.scala 11:37:@6545.4]
  assign _T_557 = _T_32 ? 4'h0 : _T_556; // @[Lookup.scala 11:37:@6546.4]
  assign _T_558 = _T_28 ? 4'h0 : _T_557; // @[Lookup.scala 11:37:@6547.4]
  assign _T_559 = _T_24 ? 4'h0 : _T_558; // @[Lookup.scala 11:37:@6548.4]
  assign _T_567 = _T_188 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@6557.4]
  assign _T_568 = _T_184 ? 2'h3 : _T_567; // @[Lookup.scala 11:37:@6558.4]
  assign _T_569 = _T_180 ? 2'h3 : _T_568; // @[Lookup.scala 11:37:@6559.4]
  assign _T_570 = _T_176 ? 2'h3 : _T_569; // @[Lookup.scala 11:37:@6560.4]
  assign _T_571 = _T_172 ? 2'h3 : _T_570; // @[Lookup.scala 11:37:@6561.4]
  assign _T_572 = _T_168 ? 2'h3 : _T_571; // @[Lookup.scala 11:37:@6562.4]
  assign _T_573 = _T_164 ? 2'h0 : _T_572; // @[Lookup.scala 11:37:@6563.4]
  assign _T_574 = _T_160 ? 2'h0 : _T_573; // @[Lookup.scala 11:37:@6564.4]
  assign _T_575 = _T_156 ? 2'h0 : _T_574; // @[Lookup.scala 11:37:@6565.4]
  assign _T_576 = _T_152 ? 2'h0 : _T_575; // @[Lookup.scala 11:37:@6566.4]
  assign _T_577 = _T_148 ? 2'h0 : _T_576; // @[Lookup.scala 11:37:@6567.4]
  assign _T_578 = _T_144 ? 2'h0 : _T_577; // @[Lookup.scala 11:37:@6568.4]
  assign _T_579 = _T_140 ? 2'h2 : _T_578; // @[Lookup.scala 11:37:@6569.4]
  assign _T_580 = _T_136 ? 2'h2 : _T_579; // @[Lookup.scala 11:37:@6570.4]
  assign _T_581 = _T_132 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@6571.4]
  assign _T_582 = _T_128 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@6572.4]
  assign _T_583 = _T_124 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@6573.4]
  assign _T_584 = _T_120 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@6574.4]
  assign _T_585 = _T_116 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@6575.4]
  assign _T_586 = _T_112 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@6576.4]
  assign _T_587 = _T_108 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@6577.4]
  assign _T_588 = _T_104 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@6578.4]
  assign _T_589 = _T_100 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@6579.4]
  assign _T_590 = _T_96 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@6580.4]
  assign _T_591 = _T_92 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@6581.4]
  assign _T_592 = _T_88 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@6582.4]
  assign _T_593 = _T_84 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@6583.4]
  assign _T_594 = _T_80 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@6584.4]
  assign _T_595 = _T_76 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@6585.4]
  assign _T_596 = _T_72 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@6586.4]
  assign _T_597 = _T_68 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@6587.4]
  assign _T_598 = _T_64 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@6588.4]
  assign _T_599 = _T_60 ? 2'h0 : _T_598; // @[Lookup.scala 11:37:@6589.4]
  assign _T_600 = _T_56 ? 2'h0 : _T_599; // @[Lookup.scala 11:37:@6590.4]
  assign _T_601 = _T_52 ? 2'h0 : _T_600; // @[Lookup.scala 11:37:@6591.4]
  assign _T_602 = _T_48 ? 2'h0 : _T_601; // @[Lookup.scala 11:37:@6592.4]
  assign _T_603 = _T_44 ? 2'h0 : _T_602; // @[Lookup.scala 11:37:@6593.4]
  assign _T_604 = _T_40 ? 2'h0 : _T_603; // @[Lookup.scala 11:37:@6594.4]
  assign _T_605 = _T_36 ? 2'h1 : _T_604; // @[Lookup.scala 11:37:@6595.4]
  assign _T_606 = _T_32 ? 2'h1 : _T_605; // @[Lookup.scala 11:37:@6596.4]
  assign _T_607 = _T_28 ? 2'h1 : _T_606; // @[Lookup.scala 11:37:@6597.4]
  assign _T_608 = _T_24 ? 2'h1 : _T_607; // @[Lookup.scala 11:37:@6598.4]
  assign _T_622 = _T_164 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@6613.4]
  assign _T_623 = _T_160 ? 1'h0 : _T_622; // @[Lookup.scala 11:37:@6614.4]
  assign _T_624 = _T_156 ? 1'h0 : _T_623; // @[Lookup.scala 11:37:@6615.4]
  assign _T_625 = _T_152 ? 1'h0 : _T_624; // @[Lookup.scala 11:37:@6616.4]
  assign _T_626 = _T_148 ? 1'h0 : _T_625; // @[Lookup.scala 11:37:@6617.4]
  assign _T_627 = _T_144 ? 1'h0 : _T_626; // @[Lookup.scala 11:37:@6618.4]
  assign _T_628 = _T_140 ? 1'h1 : _T_627; // @[Lookup.scala 11:37:@6619.4]
  assign _T_629 = _T_136 ? 1'h1 : _T_628; // @[Lookup.scala 11:37:@6620.4]
  assign _T_630 = _T_132 ? 1'h1 : _T_629; // @[Lookup.scala 11:37:@6621.4]
  assign _T_631 = _T_128 ? 1'h1 : _T_630; // @[Lookup.scala 11:37:@6622.4]
  assign _T_632 = _T_124 ? 1'h1 : _T_631; // @[Lookup.scala 11:37:@6623.4]
  assign _T_633 = _T_120 ? 1'h1 : _T_632; // @[Lookup.scala 11:37:@6624.4]
  assign _T_634 = _T_116 ? 1'h1 : _T_633; // @[Lookup.scala 11:37:@6625.4]
  assign _T_635 = _T_112 ? 1'h1 : _T_634; // @[Lookup.scala 11:37:@6626.4]
  assign _T_636 = _T_108 ? 1'h1 : _T_635; // @[Lookup.scala 11:37:@6627.4]
  assign _T_637 = _T_104 ? 1'h1 : _T_636; // @[Lookup.scala 11:37:@6628.4]
  assign _T_638 = _T_100 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:@6629.4]
  assign _T_639 = _T_96 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:@6630.4]
  assign _T_640 = _T_92 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:@6631.4]
  assign _T_641 = _T_88 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:@6632.4]
  assign _T_642 = _T_84 ? 1'h1 : _T_641; // @[Lookup.scala 11:37:@6633.4]
  assign _T_643 = _T_80 ? 1'h1 : _T_642; // @[Lookup.scala 11:37:@6634.4]
  assign _T_644 = _T_76 ? 1'h1 : _T_643; // @[Lookup.scala 11:37:@6635.4]
  assign _T_645 = _T_72 ? 1'h1 : _T_644; // @[Lookup.scala 11:37:@6636.4]
  assign _T_646 = _T_68 ? 1'h1 : _T_645; // @[Lookup.scala 11:37:@6637.4]
  assign _T_647 = _T_64 ? 1'h1 : _T_646; // @[Lookup.scala 11:37:@6638.4]
  assign _T_648 = _T_60 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:@6639.4]
  assign _T_649 = _T_56 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:@6640.4]
  assign _T_650 = _T_52 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:@6641.4]
  assign _T_651 = _T_48 ? 1'h0 : _T_650; // @[Lookup.scala 11:37:@6642.4]
  assign _T_652 = _T_44 ? 1'h0 : _T_651; // @[Lookup.scala 11:37:@6643.4]
  assign _T_653 = _T_40 ? 1'h0 : _T_652; // @[Lookup.scala 11:37:@6644.4]
  assign _T_654 = _T_36 ? 1'h1 : _T_653; // @[Lookup.scala 11:37:@6645.4]
  assign _T_655 = _T_32 ? 1'h1 : _T_654; // @[Lookup.scala 11:37:@6646.4]
  assign _T_656 = _T_28 ? 1'h1 : _T_655; // @[Lookup.scala 11:37:@6647.4]
  assign _T_657 = _T_24 ? 1'h1 : _T_656; // @[Lookup.scala 11:37:@6648.4]
  assign _T_659 = _T_212 ? 1'h0 : _T_216; // @[Lookup.scala 11:37:@6651.4]
  assign _T_660 = _T_208 ? 1'h0 : _T_659; // @[Lookup.scala 11:37:@6652.4]
  assign _T_661 = _T_204 ? 1'h0 : _T_660; // @[Lookup.scala 11:37:@6653.4]
  assign _T_662 = _T_200 ? 1'h0 : _T_661; // @[Lookup.scala 11:37:@6654.4]
  assign _T_663 = _T_196 ? 1'h0 : _T_662; // @[Lookup.scala 11:37:@6655.4]
  assign _T_664 = _T_192 ? 1'h0 : _T_663; // @[Lookup.scala 11:37:@6656.4]
  assign _T_665 = _T_188 ? 1'h0 : _T_664; // @[Lookup.scala 11:37:@6657.4]
  assign _T_666 = _T_184 ? 1'h0 : _T_665; // @[Lookup.scala 11:37:@6658.4]
  assign _T_667 = _T_180 ? 1'h0 : _T_666; // @[Lookup.scala 11:37:@6659.4]
  assign _T_668 = _T_176 ? 1'h0 : _T_667; // @[Lookup.scala 11:37:@6660.4]
  assign _T_669 = _T_172 ? 1'h0 : _T_668; // @[Lookup.scala 11:37:@6661.4]
  assign _T_670 = _T_168 ? 1'h0 : _T_669; // @[Lookup.scala 11:37:@6662.4]
  assign _T_671 = _T_164 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:@6663.4]
  assign _T_672 = _T_160 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:@6664.4]
  assign _T_673 = _T_156 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:@6665.4]
  assign _T_674 = _T_152 ? 1'h0 : _T_673; // @[Lookup.scala 11:37:@6666.4]
  assign _T_675 = _T_148 ? 1'h0 : _T_674; // @[Lookup.scala 11:37:@6667.4]
  assign _T_676 = _T_144 ? 1'h0 : _T_675; // @[Lookup.scala 11:37:@6668.4]
  assign _T_677 = _T_140 ? 1'h0 : _T_676; // @[Lookup.scala 11:37:@6669.4]
  assign _T_678 = _T_136 ? 1'h0 : _T_677; // @[Lookup.scala 11:37:@6670.4]
  assign _T_679 = _T_132 ? 1'h0 : _T_678; // @[Lookup.scala 11:37:@6671.4]
  assign _T_680 = _T_128 ? 1'h0 : _T_679; // @[Lookup.scala 11:37:@6672.4]
  assign _T_681 = _T_124 ? 1'h0 : _T_680; // @[Lookup.scala 11:37:@6673.4]
  assign _T_682 = _T_120 ? 1'h0 : _T_681; // @[Lookup.scala 11:37:@6674.4]
  assign _T_683 = _T_116 ? 1'h0 : _T_682; // @[Lookup.scala 11:37:@6675.4]
  assign _T_684 = _T_112 ? 1'h0 : _T_683; // @[Lookup.scala 11:37:@6676.4]
  assign _T_685 = _T_108 ? 1'h0 : _T_684; // @[Lookup.scala 11:37:@6677.4]
  assign _T_686 = _T_104 ? 1'h0 : _T_685; // @[Lookup.scala 11:37:@6678.4]
  assign _T_687 = _T_100 ? 1'h0 : _T_686; // @[Lookup.scala 11:37:@6679.4]
  assign _T_688 = _T_96 ? 1'h0 : _T_687; // @[Lookup.scala 11:37:@6680.4]
  assign _T_689 = _T_92 ? 1'h0 : _T_688; // @[Lookup.scala 11:37:@6681.4]
  assign _T_690 = _T_88 ? 1'h0 : _T_689; // @[Lookup.scala 11:37:@6682.4]
  assign _T_691 = _T_84 ? 1'h0 : _T_690; // @[Lookup.scala 11:37:@6683.4]
  assign _T_692 = _T_80 ? 1'h0 : _T_691; // @[Lookup.scala 11:37:@6684.4]
  assign _T_693 = _T_76 ? 1'h0 : _T_692; // @[Lookup.scala 11:37:@6685.4]
  assign _T_694 = _T_72 ? 1'h0 : _T_693; // @[Lookup.scala 11:37:@6686.4]
  assign _T_695 = _T_68 ? 1'h0 : _T_694; // @[Lookup.scala 11:37:@6687.4]
  assign _T_696 = _T_64 ? 1'h0 : _T_695; // @[Lookup.scala 11:37:@6688.4]
  assign _T_697 = _T_60 ? 1'h0 : _T_696; // @[Lookup.scala 11:37:@6689.4]
  assign _T_698 = _T_56 ? 1'h0 : _T_697; // @[Lookup.scala 11:37:@6690.4]
  assign _T_699 = _T_52 ? 1'h0 : _T_698; // @[Lookup.scala 11:37:@6691.4]
  assign _T_700 = _T_48 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:@6692.4]
  assign _T_701 = _T_44 ? 1'h1 : _T_700; // @[Lookup.scala 11:37:@6693.4]
  assign _T_702 = _T_40 ? 1'h1 : _T_701; // @[Lookup.scala 11:37:@6694.4]
  assign _T_703 = _T_36 ? 1'h1 : _T_702; // @[Lookup.scala 11:37:@6695.4]
  assign _T_704 = _T_32 ? 1'h1 : _T_703; // @[Lookup.scala 11:37:@6696.4]
  assign _T_705 = _T_28 ? 1'h1 : _T_704; // @[Lookup.scala 11:37:@6697.4]
  assign _T_706 = _T_24 ? 1'h1 : _T_705; // @[Lookup.scala 11:37:@6698.4]
  assign _T_750 = _T_44 ? 1'h1 : _T_48; // @[Lookup.scala 11:37:@6743.4]
  assign _T_751 = _T_40 ? 1'h1 : _T_750; // @[Lookup.scala 11:37:@6744.4]
  assign _T_752 = _T_36 ? 1'h0 : _T_751; // @[Lookup.scala 11:37:@6745.4]
  assign _T_753 = _T_32 ? 1'h0 : _T_752; // @[Lookup.scala 11:37:@6746.4]
  assign _T_754 = _T_28 ? 1'h0 : _T_753; // @[Lookup.scala 11:37:@6747.4]
  assign _T_755 = _T_24 ? 1'h0 : _T_754; // @[Lookup.scala 11:37:@6748.4]
  assign _T_798 = _T_48 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@6792.4]
  assign _T_799 = _T_44 ? 3'h1 : _T_798; // @[Lookup.scala 11:37:@6793.4]
  assign _T_800 = _T_40 ? 3'h3 : _T_799; // @[Lookup.scala 11:37:@6794.4]
  assign _T_801 = _T_36 ? 3'h6 : _T_800; // @[Lookup.scala 11:37:@6795.4]
  assign _T_802 = _T_32 ? 3'h2 : _T_801; // @[Lookup.scala 11:37:@6796.4]
  assign _T_803 = _T_28 ? 3'h5 : _T_802; // @[Lookup.scala 11:37:@6797.4]
  assign _T_804 = _T_24 ? 3'h1 : _T_803; // @[Lookup.scala 11:37:@6798.4]
  assign _T_808 = _T_204 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@6803.4]
  assign _T_809 = _T_200 ? 3'h4 : _T_808; // @[Lookup.scala 11:37:@6804.4]
  assign _T_810 = _T_196 ? 3'h4 : _T_809; // @[Lookup.scala 11:37:@6805.4]
  assign _T_811 = _T_192 ? 3'h4 : _T_810; // @[Lookup.scala 11:37:@6806.4]
  assign _T_812 = _T_188 ? 3'h3 : _T_811; // @[Lookup.scala 11:37:@6807.4]
  assign _T_813 = _T_184 ? 3'h3 : _T_812; // @[Lookup.scala 11:37:@6808.4]
  assign _T_814 = _T_180 ? 3'h2 : _T_813; // @[Lookup.scala 11:37:@6809.4]
  assign _T_815 = _T_176 ? 3'h1 : _T_814; // @[Lookup.scala 11:37:@6810.4]
  assign _T_816 = _T_172 ? 3'h2 : _T_815; // @[Lookup.scala 11:37:@6811.4]
  assign _T_817 = _T_168 ? 3'h1 : _T_816; // @[Lookup.scala 11:37:@6812.4]
  assign _T_818 = _T_164 ? 3'h0 : _T_817; // @[Lookup.scala 11:37:@6813.4]
  assign _T_819 = _T_160 ? 3'h0 : _T_818; // @[Lookup.scala 11:37:@6814.4]
  assign _T_820 = _T_156 ? 3'h0 : _T_819; // @[Lookup.scala 11:37:@6815.4]
  assign _T_821 = _T_152 ? 3'h0 : _T_820; // @[Lookup.scala 11:37:@6816.4]
  assign _T_822 = _T_148 ? 3'h0 : _T_821; // @[Lookup.scala 11:37:@6817.4]
  assign _T_823 = _T_144 ? 3'h0 : _T_822; // @[Lookup.scala 11:37:@6818.4]
  assign _T_824 = _T_140 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@6819.4]
  assign _T_825 = _T_136 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@6820.4]
  assign _T_826 = _T_132 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@6821.4]
  assign _T_827 = _T_128 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@6822.4]
  assign _T_828 = _T_124 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@6823.4]
  assign _T_829 = _T_120 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@6824.4]
  assign _T_830 = _T_116 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@6825.4]
  assign _T_831 = _T_112 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@6826.4]
  assign _T_832 = _T_108 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@6827.4]
  assign _T_833 = _T_104 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@6828.4]
  assign _T_834 = _T_100 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@6829.4]
  assign _T_835 = _T_96 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@6830.4]
  assign _T_836 = _T_92 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@6831.4]
  assign _T_837 = _T_88 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@6832.4]
  assign _T_838 = _T_84 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@6833.4]
  assign _T_839 = _T_80 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@6834.4]
  assign _T_840 = _T_76 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@6835.4]
  assign _T_841 = _T_72 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@6836.4]
  assign _T_842 = _T_68 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@6837.4]
  assign _T_843 = _T_64 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@6838.4]
  assign _T_844 = _T_60 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@6839.4]
  assign _T_845 = _T_56 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@6840.4]
  assign _T_846 = _T_52 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@6841.4]
  assign _T_847 = _T_48 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@6842.4]
  assign _T_848 = _T_44 ? 3'h0 : _T_847; // @[Lookup.scala 11:37:@6843.4]
  assign _T_849 = _T_40 ? 3'h0 : _T_848; // @[Lookup.scala 11:37:@6844.4]
  assign _T_850 = _T_36 ? 3'h0 : _T_849; // @[Lookup.scala 11:37:@6845.4]
  assign _T_851 = _T_32 ? 3'h0 : _T_850; // @[Lookup.scala 11:37:@6846.4]
  assign _T_852 = _T_28 ? 3'h0 : _T_851; // @[Lookup.scala 11:37:@6847.4]
  assign _T_853 = _T_24 ? 3'h0 : _T_852; // @[Lookup.scala 11:37:@6848.4]
  assign _T_905 = io_inst[19:15]; // @[InstDecoder.scala 128:25:@6915.4]
  assign _T_907 = io_inst[11:7]; // @[InstDecoder.scala 130:25:@6919.4]
  assign imm_itype = io_inst[31:20]; // @[InstDecoder.scala 133:27:@6921.4]
  assign _T_908 = io_inst[31:25]; // @[InstDecoder.scala 134:31:@6922.4]
  assign imm_stype = {_T_908,_T_907}; // @[Cat.scala 30:58:@6924.4]
  assign _T_910 = io_inst[31]; // @[InstDecoder.scala 135:31:@6925.4]
  assign _T_911 = io_inst[7]; // @[InstDecoder.scala 135:44:@6926.4]
  assign _T_912 = io_inst[30:25]; // @[InstDecoder.scala 135:56:@6927.4]
  assign _T_913 = io_inst[11:8]; // @[InstDecoder.scala 135:73:@6928.4]
  assign imm_sbtype = {_T_910,_T_911,_T_912,_T_913}; // @[Cat.scala 30:58:@6931.4]
  assign imm_utype = io_inst[31:12]; // @[InstDecoder.scala 136:27:@6932.4]
  assign _T_917 = io_inst[19:12]; // @[InstDecoder.scala 137:44:@6934.4]
  assign _T_918 = io_inst[20]; // @[InstDecoder.scala 137:60:@6935.4]
  assign _T_919 = io_inst[30:21]; // @[InstDecoder.scala 137:73:@6936.4]
  assign imm_ujtype = {_T_910,_T_917,_T_918,_T_919}; // @[Cat.scala 30:58:@6939.4]
  assign _T_922 = imm_itype[11]; // @[InstDecoder.scala 140:43:@6940.4]
  assign _T_926 = _T_922 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@6942.4]
  assign _T_928 = imm_stype[11]; // @[InstDecoder.scala 141:43:@6945.4]
  assign _T_932 = _T_928 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@6947.4]
  assign _T_934 = imm_sbtype[11]; // @[InstDecoder.scala 142:44:@6950.4]
  assign _T_938 = _T_934 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@6952.4]
  assign _T_940 = {_T_938,_T_910,_T_911,_T_912,_T_913}; // @[Cat.scala 30:58:@6953.4]
  assign _T_948 = imm_ujtype[19]; // @[InstDecoder.scala 144:44:@6959.4]
  assign _T_952 = _T_948 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@6961.4]
  assign _T_954 = {_T_952,_T_910,_T_917,_T_918,_T_919}; // @[Cat.scala 30:58:@6962.4]
  assign io_cinfo_br_type = _T_20 ? 4'h0 : _T_314; // @[InstDecoder.scala 113:20:@6900.4]
  assign io_cinfo_op1_sel = _T_20 ? 2'h0 : _T_363; // @[InstDecoder.scala 114:20:@6901.4]
  assign io_cinfo_op2_sel = _T_20 ? 3'h1 : _T_412; // @[InstDecoder.scala 115:20:@6902.4]
  assign io_cinfo_rs1_oen = _T_20 ? 1'h1 : _T_461; // @[InstDecoder.scala 116:20:@6903.4]
  assign io_cinfo_rs2_oen = _T_20 ? 1'h0 : _T_510; // @[InstDecoder.scala 117:20:@6904.4]
  assign io_cinfo_alu_fun = _T_20 ? 4'h0 : _T_559; // @[InstDecoder.scala 118:20:@6905.4]
  assign io_cinfo_wb_sel = _T_20 ? 2'h1 : _T_608; // @[InstDecoder.scala 119:20:@6906.4]
  assign io_cinfo_rf_wen = _T_20 ? 1'h1 : _T_657; // @[InstDecoder.scala 120:20:@6907.4]
  assign io_cinfo_mem_en = _T_20 ? 1'h1 : _T_706; // @[InstDecoder.scala 121:20:@6908.4]
  assign io_cinfo_mem_fcn = _T_20 ? 1'h0 : _T_755; // @[InstDecoder.scala 122:20:@6909.4]
  assign io_cinfo_mem_typ = _T_20 ? 3'h3 : _T_804; // @[InstDecoder.scala 123:20:@6910.4]
  assign io_cinfo_csr_cmd = _T_20 ? 3'h0 : _T_853; // @[InstDecoder.scala 124:20:@6911.4]
  assign io_cinfo_illegal = signals_0 == 1'h0; // @[InstDecoder.scala 125:20:@6913.4]
  assign io_dinfo_imm_i = {_T_926,imm_itype}; // @[InstDecoder.scala 140:19:@6944.4]
  assign io_dinfo_imm_s = {_T_932,imm_stype}; // @[InstDecoder.scala 141:19:@6949.4]
  assign io_dinfo_imm_sb = {_T_940,1'h0}; // @[InstDecoder.scala 142:19:@6955.4]
  assign io_dinfo_imm_u = {imm_utype,12'h0}; // @[InstDecoder.scala 143:19:@6958.4]
  assign io_dinfo_imm_uj = {_T_954,1'h0}; // @[InstDecoder.scala 144:19:@6964.4]
  assign io_dinfo_imm_z = {27'h0,_T_905}; // @[InstDecoder.scala 145:19:@6968.4]
  assign io_rs1_addr = io_inst[19:15]; // @[InstDecoder.scala 128:15:@6916.4]
  assign io_rs2_addr = io_inst[24:20]; // @[InstDecoder.scala 129:15:@6918.4]
  assign io_wbaddr = io_inst[11:7]; // @[InstDecoder.scala 130:15:@6920.4]
endmodule
module BackEnd( // @[:@7845.2]
  input         clock, // @[:@7846.4]
  input         reset, // @[:@7847.4]
  output        io_mem_req_valid, // @[:@7848.4]
  output [31:0] io_mem_req_bits_addr, // @[:@7848.4]
  output [31:0] io_mem_req_bits_data, // @[:@7848.4]
  output        io_mem_req_bits_fcn, // @[:@7848.4]
  output [2:0]  io_mem_req_bits_typ, // @[:@7848.4]
  input         io_mem_resp_valid, // @[:@7848.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@7848.4]
  output [31:0] io_cyc, // @[:@7848.4]
  output        io_front_xcpt_valid, // @[:@7848.4]
  output [31:0] io_front_xcpt_bits, // @[:@7848.4]
  output        io_front_kill, // @[:@7848.4]
  output        io_front_forward_0, // @[:@7848.4]
  output        io_front_forward_1, // @[:@7848.4]
  input         io_front_inst_0_valid, // @[:@7848.4]
  input  [31:0] io_front_inst_0_bits, // @[:@7848.4]
  input         io_front_inst_1_valid, // @[:@7848.4]
  input  [31:0] io_front_inst_1_bits, // @[:@7848.4]
  input  [31:0] io_front_pc_0, // @[:@7848.4]
  input  [31:0] io_front_pc_1, // @[:@7848.4]
  input         io_front_split, // @[:@7848.4]
  input         io_front_pred_redirect, // @[:@7848.4]
  input  [9:0]  io_front_pred_history, // @[:@7848.4]
  input         io_front_pred_diff, // @[:@7848.4]
  input  [31:0] io_front_pred_tgt, // @[:@7848.4]
  input         io_front_branch, // @[:@7848.4]
  input         io_front_call, // @[:@7848.4]
  input         io_front_retn, // @[:@7848.4]
  input         io_front_bj_sel_0, // @[:@7848.4]
  input         io_front_bj_sel_1, // @[:@7848.4]
  output        io_front_ras_pop, // @[:@7848.4]
  output        io_front_ras_push_valid, // @[:@7848.4]
  output [31:0] io_front_ras_push_bits, // @[:@7848.4]
  output [31:0] io_front_fb_pc, // @[:@7848.4]
  output [1:0]  io_front_fb_type, // @[:@7848.4]
  output        io_front_feedBack_redirect, // @[:@7848.4]
  output [9:0]  io_front_feedBack_history, // @[:@7848.4]
  output        io_front_feedBack_diff, // @[:@7848.4]
  output [31:0] io_front_feedBack_tgt, // @[:@7848.4]
  output        io_front_feedBack_valid // @[:@7848.4]
);
  wire  csr_clock; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_reset; // @[BackEnd.scala 76:19:@7850.4]
  wire [2:0] csr_io_rw_cmd; // @[BackEnd.scala 76:19:@7850.4]
  wire [11:0] csr_io_rw_addr; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_rw_rdata; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_rw_wdata; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_eret; // @[BackEnd.scala 76:19:@7850.4]
  wire [1:0] csr_io_status_prv; // @[BackEnd.scala 76:19:@7850.4]
  wire [13:0] csr_io_status_unimp5; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_status_mprv; // @[BackEnd.scala 76:19:@7850.4]
  wire [1:0] csr_io_status_unimp4; // @[BackEnd.scala 76:19:@7850.4]
  wire [1:0] csr_io_status_mpp; // @[BackEnd.scala 76:19:@7850.4]
  wire [2:0] csr_io_status_unimp3; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_status_mpie; // @[BackEnd.scala 76:19:@7850.4]
  wire [2:0] csr_io_status_unimp2; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_status_mie; // @[BackEnd.scala 76:19:@7850.4]
  wire [2:0] csr_io_status_unimp1; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_xcpt; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_cause; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_tval; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_evec; // @[BackEnd.scala 76:19:@7850.4]
  wire  csr_io_illegal; // @[BackEnd.scala 76:19:@7850.4]
  wire [1:0] csr_io_retire; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_pc; // @[BackEnd.scala 76:19:@7850.4]
  wire [31:0] csr_io_time; // @[BackEnd.scala 76:19:@7850.4]
  wire  regfile_clock; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_rs1_addr_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_rs1_addr_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_rs1_data_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_rs1_data_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_rs2_addr_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_rs2_addr_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_rs2_data_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_rs2_data_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_waddr_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [4:0] regfile_io_waddr_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_wdata_0; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] regfile_io_wdata_1; // @[BackEnd.scala 77:23:@7853.4]
  wire  regfile_io_wen_0; // @[BackEnd.scala 77:23:@7853.4]
  wire  regfile_io_wen_1; // @[BackEnd.scala 77:23:@7853.4]
  wire [31:0] ALU_io_op1; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_op2; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_pc; // @[BackEnd.scala 78:33:@7856.4]
  wire [3:0] ALU_io_ctrl_fun; // @[BackEnd.scala 78:33:@7856.4]
  wire [3:0] ALU_io_ctrl_br_type; // @[BackEnd.scala 78:33:@7856.4]
  wire [1:0] ALU_io_ctrl_wb_sel; // @[BackEnd.scala 78:33:@7856.4]
  wire [1:0] ALU_io_ctrl_pc_sel; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_rs2_data; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_result; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_target_brjmp; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_target_jpreg; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_io_target_conti; // @[BackEnd.scala 78:33:@7856.4]
  wire [31:0] ALU_1_io_op1; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_op2; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_pc; // @[BackEnd.scala 78:33:@7859.4]
  wire [3:0] ALU_1_io_ctrl_fun; // @[BackEnd.scala 78:33:@7859.4]
  wire [3:0] ALU_1_io_ctrl_br_type; // @[BackEnd.scala 78:33:@7859.4]
  wire [1:0] ALU_1_io_ctrl_wb_sel; // @[BackEnd.scala 78:33:@7859.4]
  wire [1:0] ALU_1_io_ctrl_pc_sel; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_rs2_data; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_result; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_target_brjmp; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_target_jpreg; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] ALU_1_io_target_conti; // @[BackEnd.scala 78:33:@7859.4]
  wire [31:0] InstDecoder_io_inst; // @[BackEnd.scala 79:33:@7862.4]
  wire [3:0] InstDecoder_io_cinfo_br_type; // @[BackEnd.scala 79:33:@7862.4]
  wire [1:0] InstDecoder_io_cinfo_op1_sel; // @[BackEnd.scala 79:33:@7862.4]
  wire [2:0] InstDecoder_io_cinfo_op2_sel; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 79:33:@7862.4]
  wire [3:0] InstDecoder_io_cinfo_alu_fun; // @[BackEnd.scala 79:33:@7862.4]
  wire [1:0] InstDecoder_io_cinfo_wb_sel; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_mem_en; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_mem_fcn; // @[BackEnd.scala 79:33:@7862.4]
  wire [2:0] InstDecoder_io_cinfo_mem_typ; // @[BackEnd.scala 79:33:@7862.4]
  wire [2:0] InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 79:33:@7862.4]
  wire  InstDecoder_io_cinfo_illegal; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_i; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_s; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_sb; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_u; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_uj; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_io_dinfo_imm_z; // @[BackEnd.scala 79:33:@7862.4]
  wire [4:0] InstDecoder_io_rs1_addr; // @[BackEnd.scala 79:33:@7862.4]
  wire [4:0] InstDecoder_io_rs2_addr; // @[BackEnd.scala 79:33:@7862.4]
  wire [4:0] InstDecoder_io_wbaddr; // @[BackEnd.scala 79:33:@7862.4]
  wire [31:0] InstDecoder_1_io_inst; // @[BackEnd.scala 79:33:@7865.4]
  wire [3:0] InstDecoder_1_io_cinfo_br_type; // @[BackEnd.scala 79:33:@7865.4]
  wire [1:0] InstDecoder_1_io_cinfo_op1_sel; // @[BackEnd.scala 79:33:@7865.4]
  wire [2:0] InstDecoder_1_io_cinfo_op2_sel; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_rs1_oen; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_rs2_oen; // @[BackEnd.scala 79:33:@7865.4]
  wire [3:0] InstDecoder_1_io_cinfo_alu_fun; // @[BackEnd.scala 79:33:@7865.4]
  wire [1:0] InstDecoder_1_io_cinfo_wb_sel; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_rf_wen; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_mem_en; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_mem_fcn; // @[BackEnd.scala 79:33:@7865.4]
  wire [2:0] InstDecoder_1_io_cinfo_mem_typ; // @[BackEnd.scala 79:33:@7865.4]
  wire [2:0] InstDecoder_1_io_cinfo_csr_cmd; // @[BackEnd.scala 79:33:@7865.4]
  wire  InstDecoder_1_io_cinfo_illegal; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_i; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_s; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_sb; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_u; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_uj; // @[BackEnd.scala 79:33:@7865.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_z; // @[BackEnd.scala 79:33:@7865.4]
  wire [4:0] InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 79:33:@7865.4]
  wire [4:0] InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 79:33:@7865.4]
  wire [4:0] InstDecoder_1_io_wbaddr; // @[BackEnd.scala 79:33:@7865.4]
  reg  exe_0_rf_wen; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_0;
  reg [4:0] exe_0_wbaddr; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_1;
  reg  exe_0_mem_en; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_2;
  reg [2:0] exe_0_csr_cmd; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_3;
  reg  exe_0_illegal; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_4;
  reg [31:0] exe_0_pc; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_5;
  reg [31:0] exe_0_inst; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_6;
  reg [31:0] exe_0_rs2_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_7;
  reg [1:0] exe_0_wb_sel; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_8;
  reg  exe_0_mem_fcn; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_9;
  reg [2:0] exe_0_mem_typ; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_10;
  reg [3:0] exe_0_br_type; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_11;
  reg  exe_0_bj_sel; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_12;
  reg [31:0] exe_0_op1_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_13;
  reg [31:0] exe_0_op2_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_14;
  reg [3:0] exe_0_alu_fun; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_15;
  reg  exe_1_rf_wen; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_16;
  reg [4:0] exe_1_wbaddr; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_17;
  reg  exe_1_mem_en; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_18;
  reg [2:0] exe_1_csr_cmd; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_19;
  reg  exe_1_illegal; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_20;
  reg [31:0] exe_1_pc; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_21;
  reg [31:0] exe_1_inst; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_22;
  reg [31:0] exe_1_rs2_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_23;
  reg [1:0] exe_1_wb_sel; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_24;
  reg  exe_1_mem_fcn; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_25;
  reg [2:0] exe_1_mem_typ; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_26;
  reg [3:0] exe_1_br_type; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_27;
  reg  exe_1_bj_sel; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_28;
  reg [31:0] exe_1_op1_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_29;
  reg [31:0] exe_1_op2_data; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_30;
  reg [3:0] exe_1_alu_fun; // @[BackEnd.scala 86:22:@7873.4]
  reg [31:0] _RAND_31;
  reg  exe_valid_0; // @[BackEnd.scala 87:26:@7877.4]
  reg [31:0] _RAND_32;
  reg  exe_valid_1; // @[BackEnd.scala 87:26:@7877.4]
  reg [31:0] _RAND_33;
  reg  mem_0_rf_wen; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_34;
  reg [4:0] mem_0_wbaddr; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_35;
  reg  mem_0_mem_en; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_36;
  reg [2:0] mem_0_csr_cmd; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_37;
  reg  mem_0_illegal; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_38;
  reg [31:0] mem_0_pc; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_39;
  reg [31:0] mem_0_inst; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_40;
  reg [1:0] mem_0_wb_sel; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_41;
  reg  mem_0_mem_fcn; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_42;
  reg [2:0] mem_0_mem_typ; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_43;
  reg  mem_1_rf_wen; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_44;
  reg [4:0] mem_1_wbaddr; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_45;
  reg  mem_1_mem_en; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_46;
  reg [2:0] mem_1_csr_cmd; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_47;
  reg  mem_1_illegal; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_48;
  reg [31:0] mem_1_pc; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_49;
  reg [31:0] mem_1_inst; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_50;
  reg [1:0] mem_1_wb_sel; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_51;
  reg  mem_1_mem_fcn; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_52;
  reg [2:0] mem_1_mem_typ; // @[BackEnd.scala 89:22:@7879.4]
  reg [31:0] _RAND_53;
  reg  mem_valid_0; // @[BackEnd.scala 90:26:@7883.4]
  reg [31:0] _RAND_54;
  reg  mem_valid_1; // @[BackEnd.scala 90:26:@7883.4]
  reg [31:0] _RAND_55;
  reg  wb_0_rf_wen; // @[BackEnd.scala 92:22:@7885.4]
  reg [31:0] _RAND_56;
  reg [4:0] wb_0_wbaddr; // @[BackEnd.scala 92:22:@7885.4]
  reg [31:0] _RAND_57;
  reg  wb_1_rf_wen; // @[BackEnd.scala 92:22:@7885.4]
  reg [31:0] _RAND_58;
  reg [4:0] wb_1_wbaddr; // @[BackEnd.scala 92:22:@7885.4]
  reg [31:0] _RAND_59;
  reg  wb_valid_0; // @[BackEnd.scala 93:26:@7889.4]
  reg [31:0] _RAND_60;
  reg  wb_valid_1; // @[BackEnd.scala 93:26:@7889.4]
  reg [31:0] _RAND_61;
  reg [31:0] wb_wbdata_0; // @[BackEnd.scala 98:23:@7893.4]
  reg [31:0] _RAND_62;
  reg [31:0] wb_wbdata_1; // @[BackEnd.scala 98:23:@7893.4]
  reg [31:0] _RAND_63;
  wire  dec_wire_0_rs1_oen; // @[BackEnd.scala 111:51:@7901.4]
  wire  dec_wire_0_rs2_oen; // @[BackEnd.scala 112:51:@7903.4]
  wire  _T_542; // @[BackEnd.scala 113:51:@7905.4]
  wire  _T_544; // @[BackEnd.scala 113:91:@7906.4]
  wire  dec_wire_0_rf_wen; // @[BackEnd.scala 113:74:@7907.4]
  wire [2:0] dec_wire_0_csr_cmd; // @[BackEnd.scala 114:31:@7909.4]
  wire  _T_547; // @[BackEnd.scala 122:23:@7915.4]
  wire  _T_744; // @[BackEnd.scala 204:41:@8190.4]
  wire  _T_746; // @[BackEnd.scala 204:75:@8191.4]
  wire  exe_wire_1_rf_wen; // @[BackEnd.scala 204:58:@8192.4]
  wire  _T_548; // @[BackEnd.scala 122:44:@7916.4]
  wire  _T_549; // @[BackEnd.scala 123:23:@7917.4]
  wire  _T_733; // @[BackEnd.scala 204:41:@8153.4]
  wire  _T_735; // @[BackEnd.scala 204:75:@8154.4]
  wire  exe_wire_0_rf_wen; // @[BackEnd.scala 204:58:@8155.4]
  wire  _T_550; // @[BackEnd.scala 123:44:@7918.4]
  wire  _T_551; // @[BackEnd.scala 124:23:@7919.4]
  wire  _T_870; // @[BackEnd.scala 290:41:@8365.4]
  wire  _T_872; // @[BackEnd.scala 290:75:@8366.4]
  wire  mem_wire_1_rf_wen; // @[BackEnd.scala 290:58:@8367.4]
  wire  _T_552; // @[BackEnd.scala 124:44:@7920.4]
  wire  _T_553; // @[BackEnd.scala 125:23:@7921.4]
  wire  _T_851; // @[BackEnd.scala 290:41:@8337.4]
  wire  _T_853; // @[BackEnd.scala 290:75:@8338.4]
  wire  mem_wire_0_rf_wen; // @[BackEnd.scala 290:58:@8339.4]
  wire  _T_554; // @[BackEnd.scala 125:44:@7922.4]
  wire  _T_555; // @[BackEnd.scala 126:23:@7923.4]
  wire  _T_935; // @[BackEnd.scala 363:40:@8554.4]
  wire  _T_937; // @[BackEnd.scala 363:72:@8555.4]
  wire  wb_wire_1_rf_wen; // @[BackEnd.scala 363:56:@8556.4]
  wire  _T_556; // @[BackEnd.scala 126:44:@7924.4]
  wire  _T_557; // @[BackEnd.scala 127:23:@7925.4]
  wire  _T_931; // @[BackEnd.scala 363:40:@8547.4]
  wire  _T_933; // @[BackEnd.scala 363:72:@8548.4]
  wire  wb_wire_0_rf_wen; // @[BackEnd.scala 363:56:@8549.4]
  wire  _T_558; // @[BackEnd.scala 127:44:@7926.4]
  wire [31:0] rf_rs1_data_0; // @[BackEnd.scala 106:25:@7898.4 BackEnd.scala 118:20:@7913.4]
  wire [31:0] _T_559; // @[Mux.scala 61:16:@7927.4]
  wire [31:0] _T_560; // @[Mux.scala 61:16:@7928.4]
  wire  _T_866; // @[BackEnd.scala 302:22:@8356.4]
  wire  _T_867; // @[BackEnd.scala 303:22:@8357.4]
  reg [31:0] mem_reg_wbdata_0; // @[BackEnd.scala 202:28:@8152.4]
  reg [31:0] _RAND_64;
  wire [31:0] _T_868; // @[Mux.scala 61:16:@8358.4]
  wire [31:0] mem_wbdata_0; // @[Mux.scala 61:16:@8359.4]
  wire [31:0] _T_561; // @[Mux.scala 61:16:@7929.4]
  wire  _T_885; // @[BackEnd.scala 302:22:@8384.4]
  wire  _T_886; // @[BackEnd.scala 303:22:@8385.4]
  reg [31:0] mem_reg_wbdata_1; // @[BackEnd.scala 202:28:@8152.4]
  reg [31:0] _RAND_65;
  wire [31:0] _T_887; // @[Mux.scala 61:16:@8386.4]
  wire [31:0] mem_wbdata_1; // @[Mux.scala 61:16:@8387.4]
  wire [31:0] _T_562; // @[Mux.scala 61:16:@7930.4]
  wire [31:0] exe_wbdata_0; // @[BackEnd.scala 96:24:@7891.4 BackEnd.scala 219:19:@8174.4]
  wire [31:0] _T_563; // @[Mux.scala 61:16:@7931.4]
  wire [31:0] exe_wbdata_1; // @[BackEnd.scala 96:24:@7891.4 BackEnd.scala 219:19:@8211.4]
  wire [31:0] dec_rs1_data_0; // @[Mux.scala 61:16:@7932.4]
  wire  _T_565; // @[BackEnd.scala 131:23:@7934.4]
  wire  _T_566; // @[BackEnd.scala 131:44:@7935.4]
  wire  _T_567; // @[BackEnd.scala 132:23:@7936.4]
  wire  _T_568; // @[BackEnd.scala 132:44:@7937.4]
  wire  _T_569; // @[BackEnd.scala 133:23:@7938.4]
  wire  _T_570; // @[BackEnd.scala 133:44:@7939.4]
  wire  _T_571; // @[BackEnd.scala 134:23:@7940.4]
  wire  _T_572; // @[BackEnd.scala 134:44:@7941.4]
  wire  _T_573; // @[BackEnd.scala 135:23:@7942.4]
  wire  _T_574; // @[BackEnd.scala 135:44:@7943.4]
  wire  _T_575; // @[BackEnd.scala 136:23:@7944.4]
  wire  _T_576; // @[BackEnd.scala 136:44:@7945.4]
  wire [31:0] rf_rs2_data_0; // @[BackEnd.scala 107:25:@7899.4 BackEnd.scala 119:20:@7914.4]
  wire [31:0] _T_577; // @[Mux.scala 61:16:@7946.4]
  wire [31:0] _T_578; // @[Mux.scala 61:16:@7947.4]
  wire [31:0] _T_579; // @[Mux.scala 61:16:@7948.4]
  wire [31:0] _T_580; // @[Mux.scala 61:16:@7949.4]
  wire [31:0] _T_581; // @[Mux.scala 61:16:@7950.4]
  wire [31:0] dec_rs2_data_0; // @[Mux.scala 61:16:@7951.4]
  wire  _T_583; // @[BackEnd.scala 140:29:@7953.4]
  wire  _T_584; // @[BackEnd.scala 141:29:@7954.4]
  wire [31:0] _T_585; // @[Mux.scala 61:16:@7955.4]
  wire [31:0] dec_op1_data_0; // @[Mux.scala 61:16:@7956.4]
  wire  _T_587; // @[BackEnd.scala 144:29:@7958.4]
  wire  _T_588; // @[BackEnd.scala 145:29:@7959.4]
  wire  _T_589; // @[BackEnd.scala 146:29:@7960.4]
  wire  _T_590; // @[BackEnd.scala 147:29:@7961.4]
  wire  _T_591; // @[BackEnd.scala 148:29:@7962.4]
  wire [31:0] _T_592; // @[Mux.scala 61:16:@7963.4]
  wire [31:0] _T_593; // @[Mux.scala 61:16:@7964.4]
  wire [31:0] _T_594; // @[Mux.scala 61:16:@7965.4]
  wire [31:0] _T_595; // @[Mux.scala 61:16:@7966.4]
  wire [31:0] dec_op2_data_0; // @[Mux.scala 61:16:@7967.4]
  wire  exe_wire_0_mem_en; // @[BackEnd.scala 205:41:@8157.4]
  wire  exe_wire_1_mem_en; // @[BackEnd.scala 205:41:@8194.4]
  wire  stall_1_1; // @[BackEnd.scala 405:80:@8709.4]
  wire  _T_598; // @[BackEnd.scala 150:11:@7969.4]
  wire [2:0] mem_wire_1_csr_cmd; // @[BackEnd.scala 292:31:@8371.4]
  wire  _T_881; // @[BackEnd.scala 296:39:@8379.4]
  wire  mem_wire_1_mem_en; // @[BackEnd.scala 291:41:@8369.4]
  wire  _T_882; // @[BackEnd.scala 296:49:@8380.4]
  wire  mem_wire_1_illegal; // @[BackEnd.scala 293:41:@8373.4]
  wire  _T_883; // @[BackEnd.scala 297:39:@8381.4]
  reg [31:0] mem_reg_jpnpc; // @[BackEnd.scala 260:31:@8284.4]
  reg [31:0] _RAND_66;
  wire [1:0] _T_877; // @[BackEnd.scala 294:54:@8375.4]
  wire  _T_879; // @[BackEnd.scala 294:60:@8376.4]
  wire  mem_wire_jump_1; // @[BackEnd.scala 294:38:@8377.4]
  wire  mem_sel_1; // @[BackEnd.scala 298:39:@8382.4]
  wire [2:0] mem_wire_0_csr_cmd; // @[BackEnd.scala 292:31:@8343.4]
  wire  _T_862; // @[BackEnd.scala 296:39:@8351.4]
  wire  mem_wire_0_mem_en; // @[BackEnd.scala 291:41:@8341.4]
  wire  _T_863; // @[BackEnd.scala 296:49:@8352.4]
  wire  mem_wire_0_illegal; // @[BackEnd.scala 293:41:@8345.4]
  wire  _T_864; // @[BackEnd.scala 297:39:@8353.4]
  wire  mem_wire_jump_0; // @[BackEnd.scala 294:38:@8349.4]
  wire  mem_sel_0; // @[BackEnd.scala 298:39:@8354.4]
  wire [1:0] _T_1114; // @[BackEnd.scala 407:34:@8715.4]
  wire [1:0] _T_1115; // @[BackEnd.scala 407:41:@8716.4]
  wire  _T_1117; // @[BackEnd.scala 407:41:@8717.4]
  wire  _T_1119; // @[BackEnd.scala 407:72:@8718.4]
  wire  _T_1120; // @[BackEnd.scala 407:69:@8719.4]
  wire  _T_1121; // @[BackEnd.scala 407:46:@8720.4]
  wire  stall_0_2; // @[BackEnd.scala 406:45:@8713.4]
  wire  stall_1_2; // @[BackEnd.scala 407:92:@8721.4]
  wire  _T_600; // @[BackEnd.scala 150:35:@7970.4]
  wire  _T_601; // @[BackEnd.scala 150:32:@7971.4]
  wire  _T_602; // @[BackEnd.scala 154:52:@7975.6]
  wire  _T_603; // @[BackEnd.scala 154:86:@7976.6]
  wire  _T_604; // @[BackEnd.scala 154:62:@7977.6]
  wire  _T_606; // @[BackEnd.scala 155:47:@7978.6]
  wire  _T_607; // @[BackEnd.scala 154:97:@7979.6]
  wire [2:0] _T_608; // @[BackEnd.scala 154:29:@7980.6]
  wire  dec_wire_1_rs1_oen; // @[BackEnd.scala 111:51:@7997.4]
  wire  dec_wire_1_rs2_oen; // @[BackEnd.scala 112:51:@7999.4]
  wire  _T_616; // @[BackEnd.scala 122:23:@8011.4]
  wire  _T_617; // @[BackEnd.scala 122:44:@8012.4]
  wire  _T_618; // @[BackEnd.scala 123:23:@8013.4]
  wire  _T_619; // @[BackEnd.scala 123:44:@8014.4]
  wire  _T_620; // @[BackEnd.scala 124:23:@8015.4]
  wire  _T_621; // @[BackEnd.scala 124:44:@8016.4]
  wire  _T_622; // @[BackEnd.scala 125:23:@8017.4]
  wire  _T_623; // @[BackEnd.scala 125:44:@8018.4]
  wire  _T_624; // @[BackEnd.scala 126:23:@8019.4]
  wire  _T_625; // @[BackEnd.scala 126:44:@8020.4]
  wire  _T_626; // @[BackEnd.scala 127:23:@8021.4]
  wire  _T_627; // @[BackEnd.scala 127:44:@8022.4]
  wire [31:0] rf_rs1_data_1; // @[BackEnd.scala 106:25:@7898.4 BackEnd.scala 118:20:@8009.4]
  wire [31:0] _T_628; // @[Mux.scala 61:16:@8023.4]
  wire [31:0] _T_629; // @[Mux.scala 61:16:@8024.4]
  wire [31:0] _T_630; // @[Mux.scala 61:16:@8025.4]
  wire [31:0] _T_631; // @[Mux.scala 61:16:@8026.4]
  wire [31:0] _T_632; // @[Mux.scala 61:16:@8027.4]
  wire [31:0] dec_rs1_data_1; // @[Mux.scala 61:16:@8028.4]
  wire  _T_634; // @[BackEnd.scala 131:23:@8030.4]
  wire  _T_635; // @[BackEnd.scala 131:44:@8031.4]
  wire  _T_636; // @[BackEnd.scala 132:23:@8032.4]
  wire  _T_637; // @[BackEnd.scala 132:44:@8033.4]
  wire  _T_638; // @[BackEnd.scala 133:23:@8034.4]
  wire  _T_639; // @[BackEnd.scala 133:44:@8035.4]
  wire  _T_640; // @[BackEnd.scala 134:23:@8036.4]
  wire  _T_641; // @[BackEnd.scala 134:44:@8037.4]
  wire  _T_642; // @[BackEnd.scala 135:23:@8038.4]
  wire  _T_643; // @[BackEnd.scala 135:44:@8039.4]
  wire  _T_644; // @[BackEnd.scala 136:23:@8040.4]
  wire  _T_645; // @[BackEnd.scala 136:44:@8041.4]
  wire [31:0] rf_rs2_data_1; // @[BackEnd.scala 107:25:@7899.4 BackEnd.scala 119:20:@8010.4]
  wire [31:0] _T_646; // @[Mux.scala 61:16:@8042.4]
  wire [31:0] _T_647; // @[Mux.scala 61:16:@8043.4]
  wire [31:0] _T_648; // @[Mux.scala 61:16:@8044.4]
  wire [31:0] _T_649; // @[Mux.scala 61:16:@8045.4]
  wire [31:0] _T_650; // @[Mux.scala 61:16:@8046.4]
  wire [31:0] dec_rs2_data_1; // @[Mux.scala 61:16:@8047.4]
  wire  _T_652; // @[BackEnd.scala 140:29:@8049.4]
  wire  _T_653; // @[BackEnd.scala 141:29:@8050.4]
  wire [31:0] _T_654; // @[Mux.scala 61:16:@8051.4]
  wire [31:0] dec_op1_data_1; // @[Mux.scala 61:16:@8052.4]
  wire  _T_656; // @[BackEnd.scala 144:29:@8054.4]
  wire  _T_657; // @[BackEnd.scala 145:29:@8055.4]
  wire  _T_658; // @[BackEnd.scala 146:29:@8056.4]
  wire  _T_659; // @[BackEnd.scala 147:29:@8057.4]
  wire  _T_660; // @[BackEnd.scala 148:29:@8058.4]
  wire [31:0] _T_661; // @[Mux.scala 61:16:@8059.4]
  wire [31:0] _T_662; // @[Mux.scala 61:16:@8060.4]
  wire [31:0] _T_663; // @[Mux.scala 61:16:@8061.4]
  wire [31:0] _T_664; // @[Mux.scala 61:16:@8062.4]
  wire [31:0] dec_op2_data_1; // @[Mux.scala 61:16:@8063.4]
  wire  _T_671; // @[BackEnd.scala 154:52:@8071.6]
  wire  _T_672; // @[BackEnd.scala 154:86:@8072.6]
  wire  _T_673; // @[BackEnd.scala 154:62:@8073.6]
  wire  _T_675; // @[BackEnd.scala 155:47:@8074.6]
  wire  _T_676; // @[BackEnd.scala 154:97:@8075.6]
  wire [2:0] _T_677; // @[BackEnd.scala 154:29:@8076.6]
  reg  exe_btb_redirect; // @[BackEnd.scala 171:23:@8092.4]
  reg [31:0] _RAND_67;
  reg [9:0] exe_btb_history; // @[BackEnd.scala 171:23:@8092.4]
  reg [31:0] _RAND_68;
  reg  exe_btb_diff; // @[BackEnd.scala 171:23:@8092.4]
  reg [31:0] _RAND_69;
  reg [31:0] exe_btb_tgt; // @[BackEnd.scala 171:23:@8092.4]
  reg [31:0] _RAND_70;
  reg  exe_branch; // @[BackEnd.scala 172:23:@8093.4]
  reg [31:0] _RAND_71;
  reg  exe_call; // @[BackEnd.scala 173:23:@8094.4]
  reg [31:0] _RAND_72;
  reg  exe_retn; // @[BackEnd.scala 174:23:@8095.4]
  reg [31:0] _RAND_73;
  wire  rs1_addr_N0_0; // @[BackEnd.scala 388:41:@8638.4]
  wire  _T_1048; // @[BackEnd.scala 391:42:@8643.4]
  wire  _T_1049; // @[BackEnd.scala 391:60:@8644.4]
  wire  _T_1041; // @[BackEnd.scala 387:62:@8635.4]
  wire  exe_load_inst_0; // @[BackEnd.scala 387:44:@8636.4]
  wire  _T_1050; // @[BackEnd.scala 391:83:@8645.4]
  wire  rs2_addr_N0_0; // @[BackEnd.scala 389:41:@8640.4]
  wire  _T_1052; // @[BackEnd.scala 392:42:@8647.4]
  wire  _T_1053; // @[BackEnd.scala 392:60:@8648.4]
  wire  _T_1054; // @[BackEnd.scala 392:83:@8649.4]
  wire  _T_1055; // @[BackEnd.scala 391:104:@8650.4]
  wire  _T_1057; // @[BackEnd.scala 393:42:@8652.4]
  wire  _T_1058; // @[BackEnd.scala 393:60:@8653.4]
  wire  _T_1066; // @[BackEnd.scala 387:62:@8662.4]
  wire  exe_load_inst_1; // @[BackEnd.scala 387:44:@8663.4]
  wire  _T_1059; // @[BackEnd.scala 393:83:@8654.4]
  wire  _T_1060; // @[BackEnd.scala 392:104:@8655.4]
  wire  _T_1062; // @[BackEnd.scala 394:42:@8657.4]
  wire  _T_1063; // @[BackEnd.scala 394:60:@8658.4]
  wire  _T_1064; // @[BackEnd.scala 394:83:@8659.4]
  wire  rAW_0; // @[BackEnd.scala 393:104:@8660.4]
  wire [2:0] exe_wire_0_csr_cmd; // @[BackEnd.scala 206:31:@8159.4]
  wire  _T_1091; // @[BackEnd.scala 397:56:@8689.4]
  wire  _T_1092; // @[BackEnd.scala 397:33:@8690.4]
  wire [2:0] exe_wire_1_csr_cmd; // @[BackEnd.scala 206:31:@8196.4]
  wire  _T_1093; // @[BackEnd.scala 397:89:@8691.4]
  wire  stall_0_0; // @[BackEnd.scala 397:66:@8692.4]
  wire  _T_689; // @[BackEnd.scala 184:31:@8110.4]
  wire  _T_695; // @[BackEnd.scala 184:79:@8114.4]
  wire  ma_jump; // @[BackEnd.scala 334:29:@8510.4]
  wire  mem_en; // @[BackEnd.scala 316:25:@8398.4]
  wire  mem_fcn; // @[BackEnd.scala 317:25:@8399.4]
  wire  _T_901; // @[BackEnd.scala 332:44:@8504.4]
  wire  _T_902; // @[BackEnd.scala 332:33:@8505.4]
  wire [2:0] mem_typ; // @[BackEnd.scala 318:25:@8400.4]
  wire [1:0] _T_890; // @[BackEnd.scala 327:43:@8496.4]
  wire  _T_900; // @[Mux.scala 46:19:@8502.4]
  wire [31:0] mem_exe_out; // @[BackEnd.scala 312:25:@8394.4]
  wire  _T_893; // @[BackEnd.scala 328:23:@8497.4]
  wire  _T_898; // @[Mux.scala 46:19:@8500.4]
  wire [1:0] _T_895; // @[BackEnd.scala 329:23:@8498.4]
  wire  _T_897; // @[BackEnd.scala 329:29:@8499.4]
  wire  _T_899; // @[Mux.scala 46:16:@8501.4]
  wire  ls_addr_ma_valid; // @[Mux.scala 46:16:@8503.4]
  wire  ma_load; // @[BackEnd.scala 332:54:@8506.4]
  wire  _T_922; // @[BackEnd.scala 349:25:@8526.4]
  wire  _T_904; // @[BackEnd.scala 333:33:@8508.4]
  wire  ma_store; // @[BackEnd.scala 333:54:@8509.4]
  wire  _T_923; // @[BackEnd.scala 349:36:@8527.4]
  wire  ma_illegal; // @[BackEnd.scala 335:29:@8511.4]
  wire  _T_924; // @[BackEnd.scala 349:48:@8528.4]
  wire  xcpt_valid; // @[BackEnd.scala 349:62:@8529.4]
  wire  _T_696; // @[BackEnd.scala 184:104:@8115.4]
  wire  not_expect; // @[BackEnd.scala 256:48:@8279.4]
  wire  exe_wire_0_bj_sel; // @[BackEnd.scala 208:41:@8163.4]
  wire  exe_wire_1_bj_sel; // @[BackEnd.scala 208:41:@8200.4]
  wire  exe_bj_valid; // @[BackEnd.scala 198:56:@8148.4]
  wire  mispredict; // @[BackEnd.scala 257:28:@8280.4]
  wire  _T_704; // @[BackEnd.scala 187:47:@8124.8]
  wire  _T_705; // @[BackEnd.scala 187:44:@8125.8]
  wire  _GEN_39; // @[BackEnd.scala 186:60:@8123.6]
  wire  _GEN_40; // @[BackEnd.scala 184:119:@8116.4]
  wire  _T_1095; // @[BackEnd.scala 400:20:@8694.4]
  wire  rs1_addr_N0_1; // @[BackEnd.scala 388:41:@8665.4]
  wire  _T_1096; // @[BackEnd.scala 400:40:@8695.4]
  wire  _T_1097; // @[BackEnd.scala 400:58:@8696.4]
  wire  _T_1098; // @[BackEnd.scala 400:81:@8697.4]
  wire  _T_1099; // @[BackEnd.scala 401:20:@8698.4]
  wire  rs2_addr_N0_1; // @[BackEnd.scala 389:41:@8667.4]
  wire  _T_1100; // @[BackEnd.scala 401:40:@8699.4]
  wire  _T_1101; // @[BackEnd.scala 401:58:@8700.4]
  wire  _T_1102; // @[BackEnd.scala 401:81:@8701.4]
  wire  _T_1103; // @[BackEnd.scala 400:104:@8702.4]
  wire  _T_1104; // @[BackEnd.scala 402:25:@8703.4]
  wire  _T_1105; // @[BackEnd.scala 401:104:@8704.4]
  wire  _T_1073; // @[BackEnd.scala 391:42:@8670.4]
  wire  _T_1074; // @[BackEnd.scala 391:60:@8671.4]
  wire  _T_1075; // @[BackEnd.scala 391:83:@8672.4]
  wire  _T_1077; // @[BackEnd.scala 392:42:@8674.4]
  wire  _T_1078; // @[BackEnd.scala 392:60:@8675.4]
  wire  _T_1079; // @[BackEnd.scala 392:83:@8676.4]
  wire  _T_1080; // @[BackEnd.scala 391:104:@8677.4]
  wire  _T_1082; // @[BackEnd.scala 393:42:@8679.4]
  wire  _T_1083; // @[BackEnd.scala 393:60:@8680.4]
  wire  _T_1084; // @[BackEnd.scala 393:83:@8681.4]
  wire  _T_1085; // @[BackEnd.scala 392:104:@8682.4]
  wire  _T_1087; // @[BackEnd.scala 394:42:@8684.4]
  wire  _T_1088; // @[BackEnd.scala 394:60:@8685.4]
  wire  _T_1089; // @[BackEnd.scala 394:83:@8686.4]
  wire  rAW_1; // @[BackEnd.scala 393:104:@8687.4]
  wire  _T_1106; // @[BackEnd.scala 402:35:@8705.4]
  wire  stall_1_0; // @[BackEnd.scala 402:45:@8706.4]
  wire  _T_708; // @[BackEnd.scala 190:30:@8129.4]
  wire  _T_711; // @[BackEnd.scala 190:54:@8131.4]
  wire  _T_712; // @[BackEnd.scala 190:79:@8132.4]
  wire  exe_cancel; // @[BackEnd.scala 258:28:@8282.4]
  wire  _T_713; // @[BackEnd.scala 190:93:@8133.4]
  wire  _T_722; // @[BackEnd.scala 193:44:@8143.8]
  wire  _T_724; // @[BackEnd.scala 193:62:@8144.8]
  wire  _T_725; // @[BackEnd.scala 193:59:@8145.8]
  wire  _GEN_41; // @[BackEnd.scala 192:60:@8141.6]
  wire  _GEN_42; // @[BackEnd.scala 190:108:@8134.4]
  wire  exe_wire_branch; // @[BackEnd.scala 199:38:@8149.4]
  wire  exe_wire_call; // @[BackEnd.scala 200:38:@8150.4]
  wire  exe_wire_retn; // @[BackEnd.scala 201:38:@8151.4]
  wire [31:0] target_brjmp; // @[BackEnd.scala 237:19:@8227.4]
  wire [31:0] target_jpreg; // @[BackEnd.scala 237:19:@8227.4]
  wire [31:0] target_conti; // @[BackEnd.scala 237:19:@8227.4]
  wire [1:0] pc_sel; // @[BackEnd.scala 238:19:@8228.4]
  reg  _T_759; // @[BackEnd.scala 62:27:@8230.4]
  reg [31:0] _RAND_74;
  wire  _GEN_67; // @[BackEnd.scala 64:20:@8235.6]
  wire  _GEN_68; // @[BackEnd.scala 63:20:@8231.4]
  reg  _T_767; // @[BackEnd.scala 62:27:@8241.4]
  reg [31:0] _RAND_75;
  wire  _GEN_69; // @[BackEnd.scala 64:20:@8246.6]
  wire  _GEN_70; // @[BackEnd.scala 63:20:@8242.4]
  reg  _T_775; // @[BackEnd.scala 62:27:@8253.4]
  reg [31:0] _RAND_76;
  wire  _GEN_71; // @[BackEnd.scala 64:20:@8258.6]
  wire  _GEN_72; // @[BackEnd.scala 63:20:@8254.4]
  wire  _T_779; // @[BackEnd.scala 244:40:@8263.4]
  wire  _T_780; // @[BackEnd.scala 244:63:@8264.4]
  wire [31:0] _T_784; // @[BackEnd.scala 247:8:@8269.4]
  wire [1:0] _T_790; // @[BackEnd.scala 254:8:@8276.4]
  wire [31:0] _T_802; // @[Bitwise.scala 72:12:@8289.6]
  wire [31:0] _T_803; // @[BackEnd.scala 263:47:@8290.6]
  wire [31:0] _T_808; // @[Bitwise.scala 72:12:@8293.6]
  wire [31:0] _T_809; // @[BackEnd.scala 264:47:@8294.6]
  wire [31:0] _T_810; // @[BackEnd.scala 263:63:@8295.6]
  wire [31:0] _GEN_73; // @[BackEnd.scala 261:31:@8286.4]
  wire  _T_813; // @[BackEnd.scala 267:57:@8299.4]
  wire  _T_814; // @[BackEnd.scala 267:54:@8300.4]
  wire  _T_815; // @[BackEnd.scala 267:78:@8301.4]
  wire  _GEN_74; // @[BackEnd.scala 269:37:@8307.6]
  wire  _GEN_75; // @[BackEnd.scala 267:93:@8302.4]
  wire  _T_821; // @[BackEnd.scala 273:30:@8311.4]
  wire  _T_822; // @[BackEnd.scala 273:55:@8312.4]
  wire  _T_827; // @[BackEnd.scala 276:37:@8319.8]
  wire  _T_828; // @[BackEnd.scala 276:34:@8320.8]
  wire  _GEN_76; // @[BackEnd.scala 275:37:@8318.6]
  wire  _GEN_77; // @[BackEnd.scala 273:70:@8313.4]
  wire  _T_831; // @[BackEnd.scala 279:69:@8324.4]
  wire [31:0] mem_inst; // @[BackEnd.scala 311:25:@8393.4]
  wire  _T_905; // @[BackEnd.scala 336:27:@8512.4]
  wire  _T_906; // @[BackEnd.scala 336:39:@8513.4]
  wire [2:0] _T_913; // @[Mux.scala 61:16:@8516.4]
  wire [2:0] _T_914; // @[Mux.scala 61:16:@8517.4]
  wire [2:0] _T_915; // @[Mux.scala 61:16:@8518.4]
  wire [2:0] _T_916; // @[Mux.scala 61:16:@8519.4]
  wire [31:0] _T_918; // @[Mux.scala 61:16:@8521.4]
  wire [31:0] _T_919; // @[Mux.scala 61:16:@8522.4]
  wire [31:0] _T_920; // @[Mux.scala 61:16:@8523.4]
  wire  _T_926; // @[BackEnd.scala 352:44:@8532.4]
  wire  _T_927; // @[BackEnd.scala 352:29:@8533.4]
  wire  _GEN_78; // @[BackEnd.scala 352:60:@8534.4]
  wire  _T_929; // @[BackEnd.scala 356:29:@8540.4]
  wire  _GEN_79; // @[BackEnd.scala 356:44:@8541.4]
  wire [1:0] _T_946; // @[BackEnd.scala 375:25:@8562.4]
  wire  retire_0; // @[BackEnd.scala 375:32:@8563.4]
  wire [1:0] _T_949; // @[BackEnd.scala 376:32:@8566.4]
  wire  retire_1; // @[BackEnd.scala 376:32:@8567.4]
  reg  _T_1127; // @[BackEnd.scala 62:27:@8724.4]
  reg [31:0] _RAND_77;
  wire  _GEN_80; // @[BackEnd.scala 64:20:@8729.6]
  wire  _GEN_81; // @[BackEnd.scala 63:20:@8725.4]
  wire  _T_1132; // @[BackEnd.scala 411:26:@8736.4]
  wire  _T_1135; // @[BackEnd.scala 411:47:@8738.4]
  wire  _T_1140; // @[BackEnd.scala 412:26:@8742.4]
  wire  _T_1143; // @[BackEnd.scala 412:47:@8744.4]
  wire [7:0] _T_1149; // @[BackEnd.scala 421:12:@8748.4]
  wire [7:0] _T_1157; // @[BackEnd.scala 423:12:@8750.4]
  wire  _T_1160; // @[BackEnd.scala 424:32:@8751.4]
  wire  _T_1163; // @[BackEnd.scala 425:32:@8752.4]
  wire  _T_1166; // @[BackEnd.scala 426:32:@8753.4]
  wire  _T_1169; // @[BackEnd.scala 427:32:@8754.4]
  wire [7:0] _T_1172; // @[BackEnd.scala 427:12:@8755.4]
  wire [7:0] _T_1173; // @[BackEnd.scala 426:12:@8756.4]
  wire [7:0] _T_1174; // @[BackEnd.scala 425:12:@8757.4]
  wire [7:0] _T_1175; // @[BackEnd.scala 424:12:@8758.4]
  wire [7:0] _T_1179; // @[BackEnd.scala 428:12:@8759.4]
  wire  _T_1182; // @[BackEnd.scala 429:13:@8760.4]
  wire  _T_1183; // @[BackEnd.scala 429:27:@8761.4]
  wire  _T_1189; // @[BackEnd.scala 429:72:@8765.4]
  wire [31:0] _T_1195; // @[BackEnd.scala 429:12:@8769.4]
  wire  _T_1198; // @[BackEnd.scala 416:11:@8771.4]
  wire [7:0] _T_1201; // @[BackEnd.scala 421:12:@8775.4]
  wire [7:0] _T_1205; // @[BackEnd.scala 422:12:@8776.4]
  wire [7:0] _T_1209; // @[BackEnd.scala 423:12:@8777.4]
  wire  _T_1212; // @[BackEnd.scala 424:32:@8778.4]
  wire  _T_1215; // @[BackEnd.scala 425:32:@8779.4]
  wire  _T_1218; // @[BackEnd.scala 426:32:@8780.4]
  wire  _T_1221; // @[BackEnd.scala 427:32:@8781.4]
  wire [7:0] _T_1224; // @[BackEnd.scala 427:12:@8782.4]
  wire [7:0] _T_1225; // @[BackEnd.scala 426:12:@8783.4]
  wire [7:0] _T_1226; // @[BackEnd.scala 425:12:@8784.4]
  wire [7:0] _T_1227; // @[BackEnd.scala 424:12:@8785.4]
  wire  _T_1234; // @[BackEnd.scala 429:13:@8787.4]
  wire  _T_1235; // @[BackEnd.scala 429:27:@8788.4]
  wire  _T_1240; // @[BackEnd.scala 429:41:@8791.4]
  wire  _T_1241; // @[BackEnd.scala 429:72:@8792.4]
  wire  _T_1246; // @[BackEnd.scala 430:29:@8795.4]
  wire [31:0] _T_1247; // @[BackEnd.scala 429:12:@8796.4]
  wire [31:0] _T_1257; // @[BackEnd.scala 452:12:@8817.6]
  CSRFile csr ( // @[BackEnd.scala 76:19:@7850.4]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_status_prv(csr_io_status_prv),
    .io_status_unimp5(csr_io_status_unimp5),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_unimp4(csr_io_status_unimp4),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_unimp3(csr_io_status_unimp3),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_unimp2(csr_io_status_unimp2),
    .io_status_mie(csr_io_status_mie),
    .io_status_unimp1(csr_io_status_unimp1),
    .io_xcpt(csr_io_xcpt),
    .io_cause(csr_io_cause),
    .io_tval(csr_io_tval),
    .io_evec(csr_io_evec),
    .io_illegal(csr_io_illegal),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    .io_time(csr_io_time)
  );
  Regfile regfile ( // @[BackEnd.scala 77:23:@7853.4]
    .clock(regfile_clock),
    .io_rs1_addr_0(regfile_io_rs1_addr_0),
    .io_rs1_addr_1(regfile_io_rs1_addr_1),
    .io_rs1_data_0(regfile_io_rs1_data_0),
    .io_rs1_data_1(regfile_io_rs1_data_1),
    .io_rs2_addr_0(regfile_io_rs2_addr_0),
    .io_rs2_addr_1(regfile_io_rs2_addr_1),
    .io_rs2_data_0(regfile_io_rs2_data_0),
    .io_rs2_data_1(regfile_io_rs2_data_1),
    .io_waddr_0(regfile_io_waddr_0),
    .io_waddr_1(regfile_io_waddr_1),
    .io_wdata_0(regfile_io_wdata_0),
    .io_wdata_1(regfile_io_wdata_1),
    .io_wen_0(regfile_io_wen_0),
    .io_wen_1(regfile_io_wen_1)
  );
  ALU ALU ( // @[BackEnd.scala 78:33:@7856.4]
    .io_op1(ALU_io_op1),
    .io_op2(ALU_io_op2),
    .io_pc(ALU_io_pc),
    .io_ctrl_fun(ALU_io_ctrl_fun),
    .io_ctrl_br_type(ALU_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_io_ctrl_pc_sel),
    .io_rs2_data(ALU_io_rs2_data),
    .io_result(ALU_io_result),
    .io_target_brjmp(ALU_io_target_brjmp),
    .io_target_jpreg(ALU_io_target_jpreg),
    .io_target_conti(ALU_io_target_conti)
  );
  ALU ALU_1 ( // @[BackEnd.scala 78:33:@7859.4]
    .io_op1(ALU_1_io_op1),
    .io_op2(ALU_1_io_op2),
    .io_pc(ALU_1_io_pc),
    .io_ctrl_fun(ALU_1_io_ctrl_fun),
    .io_ctrl_br_type(ALU_1_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_1_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_1_io_ctrl_pc_sel),
    .io_rs2_data(ALU_1_io_rs2_data),
    .io_result(ALU_1_io_result),
    .io_target_brjmp(ALU_1_io_target_brjmp),
    .io_target_jpreg(ALU_1_io_target_jpreg),
    .io_target_conti(ALU_1_io_target_conti)
  );
  InstDecoder InstDecoder ( // @[BackEnd.scala 79:33:@7862.4]
    .io_inst(InstDecoder_io_inst),
    .io_cinfo_br_type(InstDecoder_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_io_cinfo_illegal),
    .io_dinfo_imm_i(InstDecoder_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_io_dinfo_imm_z),
    .io_rs1_addr(InstDecoder_io_rs1_addr),
    .io_rs2_addr(InstDecoder_io_rs2_addr),
    .io_wbaddr(InstDecoder_io_wbaddr)
  );
  InstDecoder InstDecoder_1 ( // @[BackEnd.scala 79:33:@7865.4]
    .io_inst(InstDecoder_1_io_inst),
    .io_cinfo_br_type(InstDecoder_1_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_1_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_1_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_1_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_1_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_1_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_1_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_1_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_1_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_1_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_1_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_1_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_1_io_cinfo_illegal),
    .io_dinfo_imm_i(InstDecoder_1_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_1_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_1_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_1_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_1_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_1_io_dinfo_imm_z),
    .io_rs1_addr(InstDecoder_1_io_rs1_addr),
    .io_rs2_addr(InstDecoder_1_io_rs2_addr),
    .io_wbaddr(InstDecoder_1_io_wbaddr)
  );
  assign dec_wire_0_rs1_oen = io_front_inst_0_valid & InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 111:51:@7901.4]
  assign dec_wire_0_rs2_oen = io_front_inst_0_valid & InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 112:51:@7903.4]
  assign _T_542 = io_front_inst_0_valid & InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 113:51:@7905.4]
  assign _T_544 = InstDecoder_io_wbaddr != 5'h0; // @[BackEnd.scala 113:91:@7906.4]
  assign dec_wire_0_rf_wen = _T_542 & _T_544; // @[BackEnd.scala 113:74:@7907.4]
  assign dec_wire_0_csr_cmd = io_front_inst_0_valid ? InstDecoder_io_cinfo_csr_cmd : 3'h0; // @[BackEnd.scala 114:31:@7909.4]
  assign _T_547 = exe_1_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 122:23:@7915.4]
  assign _T_744 = exe_valid_1 & exe_1_rf_wen; // @[BackEnd.scala 204:41:@8190.4]
  assign _T_746 = exe_1_wbaddr != 5'h0; // @[BackEnd.scala 204:75:@8191.4]
  assign exe_wire_1_rf_wen = _T_744 & _T_746; // @[BackEnd.scala 204:58:@8192.4]
  assign _T_548 = _T_547 & exe_wire_1_rf_wen; // @[BackEnd.scala 122:44:@7916.4]
  assign _T_549 = exe_0_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 123:23:@7917.4]
  assign _T_733 = exe_valid_0 & exe_0_rf_wen; // @[BackEnd.scala 204:41:@8153.4]
  assign _T_735 = exe_0_wbaddr != 5'h0; // @[BackEnd.scala 204:75:@8154.4]
  assign exe_wire_0_rf_wen = _T_733 & _T_735; // @[BackEnd.scala 204:58:@8155.4]
  assign _T_550 = _T_549 & exe_wire_0_rf_wen; // @[BackEnd.scala 123:44:@7918.4]
  assign _T_551 = mem_1_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 124:23:@7919.4]
  assign _T_870 = mem_valid_1 & mem_1_rf_wen; // @[BackEnd.scala 290:41:@8365.4]
  assign _T_872 = mem_1_wbaddr != 5'h0; // @[BackEnd.scala 290:75:@8366.4]
  assign mem_wire_1_rf_wen = _T_870 & _T_872; // @[BackEnd.scala 290:58:@8367.4]
  assign _T_552 = _T_551 & mem_wire_1_rf_wen; // @[BackEnd.scala 124:44:@7920.4]
  assign _T_553 = mem_0_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 125:23:@7921.4]
  assign _T_851 = mem_valid_0 & mem_0_rf_wen; // @[BackEnd.scala 290:41:@8337.4]
  assign _T_853 = mem_0_wbaddr != 5'h0; // @[BackEnd.scala 290:75:@8338.4]
  assign mem_wire_0_rf_wen = _T_851 & _T_853; // @[BackEnd.scala 290:58:@8339.4]
  assign _T_554 = _T_553 & mem_wire_0_rf_wen; // @[BackEnd.scala 125:44:@7922.4]
  assign _T_555 = wb_1_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 126:23:@7923.4]
  assign _T_935 = wb_valid_1 & wb_1_rf_wen; // @[BackEnd.scala 363:40:@8554.4]
  assign _T_937 = wb_1_wbaddr != 5'h0; // @[BackEnd.scala 363:72:@8555.4]
  assign wb_wire_1_rf_wen = _T_935 & _T_937; // @[BackEnd.scala 363:56:@8556.4]
  assign _T_556 = _T_555 & wb_wire_1_rf_wen; // @[BackEnd.scala 126:44:@7924.4]
  assign _T_557 = wb_0_wbaddr == InstDecoder_io_rs1_addr; // @[BackEnd.scala 127:23:@7925.4]
  assign _T_931 = wb_valid_0 & wb_0_rf_wen; // @[BackEnd.scala 363:40:@8547.4]
  assign _T_933 = wb_0_wbaddr != 5'h0; // @[BackEnd.scala 363:72:@8548.4]
  assign wb_wire_0_rf_wen = _T_931 & _T_933; // @[BackEnd.scala 363:56:@8549.4]
  assign _T_558 = _T_557 & wb_wire_0_rf_wen; // @[BackEnd.scala 127:44:@7926.4]
  assign rf_rs1_data_0 = regfile_io_rs1_data_0; // @[BackEnd.scala 106:25:@7898.4 BackEnd.scala 118:20:@7913.4]
  assign _T_559 = _T_558 ? wb_wbdata_0 : rf_rs1_data_0; // @[Mux.scala 61:16:@7927.4]
  assign _T_560 = _T_556 ? wb_wbdata_1 : _T_559; // @[Mux.scala 61:16:@7928.4]
  assign _T_866 = mem_0_wb_sel == 2'h1; // @[BackEnd.scala 302:22:@8356.4]
  assign _T_867 = mem_0_wb_sel == 2'h3; // @[BackEnd.scala 303:22:@8357.4]
  assign _T_868 = _T_867 ? csr_io_rw_rdata : mem_reg_wbdata_0; // @[Mux.scala 61:16:@8358.4]
  assign mem_wbdata_0 = _T_866 ? io_mem_resp_bits_data : _T_868; // @[Mux.scala 61:16:@8359.4]
  assign _T_561 = _T_554 ? mem_wbdata_0 : _T_560; // @[Mux.scala 61:16:@7929.4]
  assign _T_885 = mem_1_wb_sel == 2'h1; // @[BackEnd.scala 302:22:@8384.4]
  assign _T_886 = mem_1_wb_sel == 2'h3; // @[BackEnd.scala 303:22:@8385.4]
  assign _T_887 = _T_886 ? csr_io_rw_rdata : mem_reg_wbdata_1; // @[Mux.scala 61:16:@8386.4]
  assign mem_wbdata_1 = _T_885 ? io_mem_resp_bits_data : _T_887; // @[Mux.scala 61:16:@8387.4]
  assign _T_562 = _T_552 ? mem_wbdata_1 : _T_561; // @[Mux.scala 61:16:@7930.4]
  assign exe_wbdata_0 = ALU_io_result; // @[BackEnd.scala 96:24:@7891.4 BackEnd.scala 219:19:@8174.4]
  assign _T_563 = _T_550 ? exe_wbdata_0 : _T_562; // @[Mux.scala 61:16:@7931.4]
  assign exe_wbdata_1 = ALU_1_io_result; // @[BackEnd.scala 96:24:@7891.4 BackEnd.scala 219:19:@8211.4]
  assign dec_rs1_data_0 = _T_548 ? exe_wbdata_1 : _T_563; // @[Mux.scala 61:16:@7932.4]
  assign _T_565 = exe_1_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 131:23:@7934.4]
  assign _T_566 = _T_565 & exe_wire_1_rf_wen; // @[BackEnd.scala 131:44:@7935.4]
  assign _T_567 = exe_0_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 132:23:@7936.4]
  assign _T_568 = _T_567 & exe_wire_0_rf_wen; // @[BackEnd.scala 132:44:@7937.4]
  assign _T_569 = mem_1_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 133:23:@7938.4]
  assign _T_570 = _T_569 & mem_wire_1_rf_wen; // @[BackEnd.scala 133:44:@7939.4]
  assign _T_571 = mem_0_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 134:23:@7940.4]
  assign _T_572 = _T_571 & mem_wire_0_rf_wen; // @[BackEnd.scala 134:44:@7941.4]
  assign _T_573 = wb_1_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 135:23:@7942.4]
  assign _T_574 = _T_573 & wb_wire_1_rf_wen; // @[BackEnd.scala 135:44:@7943.4]
  assign _T_575 = wb_0_wbaddr == InstDecoder_io_rs2_addr; // @[BackEnd.scala 136:23:@7944.4]
  assign _T_576 = _T_575 & wb_wire_0_rf_wen; // @[BackEnd.scala 136:44:@7945.4]
  assign rf_rs2_data_0 = regfile_io_rs2_data_0; // @[BackEnd.scala 107:25:@7899.4 BackEnd.scala 119:20:@7914.4]
  assign _T_577 = _T_576 ? wb_wbdata_0 : rf_rs2_data_0; // @[Mux.scala 61:16:@7946.4]
  assign _T_578 = _T_574 ? wb_wbdata_1 : _T_577; // @[Mux.scala 61:16:@7947.4]
  assign _T_579 = _T_572 ? mem_wbdata_0 : _T_578; // @[Mux.scala 61:16:@7948.4]
  assign _T_580 = _T_570 ? mem_wbdata_1 : _T_579; // @[Mux.scala 61:16:@7949.4]
  assign _T_581 = _T_568 ? exe_wbdata_0 : _T_580; // @[Mux.scala 61:16:@7950.4]
  assign dec_rs2_data_0 = _T_566 ? exe_wbdata_1 : _T_581; // @[Mux.scala 61:16:@7951.4]
  assign _T_583 = InstDecoder_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 140:29:@7953.4]
  assign _T_584 = InstDecoder_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 141:29:@7954.4]
  assign _T_585 = _T_584 ? io_front_pc_0 : dec_rs1_data_0; // @[Mux.scala 61:16:@7955.4]
  assign dec_op1_data_0 = _T_583 ? InstDecoder_io_dinfo_imm_z : _T_585; // @[Mux.scala 61:16:@7956.4]
  assign _T_587 = InstDecoder_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 144:29:@7958.4]
  assign _T_588 = InstDecoder_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 145:29:@7959.4]
  assign _T_589 = InstDecoder_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 146:29:@7960.4]
  assign _T_590 = InstDecoder_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 147:29:@7961.4]
  assign _T_591 = InstDecoder_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 148:29:@7962.4]
  assign _T_592 = _T_591 ? InstDecoder_io_dinfo_imm_uj : dec_rs2_data_0; // @[Mux.scala 61:16:@7963.4]
  assign _T_593 = _T_590 ? InstDecoder_io_dinfo_imm_u : _T_592; // @[Mux.scala 61:16:@7964.4]
  assign _T_594 = _T_589 ? InstDecoder_io_dinfo_imm_sb : _T_593; // @[Mux.scala 61:16:@7965.4]
  assign _T_595 = _T_588 ? InstDecoder_io_dinfo_imm_s : _T_594; // @[Mux.scala 61:16:@7966.4]
  assign dec_op2_data_0 = _T_587 ? InstDecoder_io_dinfo_imm_i : _T_595; // @[Mux.scala 61:16:@7967.4]
  assign exe_wire_0_mem_en = exe_valid_0 & exe_0_mem_en; // @[BackEnd.scala 205:41:@8157.4]
  assign exe_wire_1_mem_en = exe_valid_1 & exe_1_mem_en; // @[BackEnd.scala 205:41:@8194.4]
  assign stall_1_1 = exe_wire_0_mem_en & exe_wire_1_mem_en; // @[BackEnd.scala 405:80:@8709.4]
  assign _T_598 = stall_1_1 == 1'h0; // @[BackEnd.scala 150:11:@7969.4]
  assign mem_wire_1_csr_cmd = mem_valid_1 ? mem_1_csr_cmd : 3'h0; // @[BackEnd.scala 292:31:@8371.4]
  assign _T_881 = mem_wire_1_csr_cmd != 3'h0; // @[BackEnd.scala 296:39:@8379.4]
  assign mem_wire_1_mem_en = mem_valid_1 & mem_1_mem_en; // @[BackEnd.scala 291:41:@8369.4]
  assign _T_882 = _T_881 | mem_wire_1_mem_en; // @[BackEnd.scala 296:49:@8380.4]
  assign mem_wire_1_illegal = mem_valid_1 & mem_1_illegal; // @[BackEnd.scala 293:41:@8373.4]
  assign _T_883 = _T_882 | mem_wire_1_illegal; // @[BackEnd.scala 297:39:@8381.4]
  assign _T_877 = mem_reg_jpnpc[1:0]; // @[BackEnd.scala 294:54:@8375.4]
  assign _T_879 = _T_877 != 2'h0; // @[BackEnd.scala 294:60:@8376.4]
  assign mem_wire_jump_1 = mem_valid_1 & _T_879; // @[BackEnd.scala 294:38:@8377.4]
  assign mem_sel_1 = _T_883 | mem_wire_jump_1; // @[BackEnd.scala 298:39:@8382.4]
  assign mem_wire_0_csr_cmd = mem_valid_0 ? mem_0_csr_cmd : 3'h0; // @[BackEnd.scala 292:31:@8343.4]
  assign _T_862 = mem_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 296:39:@8351.4]
  assign mem_wire_0_mem_en = mem_valid_0 & mem_0_mem_en; // @[BackEnd.scala 291:41:@8341.4]
  assign _T_863 = _T_862 | mem_wire_0_mem_en; // @[BackEnd.scala 296:49:@8352.4]
  assign mem_wire_0_illegal = mem_valid_0 & mem_0_illegal; // @[BackEnd.scala 293:41:@8345.4]
  assign _T_864 = _T_863 | mem_wire_0_illegal; // @[BackEnd.scala 297:39:@8353.4]
  assign mem_wire_jump_0 = mem_valid_0 & _T_879; // @[BackEnd.scala 294:38:@8349.4]
  assign mem_sel_0 = _T_864 | mem_wire_jump_0; // @[BackEnd.scala 298:39:@8354.4]
  assign _T_1114 = {mem_sel_1,mem_sel_0}; // @[BackEnd.scala 407:34:@8715.4]
  assign _T_1115 = ~ _T_1114; // @[BackEnd.scala 407:41:@8716.4]
  assign _T_1117 = _T_1115 == 2'h0; // @[BackEnd.scala 407:41:@8717.4]
  assign _T_1119 = io_mem_resp_valid == 1'h0; // @[BackEnd.scala 407:72:@8718.4]
  assign _T_1120 = mem_wire_1_mem_en & _T_1119; // @[BackEnd.scala 407:69:@8719.4]
  assign _T_1121 = _T_1117 | _T_1120; // @[BackEnd.scala 407:46:@8720.4]
  assign stall_0_2 = mem_wire_0_mem_en & _T_1119; // @[BackEnd.scala 406:45:@8713.4]
  assign stall_1_2 = _T_1121 | stall_0_2; // @[BackEnd.scala 407:92:@8721.4]
  assign _T_600 = stall_1_2 == 1'h0; // @[BackEnd.scala 150:35:@7970.4]
  assign _T_601 = _T_598 & _T_600; // @[BackEnd.scala 150:32:@7971.4]
  assign _T_602 = InstDecoder_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 154:52:@7975.6]
  assign _T_603 = InstDecoder_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 154:86:@7976.6]
  assign _T_604 = _T_602 | _T_603; // @[BackEnd.scala 154:62:@7977.6]
  assign _T_606 = InstDecoder_io_rs1_addr == 5'h0; // @[BackEnd.scala 155:47:@7978.6]
  assign _T_607 = _T_604 & _T_606; // @[BackEnd.scala 154:97:@7979.6]
  assign _T_608 = _T_607 ? 3'h5 : InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 154:29:@7980.6]
  assign dec_wire_1_rs1_oen = io_front_inst_1_valid & InstDecoder_1_io_cinfo_rs1_oen; // @[BackEnd.scala 111:51:@7997.4]
  assign dec_wire_1_rs2_oen = io_front_inst_1_valid & InstDecoder_1_io_cinfo_rs2_oen; // @[BackEnd.scala 112:51:@7999.4]
  assign _T_616 = exe_1_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 122:23:@8011.4]
  assign _T_617 = _T_616 & exe_wire_1_rf_wen; // @[BackEnd.scala 122:44:@8012.4]
  assign _T_618 = exe_0_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 123:23:@8013.4]
  assign _T_619 = _T_618 & exe_wire_0_rf_wen; // @[BackEnd.scala 123:44:@8014.4]
  assign _T_620 = mem_1_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 124:23:@8015.4]
  assign _T_621 = _T_620 & mem_wire_1_rf_wen; // @[BackEnd.scala 124:44:@8016.4]
  assign _T_622 = mem_0_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 125:23:@8017.4]
  assign _T_623 = _T_622 & mem_wire_0_rf_wen; // @[BackEnd.scala 125:44:@8018.4]
  assign _T_624 = wb_1_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 126:23:@8019.4]
  assign _T_625 = _T_624 & wb_wire_1_rf_wen; // @[BackEnd.scala 126:44:@8020.4]
  assign _T_626 = wb_0_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 127:23:@8021.4]
  assign _T_627 = _T_626 & wb_wire_0_rf_wen; // @[BackEnd.scala 127:44:@8022.4]
  assign rf_rs1_data_1 = regfile_io_rs1_data_1; // @[BackEnd.scala 106:25:@7898.4 BackEnd.scala 118:20:@8009.4]
  assign _T_628 = _T_627 ? wb_wbdata_0 : rf_rs1_data_1; // @[Mux.scala 61:16:@8023.4]
  assign _T_629 = _T_625 ? wb_wbdata_1 : _T_628; // @[Mux.scala 61:16:@8024.4]
  assign _T_630 = _T_623 ? mem_wbdata_0 : _T_629; // @[Mux.scala 61:16:@8025.4]
  assign _T_631 = _T_621 ? mem_wbdata_1 : _T_630; // @[Mux.scala 61:16:@8026.4]
  assign _T_632 = _T_619 ? exe_wbdata_0 : _T_631; // @[Mux.scala 61:16:@8027.4]
  assign dec_rs1_data_1 = _T_617 ? exe_wbdata_1 : _T_632; // @[Mux.scala 61:16:@8028.4]
  assign _T_634 = exe_1_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 131:23:@8030.4]
  assign _T_635 = _T_634 & exe_wire_1_rf_wen; // @[BackEnd.scala 131:44:@8031.4]
  assign _T_636 = exe_0_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 132:23:@8032.4]
  assign _T_637 = _T_636 & exe_wire_0_rf_wen; // @[BackEnd.scala 132:44:@8033.4]
  assign _T_638 = mem_1_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 133:23:@8034.4]
  assign _T_639 = _T_638 & mem_wire_1_rf_wen; // @[BackEnd.scala 133:44:@8035.4]
  assign _T_640 = mem_0_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 134:23:@8036.4]
  assign _T_641 = _T_640 & mem_wire_0_rf_wen; // @[BackEnd.scala 134:44:@8037.4]
  assign _T_642 = wb_1_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 135:23:@8038.4]
  assign _T_643 = _T_642 & wb_wire_1_rf_wen; // @[BackEnd.scala 135:44:@8039.4]
  assign _T_644 = wb_0_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 136:23:@8040.4]
  assign _T_645 = _T_644 & wb_wire_0_rf_wen; // @[BackEnd.scala 136:44:@8041.4]
  assign rf_rs2_data_1 = regfile_io_rs2_data_1; // @[BackEnd.scala 107:25:@7899.4 BackEnd.scala 119:20:@8010.4]
  assign _T_646 = _T_645 ? wb_wbdata_0 : rf_rs2_data_1; // @[Mux.scala 61:16:@8042.4]
  assign _T_647 = _T_643 ? wb_wbdata_1 : _T_646; // @[Mux.scala 61:16:@8043.4]
  assign _T_648 = _T_641 ? mem_wbdata_0 : _T_647; // @[Mux.scala 61:16:@8044.4]
  assign _T_649 = _T_639 ? mem_wbdata_1 : _T_648; // @[Mux.scala 61:16:@8045.4]
  assign _T_650 = _T_637 ? exe_wbdata_0 : _T_649; // @[Mux.scala 61:16:@8046.4]
  assign dec_rs2_data_1 = _T_635 ? exe_wbdata_1 : _T_650; // @[Mux.scala 61:16:@8047.4]
  assign _T_652 = InstDecoder_1_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 140:29:@8049.4]
  assign _T_653 = InstDecoder_1_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 141:29:@8050.4]
  assign _T_654 = _T_653 ? io_front_pc_1 : dec_rs1_data_1; // @[Mux.scala 61:16:@8051.4]
  assign dec_op1_data_1 = _T_652 ? InstDecoder_1_io_dinfo_imm_z : _T_654; // @[Mux.scala 61:16:@8052.4]
  assign _T_656 = InstDecoder_1_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 144:29:@8054.4]
  assign _T_657 = InstDecoder_1_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 145:29:@8055.4]
  assign _T_658 = InstDecoder_1_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 146:29:@8056.4]
  assign _T_659 = InstDecoder_1_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 147:29:@8057.4]
  assign _T_660 = InstDecoder_1_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 148:29:@8058.4]
  assign _T_661 = _T_660 ? InstDecoder_1_io_dinfo_imm_uj : dec_rs2_data_1; // @[Mux.scala 61:16:@8059.4]
  assign _T_662 = _T_659 ? InstDecoder_1_io_dinfo_imm_u : _T_661; // @[Mux.scala 61:16:@8060.4]
  assign _T_663 = _T_658 ? InstDecoder_1_io_dinfo_imm_sb : _T_662; // @[Mux.scala 61:16:@8061.4]
  assign _T_664 = _T_657 ? InstDecoder_1_io_dinfo_imm_s : _T_663; // @[Mux.scala 61:16:@8062.4]
  assign dec_op2_data_1 = _T_656 ? InstDecoder_1_io_dinfo_imm_i : _T_664; // @[Mux.scala 61:16:@8063.4]
  assign _T_671 = InstDecoder_1_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 154:52:@8071.6]
  assign _T_672 = InstDecoder_1_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 154:86:@8072.6]
  assign _T_673 = _T_671 | _T_672; // @[BackEnd.scala 154:62:@8073.6]
  assign _T_675 = InstDecoder_1_io_rs1_addr == 5'h0; // @[BackEnd.scala 155:47:@8074.6]
  assign _T_676 = _T_673 & _T_675; // @[BackEnd.scala 154:97:@8075.6]
  assign _T_677 = _T_676 ? 3'h5 : InstDecoder_1_io_cinfo_csr_cmd; // @[BackEnd.scala 154:29:@8076.6]
  assign rs1_addr_N0_0 = InstDecoder_io_rs1_addr != 5'h0; // @[BackEnd.scala 388:41:@8638.4]
  assign _T_1048 = _T_549 & rs1_addr_N0_0; // @[BackEnd.scala 391:42:@8643.4]
  assign _T_1049 = _T_1048 & dec_wire_0_rs1_oen; // @[BackEnd.scala 391:60:@8644.4]
  assign _T_1041 = exe_0_mem_fcn == 1'h0; // @[BackEnd.scala 387:62:@8635.4]
  assign exe_load_inst_0 = exe_wire_0_mem_en & _T_1041; // @[BackEnd.scala 387:44:@8636.4]
  assign _T_1050 = _T_1049 & exe_load_inst_0; // @[BackEnd.scala 391:83:@8645.4]
  assign rs2_addr_N0_0 = InstDecoder_io_rs2_addr != 5'h0; // @[BackEnd.scala 389:41:@8640.4]
  assign _T_1052 = _T_567 & rs2_addr_N0_0; // @[BackEnd.scala 392:42:@8647.4]
  assign _T_1053 = _T_1052 & dec_wire_0_rs2_oen; // @[BackEnd.scala 392:60:@8648.4]
  assign _T_1054 = _T_1053 & exe_load_inst_0; // @[BackEnd.scala 392:83:@8649.4]
  assign _T_1055 = _T_1050 | _T_1054; // @[BackEnd.scala 391:104:@8650.4]
  assign _T_1057 = _T_547 & rs1_addr_N0_0; // @[BackEnd.scala 393:42:@8652.4]
  assign _T_1058 = _T_1057 & dec_wire_0_rs1_oen; // @[BackEnd.scala 393:60:@8653.4]
  assign _T_1066 = exe_1_mem_fcn == 1'h0; // @[BackEnd.scala 387:62:@8662.4]
  assign exe_load_inst_1 = exe_wire_1_mem_en & _T_1066; // @[BackEnd.scala 387:44:@8663.4]
  assign _T_1059 = _T_1058 & exe_load_inst_1; // @[BackEnd.scala 393:83:@8654.4]
  assign _T_1060 = _T_1055 | _T_1059; // @[BackEnd.scala 392:104:@8655.4]
  assign _T_1062 = _T_565 & rs2_addr_N0_0; // @[BackEnd.scala 394:42:@8657.4]
  assign _T_1063 = _T_1062 & dec_wire_0_rs2_oen; // @[BackEnd.scala 394:60:@8658.4]
  assign _T_1064 = _T_1063 & exe_load_inst_1; // @[BackEnd.scala 394:83:@8659.4]
  assign rAW_0 = _T_1060 | _T_1064; // @[BackEnd.scala 393:104:@8660.4]
  assign exe_wire_0_csr_cmd = exe_valid_0 ? exe_0_csr_cmd : 3'h0; // @[BackEnd.scala 206:31:@8159.4]
  assign _T_1091 = exe_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 397:56:@8689.4]
  assign _T_1092 = rAW_0 | _T_1091; // @[BackEnd.scala 397:33:@8690.4]
  assign exe_wire_1_csr_cmd = exe_valid_1 ? exe_1_csr_cmd : 3'h0; // @[BackEnd.scala 206:31:@8196.4]
  assign _T_1093 = exe_wire_1_csr_cmd != 3'h0; // @[BackEnd.scala 397:89:@8691.4]
  assign stall_0_0 = _T_1092 | _T_1093; // @[BackEnd.scala 397:66:@8692.4]
  assign _T_689 = stall_0_0 | stall_1_1; // @[BackEnd.scala 184:31:@8110.4]
  assign _T_695 = _T_689 & _T_600; // @[BackEnd.scala 184:79:@8114.4]
  assign ma_jump = mem_sel_0 ? mem_wire_jump_0 : mem_wire_jump_1; // @[BackEnd.scala 334:29:@8510.4]
  assign mem_en = mem_sel_0 ? mem_wire_0_mem_en : mem_wire_1_mem_en; // @[BackEnd.scala 316:25:@8398.4]
  assign mem_fcn = mem_sel_0 ? mem_0_mem_fcn : mem_1_mem_fcn; // @[BackEnd.scala 317:25:@8399.4]
  assign _T_901 = mem_fcn == 1'h0; // @[BackEnd.scala 332:44:@8504.4]
  assign _T_902 = mem_en & _T_901; // @[BackEnd.scala 332:33:@8505.4]
  assign mem_typ = mem_sel_0 ? mem_0_mem_typ : mem_1_mem_typ; // @[BackEnd.scala 318:25:@8400.4]
  assign _T_890 = mem_typ[1:0]; // @[BackEnd.scala 327:43:@8496.4]
  assign _T_900 = 2'h2 == _T_890; // @[Mux.scala 46:19:@8502.4]
  assign mem_exe_out = mem_sel_0 ? mem_reg_wbdata_0 : mem_reg_wbdata_1; // @[BackEnd.scala 312:25:@8394.4]
  assign _T_893 = mem_exe_out[0]; // @[BackEnd.scala 328:23:@8497.4]
  assign _T_898 = 2'h3 == _T_890; // @[Mux.scala 46:19:@8500.4]
  assign _T_895 = mem_exe_out[1:0]; // @[BackEnd.scala 329:23:@8498.4]
  assign _T_897 = _T_895 != 2'h0; // @[BackEnd.scala 329:29:@8499.4]
  assign _T_899 = _T_898 ? _T_897 : 1'h0; // @[Mux.scala 46:16:@8501.4]
  assign ls_addr_ma_valid = _T_900 ? _T_893 : _T_899; // @[Mux.scala 46:16:@8503.4]
  assign ma_load = _T_902 & ls_addr_ma_valid; // @[BackEnd.scala 332:54:@8506.4]
  assign _T_922 = ma_jump | ma_load; // @[BackEnd.scala 349:25:@8526.4]
  assign _T_904 = mem_en & mem_fcn; // @[BackEnd.scala 333:33:@8508.4]
  assign ma_store = _T_904 & ls_addr_ma_valid; // @[BackEnd.scala 333:54:@8509.4]
  assign _T_923 = _T_922 | ma_store; // @[BackEnd.scala 349:36:@8527.4]
  assign ma_illegal = mem_sel_0 ? mem_wire_0_illegal : mem_wire_1_illegal; // @[BackEnd.scala 335:29:@8511.4]
  assign _T_924 = _T_923 | ma_illegal; // @[BackEnd.scala 349:48:@8528.4]
  assign xcpt_valid = _T_924 | csr_io_eret; // @[BackEnd.scala 349:62:@8529.4]
  assign _T_696 = _T_695 | xcpt_valid; // @[BackEnd.scala 184:104:@8115.4]
  assign not_expect = io_front_feedBack_tgt != exe_btb_tgt; // @[BackEnd.scala 256:48:@8279.4]
  assign exe_wire_0_bj_sel = exe_valid_0 & exe_0_bj_sel; // @[BackEnd.scala 208:41:@8163.4]
  assign exe_wire_1_bj_sel = exe_valid_1 & exe_1_bj_sel; // @[BackEnd.scala 208:41:@8200.4]
  assign exe_bj_valid = exe_wire_0_bj_sel | exe_wire_1_bj_sel; // @[BackEnd.scala 198:56:@8148.4]
  assign mispredict = not_expect & exe_bj_valid; // @[BackEnd.scala 257:28:@8280.4]
  assign _T_704 = mispredict == 1'h0; // @[BackEnd.scala 187:47:@8124.8]
  assign _T_705 = io_front_inst_0_valid & _T_704; // @[BackEnd.scala 187:44:@8125.8]
  assign _GEN_39 = _T_601 ? _T_705 : exe_valid_0; // @[BackEnd.scala 186:60:@8123.6]
  assign _GEN_40 = _T_696 ? 1'h0 : _GEN_39; // @[BackEnd.scala 184:119:@8116.4]
  assign _T_1095 = InstDecoder_io_wbaddr == InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 400:20:@8694.4]
  assign rs1_addr_N0_1 = InstDecoder_1_io_rs1_addr != 5'h0; // @[BackEnd.scala 388:41:@8665.4]
  assign _T_1096 = _T_1095 & rs1_addr_N0_1; // @[BackEnd.scala 400:40:@8695.4]
  assign _T_1097 = _T_1096 & dec_wire_1_rs1_oen; // @[BackEnd.scala 400:58:@8696.4]
  assign _T_1098 = _T_1097 & dec_wire_0_rf_wen; // @[BackEnd.scala 400:81:@8697.4]
  assign _T_1099 = InstDecoder_io_wbaddr == InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 401:20:@8698.4]
  assign rs2_addr_N0_1 = InstDecoder_1_io_rs2_addr != 5'h0; // @[BackEnd.scala 389:41:@8667.4]
  assign _T_1100 = _T_1099 & rs2_addr_N0_1; // @[BackEnd.scala 401:40:@8699.4]
  assign _T_1101 = _T_1100 & dec_wire_1_rs2_oen; // @[BackEnd.scala 401:58:@8700.4]
  assign _T_1102 = _T_1101 & dec_wire_0_rf_wen; // @[BackEnd.scala 401:81:@8701.4]
  assign _T_1103 = _T_1098 | _T_1102; // @[BackEnd.scala 400:104:@8702.4]
  assign _T_1104 = dec_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 402:25:@8703.4]
  assign _T_1105 = _T_1103 | _T_1104; // @[BackEnd.scala 401:104:@8704.4]
  assign _T_1073 = _T_618 & rs1_addr_N0_1; // @[BackEnd.scala 391:42:@8670.4]
  assign _T_1074 = _T_1073 & dec_wire_1_rs1_oen; // @[BackEnd.scala 391:60:@8671.4]
  assign _T_1075 = _T_1074 & exe_load_inst_0; // @[BackEnd.scala 391:83:@8672.4]
  assign _T_1077 = _T_636 & rs2_addr_N0_1; // @[BackEnd.scala 392:42:@8674.4]
  assign _T_1078 = _T_1077 & dec_wire_1_rs2_oen; // @[BackEnd.scala 392:60:@8675.4]
  assign _T_1079 = _T_1078 & exe_load_inst_0; // @[BackEnd.scala 392:83:@8676.4]
  assign _T_1080 = _T_1075 | _T_1079; // @[BackEnd.scala 391:104:@8677.4]
  assign _T_1082 = _T_616 & rs1_addr_N0_1; // @[BackEnd.scala 393:42:@8679.4]
  assign _T_1083 = _T_1082 & dec_wire_1_rs1_oen; // @[BackEnd.scala 393:60:@8680.4]
  assign _T_1084 = _T_1083 & exe_load_inst_1; // @[BackEnd.scala 393:83:@8681.4]
  assign _T_1085 = _T_1080 | _T_1084; // @[BackEnd.scala 392:104:@8682.4]
  assign _T_1087 = _T_634 & rs2_addr_N0_1; // @[BackEnd.scala 394:42:@8684.4]
  assign _T_1088 = _T_1087 & dec_wire_1_rs2_oen; // @[BackEnd.scala 394:60:@8685.4]
  assign _T_1089 = _T_1088 & exe_load_inst_1; // @[BackEnd.scala 394:83:@8686.4]
  assign rAW_1 = _T_1085 | _T_1089; // @[BackEnd.scala 393:104:@8687.4]
  assign _T_1106 = _T_1105 | rAW_1; // @[BackEnd.scala 402:35:@8705.4]
  assign stall_1_0 = _T_1106 | stall_0_0; // @[BackEnd.scala 402:45:@8706.4]
  assign _T_708 = stall_1_0 & _T_598; // @[BackEnd.scala 190:30:@8129.4]
  assign _T_711 = _T_708 & _T_600; // @[BackEnd.scala 190:54:@8131.4]
  assign _T_712 = _T_711 | xcpt_valid; // @[BackEnd.scala 190:79:@8132.4]
  assign exe_cancel = not_expect & exe_wire_0_bj_sel; // @[BackEnd.scala 258:28:@8282.4]
  assign _T_713 = _T_712 | exe_cancel; // @[BackEnd.scala 190:93:@8133.4]
  assign _T_722 = io_front_inst_1_valid & _T_704; // @[BackEnd.scala 193:44:@8143.8]
  assign _T_724 = io_front_split == 1'h0; // @[BackEnd.scala 193:62:@8144.8]
  assign _T_725 = _T_722 & _T_724; // @[BackEnd.scala 193:59:@8145.8]
  assign _GEN_41 = _T_601 ? _T_725 : exe_valid_1; // @[BackEnd.scala 192:60:@8141.6]
  assign _GEN_42 = _T_713 ? 1'h0 : _GEN_41; // @[BackEnd.scala 190:108:@8134.4]
  assign exe_wire_branch = exe_bj_valid & exe_branch; // @[BackEnd.scala 199:38:@8149.4]
  assign exe_wire_call = exe_bj_valid & exe_call; // @[BackEnd.scala 200:38:@8150.4]
  assign exe_wire_retn = exe_bj_valid & exe_retn; // @[BackEnd.scala 201:38:@8151.4]
  assign target_brjmp = exe_wire_0_bj_sel ? ALU_io_target_brjmp : ALU_1_io_target_brjmp; // @[BackEnd.scala 237:19:@8227.4]
  assign target_jpreg = exe_wire_0_bj_sel ? ALU_io_target_jpreg : ALU_1_io_target_jpreg; // @[BackEnd.scala 237:19:@8227.4]
  assign target_conti = exe_wire_0_bj_sel ? ALU_io_target_conti : ALU_1_io_target_conti; // @[BackEnd.scala 237:19:@8227.4]
  assign pc_sel = exe_wire_0_bj_sel ? ALU_io_ctrl_pc_sel : ALU_1_io_ctrl_pc_sel; // @[BackEnd.scala 238:19:@8228.4]
  assign _GEN_67 = exe_wire_retn ? 1'h0 : _T_759; // @[BackEnd.scala 64:20:@8235.6]
  assign _GEN_68 = _T_600 ? 1'h1 : _GEN_67; // @[BackEnd.scala 63:20:@8231.4]
  assign _GEN_69 = exe_wire_call ? 1'h0 : _T_767; // @[BackEnd.scala 64:20:@8246.6]
  assign _GEN_70 = _T_600 ? 1'h1 : _GEN_69; // @[BackEnd.scala 63:20:@8242.4]
  assign _GEN_71 = exe_bj_valid ? 1'h0 : _T_775; // @[BackEnd.scala 64:20:@8258.6]
  assign _GEN_72 = _T_600 ? 1'h1 : _GEN_71; // @[BackEnd.scala 63:20:@8254.4]
  assign _T_779 = pc_sel == 2'h1; // @[BackEnd.scala 244:40:@8263.4]
  assign _T_780 = pc_sel == 2'h2; // @[BackEnd.scala 244:63:@8264.4]
  assign _T_784 = _T_780 ? target_jpreg : target_conti; // @[BackEnd.scala 247:8:@8269.4]
  assign _T_790 = exe_wire_retn ? 2'h1 : 2'h3; // @[BackEnd.scala 254:8:@8276.4]
  assign _T_802 = _T_779 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@8289.6]
  assign _T_803 = _T_802 & target_brjmp; // @[BackEnd.scala 263:47:@8290.6]
  assign _T_808 = _T_780 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@8293.6]
  assign _T_809 = _T_808 & target_jpreg; // @[BackEnd.scala 264:47:@8294.6]
  assign _T_810 = _T_803 | _T_809; // @[BackEnd.scala 263:63:@8295.6]
  assign _GEN_73 = _T_600 ? _T_810 : mem_reg_jpnpc; // @[BackEnd.scala 261:31:@8286.4]
  assign _T_813 = stall_0_2 == 1'h0; // @[BackEnd.scala 267:57:@8299.4]
  assign _T_814 = stall_1_2 & _T_813; // @[BackEnd.scala 267:54:@8300.4]
  assign _T_815 = _T_814 | xcpt_valid; // @[BackEnd.scala 267:78:@8301.4]
  assign _GEN_74 = _T_600 ? exe_valid_0 : mem_valid_0; // @[BackEnd.scala 269:37:@8307.6]
  assign _GEN_75 = _T_815 ? 1'h0 : _GEN_74; // @[BackEnd.scala 267:93:@8302.4]
  assign _T_821 = stall_1_1 & _T_600; // @[BackEnd.scala 273:30:@8311.4]
  assign _T_822 = _T_821 | xcpt_valid; // @[BackEnd.scala 273:55:@8312.4]
  assign _T_827 = exe_cancel == 1'h0; // @[BackEnd.scala 276:37:@8319.8]
  assign _T_828 = exe_valid_1 & _T_827; // @[BackEnd.scala 276:34:@8320.8]
  assign _GEN_76 = _T_600 ? _T_828 : mem_valid_1; // @[BackEnd.scala 275:37:@8318.6]
  assign _GEN_77 = _T_822 ? 1'h0 : _GEN_76; // @[BackEnd.scala 273:70:@8313.4]
  assign _T_831 = exe_wire_1_mem_en & _T_827; // @[BackEnd.scala 279:69:@8324.4]
  assign mem_inst = mem_sel_0 ? mem_0_inst : mem_1_inst; // @[BackEnd.scala 311:25:@8393.4]
  assign _T_905 = ma_load | ma_store; // @[BackEnd.scala 336:27:@8512.4]
  assign _T_906 = _T_905 | ma_jump; // @[BackEnd.scala 336:39:@8513.4]
  assign _T_913 = ma_store ? 3'h6 : 3'h0; // @[Mux.scala 61:16:@8516.4]
  assign _T_914 = ma_load ? 3'h4 : _T_913; // @[Mux.scala 61:16:@8517.4]
  assign _T_915 = ma_illegal ? 3'h2 : _T_914; // @[Mux.scala 61:16:@8518.4]
  assign _T_916 = ma_jump ? 3'h0 : _T_915; // @[Mux.scala 61:16:@8519.4]
  assign _T_918 = ma_store ? mem_exe_out : 32'h0; // @[Mux.scala 61:16:@8521.4]
  assign _T_919 = ma_load ? mem_exe_out : _T_918; // @[Mux.scala 61:16:@8522.4]
  assign _T_920 = ma_illegal ? mem_inst : _T_919; // @[Mux.scala 61:16:@8523.4]
  assign _T_926 = xcpt_valid & mem_sel_0; // @[BackEnd.scala 352:44:@8532.4]
  assign _T_927 = stall_0_2 | _T_926; // @[BackEnd.scala 352:29:@8533.4]
  assign _GEN_78 = _T_927 ? 1'h0 : mem_valid_0; // @[BackEnd.scala 352:60:@8534.4]
  assign _T_929 = stall_1_2 | xcpt_valid; // @[BackEnd.scala 356:29:@8540.4]
  assign _GEN_79 = _T_929 ? 1'h0 : mem_valid_1; // @[BackEnd.scala 356:44:@8541.4]
  assign _T_946 = {wb_valid_1,wb_valid_0}; // @[BackEnd.scala 375:25:@8562.4]
  assign retire_0 = ^_T_946; // @[BackEnd.scala 375:32:@8563.4]
  assign _T_949 = ~ _T_946; // @[BackEnd.scala 376:32:@8566.4]
  assign retire_1 = _T_949 == 2'h0; // @[BackEnd.scala 376:32:@8567.4]
  assign _GEN_80 = mispredict ? 1'h0 : _T_1127; // @[BackEnd.scala 64:20:@8729.6]
  assign _GEN_81 = _T_600 ? 1'h1 : _GEN_80; // @[BackEnd.scala 63:20:@8725.4]
  assign _T_1132 = stall_0_0 == 1'h0; // @[BackEnd.scala 411:26:@8736.4]
  assign _T_1135 = _T_1132 & _T_598; // @[BackEnd.scala 411:47:@8738.4]
  assign _T_1140 = stall_1_0 == 1'h0; // @[BackEnd.scala 412:26:@8742.4]
  assign _T_1143 = _T_1140 & _T_598; // @[BackEnd.scala 412:47:@8744.4]
  assign _T_1149 = stall_0_2 ? 8'h4d : 8'h20; // @[BackEnd.scala 421:12:@8748.4]
  assign _T_1157 = stall_0_0 ? 8'h44 : 8'h20; // @[BackEnd.scala 423:12:@8750.4]
  assign _T_1160 = ALU_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 424:32:@8751.4]
  assign _T_1163 = ALU_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 425:32:@8752.4]
  assign _T_1166 = ALU_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 426:32:@8753.4]
  assign _T_1169 = ALU_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 427:32:@8754.4]
  assign _T_1172 = _T_1169 ? 8'h20 : 8'h3f; // @[BackEnd.scala 427:12:@8755.4]
  assign _T_1173 = _T_1166 ? 8'h45 : _T_1172; // @[BackEnd.scala 426:12:@8756.4]
  assign _T_1174 = _T_1163 ? 8'h4a : _T_1173; // @[BackEnd.scala 425:12:@8757.4]
  assign _T_1175 = _T_1160 ? 8'h42 : _T_1174; // @[BackEnd.scala 424:12:@8758.4]
  assign _T_1179 = csr_io_illegal ? 8'h58 : 8'h20; // @[BackEnd.scala 428:12:@8759.4]
  assign _T_1182 = exe_valid_0 == 1'h0; // @[BackEnd.scala 429:13:@8760.4]
  assign _T_1183 = _T_1182 | xcpt_valid; // @[BackEnd.scala 429:27:@8761.4]
  assign _T_1189 = _T_1183 | stall_1_2; // @[BackEnd.scala 429:72:@8765.4]
  assign _T_1195 = _T_1189 ? 32'h4033 : exe_0_inst; // @[BackEnd.scala 429:12:@8769.4]
  assign _T_1198 = reset == 1'h0; // @[BackEnd.scala 416:11:@8771.4]
  assign _T_1201 = stall_1_2 ? 8'h4d : 8'h20; // @[BackEnd.scala 421:12:@8775.4]
  assign _T_1205 = stall_1_1 ? 8'h45 : 8'h20; // @[BackEnd.scala 422:12:@8776.4]
  assign _T_1209 = stall_1_0 ? 8'h44 : 8'h20; // @[BackEnd.scala 423:12:@8777.4]
  assign _T_1212 = ALU_1_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 424:32:@8778.4]
  assign _T_1215 = ALU_1_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 425:32:@8779.4]
  assign _T_1218 = ALU_1_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 426:32:@8780.4]
  assign _T_1221 = ALU_1_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 427:32:@8781.4]
  assign _T_1224 = _T_1221 ? 8'h20 : 8'h3f; // @[BackEnd.scala 427:12:@8782.4]
  assign _T_1225 = _T_1218 ? 8'h45 : _T_1224; // @[BackEnd.scala 426:12:@8783.4]
  assign _T_1226 = _T_1215 ? 8'h4a : _T_1225; // @[BackEnd.scala 425:12:@8784.4]
  assign _T_1227 = _T_1212 ? 8'h42 : _T_1226; // @[BackEnd.scala 424:12:@8785.4]
  assign _T_1234 = exe_valid_1 == 1'h0; // @[BackEnd.scala 429:13:@8787.4]
  assign _T_1235 = _T_1234 | xcpt_valid; // @[BackEnd.scala 429:27:@8788.4]
  assign _T_1240 = _T_1235 | exe_cancel; // @[BackEnd.scala 429:41:@8791.4]
  assign _T_1241 = _T_1240 | stall_1_2; // @[BackEnd.scala 429:72:@8792.4]
  assign _T_1246 = _T_1241 | stall_1_1; // @[BackEnd.scala 430:29:@8795.4]
  assign _T_1247 = _T_1246 ? 32'h4033 : exe_1_inst; // @[BackEnd.scala 429:12:@8796.4]
  assign _T_1257 = exe_wire_0_bj_sel ? exe_0_inst : exe_1_inst; // @[BackEnd.scala 452:12:@8817.6]
  assign io_mem_req_valid = exe_wire_0_mem_en | _T_831; // @[BackEnd.scala 279:24:@8326.4]
  assign io_mem_req_bits_addr = exe_wire_0_mem_en ? exe_wbdata_0 : exe_wbdata_1; // @[BackEnd.scala 280:24:@8328.4]
  assign io_mem_req_bits_data = exe_wire_0_mem_en ? exe_0_rs2_data : exe_1_rs2_data; // @[BackEnd.scala 283:24:@8334.4]
  assign io_mem_req_bits_fcn = exe_wire_0_mem_en ? exe_0_mem_fcn : exe_1_mem_fcn; // @[BackEnd.scala 281:24:@8330.4]
  assign io_mem_req_bits_typ = exe_wire_0_mem_en ? exe_0_mem_typ : exe_1_mem_typ; // @[BackEnd.scala 282:24:@8332.4]
  assign io_cyc = csr_io_time; // @[BackEnd.scala 80:10:@7869.4]
  assign io_front_xcpt_valid = _T_924 | csr_io_eret; // @[BackEnd.scala 410:17:@8735.4]
  assign io_front_xcpt_bits = csr_io_evec; // @[BackEnd.scala 410:17:@8734.4]
  assign io_front_kill = mispredict & _T_1127; // @[BackEnd.scala 409:17:@8733.4]
  assign io_front_forward_0 = _T_1135 & _T_600; // @[BackEnd.scala 411:23:@8741.4]
  assign io_front_forward_1 = _T_1143 & _T_600; // @[BackEnd.scala 412:23:@8747.4]
  assign io_front_ras_pop = exe_wire_retn & _T_759; // @[BackEnd.scala 240:20:@8239.4]
  assign io_front_ras_push_valid = exe_wire_call & _T_767; // @[BackEnd.scala 241:27:@8250.4]
  assign io_front_ras_push_bits = exe_wire_0_bj_sel ? ALU_io_target_conti : ALU_1_io_target_conti; // @[BackEnd.scala 242:27:@8251.4]
  assign io_front_fb_pc = exe_wire_0_bj_sel ? exe_0_pc : exe_1_pc; // @[BackEnd.scala 252:18:@8275.4]
  assign io_front_fb_type = exe_wire_branch ? 2'h2 : _T_790; // @[BackEnd.scala 253:20:@8278.4]
  assign io_front_feedBack_redirect = _T_779 | _T_780; // @[BackEnd.scala 244:30:@8266.4]
  assign io_front_feedBack_history = exe_btb_history; // @[BackEnd.scala 250:30:@8272.4]
  assign io_front_feedBack_diff = exe_btb_diff; // @[BackEnd.scala 251:30:@8273.4]
  assign io_front_feedBack_tgt = _T_779 ? target_brjmp : _T_784; // @[BackEnd.scala 245:25:@8271.4]
  assign io_front_feedBack_valid = exe_bj_valid & _T_775; // @[BackEnd.scala 243:27:@8262.4]
  assign csr_clock = clock; // @[:@7851.4]
  assign csr_reset = reset; // @[:@7852.4]
  assign csr_io_rw_cmd = mem_sel_0 ? mem_wire_0_csr_cmd : mem_wire_1_csr_cmd; // @[BackEnd.scala 324:19:@8494.4]
  assign csr_io_rw_addr = mem_inst[31:20]; // @[BackEnd.scala 322:19:@8492.4]
  assign csr_io_rw_wdata = mem_sel_0 ? mem_reg_wbdata_0 : mem_reg_wbdata_1; // @[BackEnd.scala 323:19:@8493.4]
  assign csr_io_xcpt = _T_906 | ma_illegal; // @[BackEnd.scala 336:16:@8515.4]
  assign csr_io_cause = {{29'd0}, _T_916}; // @[BackEnd.scala 337:16:@8520.4]
  assign csr_io_tval = ma_jump ? mem_reg_jpnpc : _T_920; // @[BackEnd.scala 343:16:@8525.4]
  assign csr_io_illegal = 1'h0;
  assign csr_io_retire = {retire_1,retire_0}; // @[BackEnd.scala 377:17:@8570.4]
  assign csr_io_pc = mem_sel_0 ? mem_0_pc : mem_1_pc; // @[BackEnd.scala 325:19:@8495.4]
  assign regfile_clock = clock; // @[:@7854.4]
  assign regfile_io_rs1_addr_0 = InstDecoder_io_rs1_addr; // @[BackEnd.scala 116:28:@7911.4]
  assign regfile_io_rs1_addr_1 = InstDecoder_1_io_rs1_addr; // @[BackEnd.scala 116:28:@8007.4]
  assign regfile_io_rs2_addr_0 = InstDecoder_io_rs2_addr; // @[BackEnd.scala 117:28:@7912.4]
  assign regfile_io_rs2_addr_1 = InstDecoder_1_io_rs2_addr; // @[BackEnd.scala 117:28:@8008.4]
  assign regfile_io_waddr_0 = wb_0_wbaddr; // @[BackEnd.scala 364:25:@8551.4]
  assign regfile_io_waddr_1 = wb_1_wbaddr; // @[BackEnd.scala 364:25:@8558.4]
  assign regfile_io_wdata_0 = wb_wbdata_0; // @[BackEnd.scala 365:25:@8552.4]
  assign regfile_io_wdata_1 = wb_wbdata_1; // @[BackEnd.scala 365:25:@8559.4]
  assign regfile_io_wen_0 = _T_931 & _T_933; // @[BackEnd.scala 366:25:@8553.4]
  assign regfile_io_wen_1 = _T_935 & _T_937; // @[BackEnd.scala 366:25:@8560.4]
  assign ALU_io_op1 = exe_0_op1_data; // @[BackEnd.scala 211:25:@8167.4]
  assign ALU_io_op2 = exe_0_op2_data; // @[BackEnd.scala 212:25:@8168.4]
  assign ALU_io_pc = exe_0_pc; // @[BackEnd.scala 213:25:@8169.4]
  assign ALU_io_ctrl_fun = exe_0_alu_fun; // @[BackEnd.scala 215:25:@8171.4]
  assign ALU_io_ctrl_br_type = exe_valid_0 ? exe_0_br_type : 4'h0; // @[BackEnd.scala 216:25:@8172.4]
  assign ALU_io_ctrl_wb_sel = exe_0_wb_sel; // @[BackEnd.scala 217:25:@8173.4]
  assign ALU_io_rs2_data = exe_0_rs2_data; // @[BackEnd.scala 214:25:@8170.4]
  assign ALU_1_io_op1 = exe_1_op1_data; // @[BackEnd.scala 211:25:@8204.4]
  assign ALU_1_io_op2 = exe_1_op2_data; // @[BackEnd.scala 212:25:@8205.4]
  assign ALU_1_io_pc = exe_1_pc; // @[BackEnd.scala 213:25:@8206.4]
  assign ALU_1_io_ctrl_fun = exe_1_alu_fun; // @[BackEnd.scala 215:25:@8208.4]
  assign ALU_1_io_ctrl_br_type = exe_valid_1 ? exe_1_br_type : 4'h0; // @[BackEnd.scala 216:25:@8209.4]
  assign ALU_1_io_ctrl_wb_sel = exe_1_wb_sel; // @[BackEnd.scala 217:25:@8210.4]
  assign ALU_1_io_rs2_data = exe_1_rs2_data; // @[BackEnd.scala 214:25:@8207.4]
  assign InstDecoder_io_inst = io_front_inst_0_bits; // @[BackEnd.scala 110:18:@7900.4]
  assign InstDecoder_1_io_inst = io_front_inst_1_bits; // @[BackEnd.scala 110:18:@7996.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exe_0_rf_wen = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  exe_0_wbaddr = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  exe_0_mem_en = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  exe_0_csr_cmd = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  exe_0_illegal = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  exe_0_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  exe_0_inst = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  exe_0_rs2_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  exe_0_wb_sel = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  exe_0_mem_fcn = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  exe_0_mem_typ = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  exe_0_br_type = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  exe_0_bj_sel = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  exe_0_op1_data = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  exe_0_op2_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  exe_0_alu_fun = _RAND_15[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  exe_1_rf_wen = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  exe_1_wbaddr = _RAND_17[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  exe_1_mem_en = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  exe_1_csr_cmd = _RAND_19[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  exe_1_illegal = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  exe_1_pc = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  exe_1_inst = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  exe_1_rs2_data = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  exe_1_wb_sel = _RAND_24[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  exe_1_mem_fcn = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  exe_1_mem_typ = _RAND_26[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  exe_1_br_type = _RAND_27[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  exe_1_bj_sel = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  exe_1_op1_data = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  exe_1_op2_data = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  exe_1_alu_fun = _RAND_31[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  exe_valid_0 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  exe_valid_1 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mem_0_rf_wen = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  mem_0_wbaddr = _RAND_35[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_0_mem_en = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_0_csr_cmd = _RAND_37[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mem_0_illegal = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  mem_0_pc = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  mem_0_inst = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  mem_0_wb_sel = _RAND_41[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  mem_0_mem_fcn = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  mem_0_mem_typ = _RAND_43[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  mem_1_rf_wen = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  mem_1_wbaddr = _RAND_45[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  mem_1_mem_en = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  mem_1_csr_cmd = _RAND_47[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  mem_1_illegal = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  mem_1_pc = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  mem_1_inst = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  mem_1_wb_sel = _RAND_51[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_1_mem_fcn = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_1_mem_typ = _RAND_53[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_valid_0 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_valid_1 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  wb_0_rf_wen = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  wb_0_wbaddr = _RAND_57[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  wb_1_rf_wen = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  wb_1_wbaddr = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  wb_valid_0 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  wb_valid_1 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  wb_wbdata_0 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  wb_wbdata_1 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  mem_reg_wbdata_0 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  mem_reg_wbdata_1 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_reg_jpnpc = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  exe_btb_redirect = _RAND_67[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  exe_btb_history = _RAND_68[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  exe_btb_diff = _RAND_69[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  exe_btb_tgt = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  exe_branch = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  exe_call = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  exe_retn = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_759 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_767 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_775 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  _T_1127 = _RAND_77[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_601) begin
      exe_0_rf_wen <= InstDecoder_io_cinfo_rf_wen;
    end
    if (_T_601) begin
      exe_0_wbaddr <= InstDecoder_io_wbaddr;
    end
    if (_T_601) begin
      exe_0_mem_en <= InstDecoder_io_cinfo_mem_en;
    end
    if (_T_601) begin
      if (_T_607) begin
        exe_0_csr_cmd <= 3'h5;
      end else begin
        exe_0_csr_cmd <= InstDecoder_io_cinfo_csr_cmd;
      end
    end
    if (_T_601) begin
      exe_0_illegal <= InstDecoder_io_cinfo_illegal;
    end
    if (_T_601) begin
      exe_0_pc <= io_front_pc_0;
    end
    if (_T_601) begin
      exe_0_inst <= InstDecoder_io_inst;
    end
    if (_T_601) begin
      if (_T_566) begin
        exe_0_rs2_data <= exe_wbdata_1;
      end else begin
        if (_T_568) begin
          exe_0_rs2_data <= exe_wbdata_0;
        end else begin
          if (_T_570) begin
            if (_T_885) begin
              exe_0_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_886) begin
                exe_0_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_0_rs2_data <= mem_reg_wbdata_1;
              end
            end
          end else begin
            if (_T_572) begin
              if (_T_866) begin
                exe_0_rs2_data <= io_mem_resp_bits_data;
              end else begin
                if (_T_867) begin
                  exe_0_rs2_data <= csr_io_rw_rdata;
                end else begin
                  exe_0_rs2_data <= mem_reg_wbdata_0;
                end
              end
            end else begin
              if (_T_574) begin
                exe_0_rs2_data <= wb_wbdata_1;
              end else begin
                if (_T_576) begin
                  exe_0_rs2_data <= wb_wbdata_0;
                end else begin
                  exe_0_rs2_data <= rf_rs2_data_0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      exe_0_wb_sel <= InstDecoder_io_cinfo_wb_sel;
    end
    if (_T_601) begin
      exe_0_mem_fcn <= InstDecoder_io_cinfo_mem_fcn;
    end
    if (_T_601) begin
      exe_0_mem_typ <= InstDecoder_io_cinfo_mem_typ;
    end
    if (_T_601) begin
      exe_0_br_type <= InstDecoder_io_cinfo_br_type;
    end
    if (_T_601) begin
      exe_0_bj_sel <= io_front_bj_sel_0;
    end
    if (_T_601) begin
      if (_T_583) begin
        exe_0_op1_data <= InstDecoder_io_dinfo_imm_z;
      end else begin
        if (_T_584) begin
          exe_0_op1_data <= io_front_pc_0;
        end else begin
          if (_T_548) begin
            exe_0_op1_data <= exe_wbdata_1;
          end else begin
            if (_T_550) begin
              exe_0_op1_data <= exe_wbdata_0;
            end else begin
              if (_T_552) begin
                if (_T_885) begin
                  exe_0_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_886) begin
                    exe_0_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_0_op1_data <= mem_reg_wbdata_1;
                  end
                end
              end else begin
                if (_T_554) begin
                  if (_T_866) begin
                    exe_0_op1_data <= io_mem_resp_bits_data;
                  end else begin
                    if (_T_867) begin
                      exe_0_op1_data <= csr_io_rw_rdata;
                    end else begin
                      exe_0_op1_data <= mem_reg_wbdata_0;
                    end
                  end
                end else begin
                  if (_T_556) begin
                    exe_0_op1_data <= wb_wbdata_1;
                  end else begin
                    if (_T_558) begin
                      exe_0_op1_data <= wb_wbdata_0;
                    end else begin
                      exe_0_op1_data <= rf_rs1_data_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      if (_T_587) begin
        exe_0_op2_data <= InstDecoder_io_dinfo_imm_i;
      end else begin
        if (_T_588) begin
          exe_0_op2_data <= InstDecoder_io_dinfo_imm_s;
        end else begin
          if (_T_589) begin
            exe_0_op2_data <= InstDecoder_io_dinfo_imm_sb;
          end else begin
            if (_T_590) begin
              exe_0_op2_data <= InstDecoder_io_dinfo_imm_u;
            end else begin
              if (_T_591) begin
                exe_0_op2_data <= InstDecoder_io_dinfo_imm_uj;
              end else begin
                if (_T_566) begin
                  exe_0_op2_data <= exe_wbdata_1;
                end else begin
                  if (_T_568) begin
                    exe_0_op2_data <= exe_wbdata_0;
                  end else begin
                    if (_T_570) begin
                      if (_T_885) begin
                        exe_0_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_886) begin
                          exe_0_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_0_op2_data <= mem_reg_wbdata_1;
                        end
                      end
                    end else begin
                      if (_T_572) begin
                        if (_T_866) begin
                          exe_0_op2_data <= io_mem_resp_bits_data;
                        end else begin
                          if (_T_867) begin
                            exe_0_op2_data <= csr_io_rw_rdata;
                          end else begin
                            exe_0_op2_data <= mem_reg_wbdata_0;
                          end
                        end
                      end else begin
                        if (_T_574) begin
                          exe_0_op2_data <= wb_wbdata_1;
                        end else begin
                          if (_T_576) begin
                            exe_0_op2_data <= wb_wbdata_0;
                          end else begin
                            exe_0_op2_data <= rf_rs2_data_0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      exe_0_alu_fun <= InstDecoder_io_cinfo_alu_fun;
    end
    if (_T_601) begin
      exe_1_rf_wen <= InstDecoder_1_io_cinfo_rf_wen;
    end
    if (_T_601) begin
      exe_1_wbaddr <= InstDecoder_1_io_wbaddr;
    end
    if (_T_601) begin
      exe_1_mem_en <= InstDecoder_1_io_cinfo_mem_en;
    end
    if (_T_601) begin
      if (_T_676) begin
        exe_1_csr_cmd <= 3'h5;
      end else begin
        exe_1_csr_cmd <= InstDecoder_1_io_cinfo_csr_cmd;
      end
    end
    if (_T_601) begin
      exe_1_illegal <= InstDecoder_1_io_cinfo_illegal;
    end
    if (_T_601) begin
      exe_1_pc <= io_front_pc_1;
    end
    if (_T_601) begin
      exe_1_inst <= InstDecoder_1_io_inst;
    end
    if (_T_601) begin
      if (_T_635) begin
        exe_1_rs2_data <= exe_wbdata_1;
      end else begin
        if (_T_637) begin
          exe_1_rs2_data <= exe_wbdata_0;
        end else begin
          if (_T_639) begin
            if (_T_885) begin
              exe_1_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_886) begin
                exe_1_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_1_rs2_data <= mem_reg_wbdata_1;
              end
            end
          end else begin
            if (_T_641) begin
              if (_T_866) begin
                exe_1_rs2_data <= io_mem_resp_bits_data;
              end else begin
                if (_T_867) begin
                  exe_1_rs2_data <= csr_io_rw_rdata;
                end else begin
                  exe_1_rs2_data <= mem_reg_wbdata_0;
                end
              end
            end else begin
              if (_T_643) begin
                exe_1_rs2_data <= wb_wbdata_1;
              end else begin
                if (_T_645) begin
                  exe_1_rs2_data <= wb_wbdata_0;
                end else begin
                  exe_1_rs2_data <= rf_rs2_data_1;
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      exe_1_wb_sel <= InstDecoder_1_io_cinfo_wb_sel;
    end
    if (_T_601) begin
      exe_1_mem_fcn <= InstDecoder_1_io_cinfo_mem_fcn;
    end
    if (_T_601) begin
      exe_1_mem_typ <= InstDecoder_1_io_cinfo_mem_typ;
    end
    if (_T_601) begin
      exe_1_br_type <= InstDecoder_1_io_cinfo_br_type;
    end
    if (_T_601) begin
      exe_1_bj_sel <= io_front_bj_sel_1;
    end
    if (_T_601) begin
      if (_T_652) begin
        exe_1_op1_data <= InstDecoder_1_io_dinfo_imm_z;
      end else begin
        if (_T_653) begin
          exe_1_op1_data <= io_front_pc_1;
        end else begin
          if (_T_617) begin
            exe_1_op1_data <= exe_wbdata_1;
          end else begin
            if (_T_619) begin
              exe_1_op1_data <= exe_wbdata_0;
            end else begin
              if (_T_621) begin
                if (_T_885) begin
                  exe_1_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_886) begin
                    exe_1_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_1_op1_data <= mem_reg_wbdata_1;
                  end
                end
              end else begin
                if (_T_623) begin
                  if (_T_866) begin
                    exe_1_op1_data <= io_mem_resp_bits_data;
                  end else begin
                    if (_T_867) begin
                      exe_1_op1_data <= csr_io_rw_rdata;
                    end else begin
                      exe_1_op1_data <= mem_reg_wbdata_0;
                    end
                  end
                end else begin
                  if (_T_625) begin
                    exe_1_op1_data <= wb_wbdata_1;
                  end else begin
                    if (_T_627) begin
                      exe_1_op1_data <= wb_wbdata_0;
                    end else begin
                      exe_1_op1_data <= rf_rs1_data_1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      if (_T_656) begin
        exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_i;
      end else begin
        if (_T_657) begin
          exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_s;
        end else begin
          if (_T_658) begin
            exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_sb;
          end else begin
            if (_T_659) begin
              exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_u;
            end else begin
              if (_T_660) begin
                exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_uj;
              end else begin
                if (_T_635) begin
                  exe_1_op2_data <= exe_wbdata_1;
                end else begin
                  if (_T_637) begin
                    exe_1_op2_data <= exe_wbdata_0;
                  end else begin
                    if (_T_639) begin
                      if (_T_885) begin
                        exe_1_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_886) begin
                          exe_1_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_1_op2_data <= mem_reg_wbdata_1;
                        end
                      end
                    end else begin
                      if (_T_641) begin
                        if (_T_866) begin
                          exe_1_op2_data <= io_mem_resp_bits_data;
                        end else begin
                          if (_T_867) begin
                            exe_1_op2_data <= csr_io_rw_rdata;
                          end else begin
                            exe_1_op2_data <= mem_reg_wbdata_0;
                          end
                        end
                      end else begin
                        if (_T_643) begin
                          exe_1_op2_data <= wb_wbdata_1;
                        end else begin
                          if (_T_645) begin
                            exe_1_op2_data <= wb_wbdata_0;
                          end else begin
                            exe_1_op2_data <= rf_rs2_data_1;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_601) begin
      exe_1_alu_fun <= InstDecoder_1_io_cinfo_alu_fun;
    end
    if (reset) begin
      exe_valid_0 <= 1'h0;
    end else begin
      if (_T_696) begin
        exe_valid_0 <= 1'h0;
      end else begin
        if (_T_601) begin
          exe_valid_0 <= _T_705;
        end
      end
    end
    if (reset) begin
      exe_valid_1 <= 1'h0;
    end else begin
      if (_T_713) begin
        exe_valid_1 <= 1'h0;
      end else begin
        if (_T_601) begin
          exe_valid_1 <= _T_725;
        end
      end
    end
    if (_T_600) begin
      mem_0_rf_wen <= exe_0_rf_wen;
    end
    if (_T_600) begin
      mem_0_wbaddr <= exe_0_wbaddr;
    end
    if (_T_600) begin
      mem_0_mem_en <= exe_0_mem_en;
    end
    if (_T_600) begin
      mem_0_csr_cmd <= exe_0_csr_cmd;
    end
    if (_T_600) begin
      mem_0_illegal <= exe_0_illegal;
    end
    if (_T_600) begin
      mem_0_pc <= exe_0_pc;
    end
    if (_T_600) begin
      mem_0_inst <= exe_0_inst;
    end
    if (_T_600) begin
      mem_0_wb_sel <= exe_0_wb_sel;
    end
    if (_T_600) begin
      mem_0_mem_fcn <= exe_0_mem_fcn;
    end
    if (_T_600) begin
      mem_0_mem_typ <= exe_0_mem_typ;
    end
    if (_T_600) begin
      mem_1_rf_wen <= exe_1_rf_wen;
    end
    if (_T_600) begin
      mem_1_wbaddr <= exe_1_wbaddr;
    end
    if (_T_600) begin
      mem_1_mem_en <= exe_1_mem_en;
    end
    if (_T_600) begin
      mem_1_csr_cmd <= exe_1_csr_cmd;
    end
    if (_T_600) begin
      mem_1_illegal <= exe_1_illegal;
    end
    if (_T_600) begin
      mem_1_pc <= exe_1_pc;
    end
    if (_T_600) begin
      mem_1_inst <= exe_1_inst;
    end
    if (_T_600) begin
      mem_1_wb_sel <= exe_1_wb_sel;
    end
    if (_T_600) begin
      mem_1_mem_fcn <= exe_1_mem_fcn;
    end
    if (_T_600) begin
      mem_1_mem_typ <= exe_1_mem_typ;
    end
    if (reset) begin
      mem_valid_0 <= 1'h0;
    end else begin
      if (_T_815) begin
        mem_valid_0 <= 1'h0;
      end else begin
        if (_T_600) begin
          mem_valid_0 <= exe_valid_0;
        end
      end
    end
    if (reset) begin
      mem_valid_1 <= 1'h0;
    end else begin
      if (_T_822) begin
        mem_valid_1 <= 1'h0;
      end else begin
        if (_T_600) begin
          mem_valid_1 <= _T_828;
        end
      end
    end
    wb_0_rf_wen <= mem_0_rf_wen;
    wb_0_wbaddr <= mem_0_wbaddr;
    wb_1_rf_wen <= mem_1_rf_wen;
    wb_1_wbaddr <= mem_1_wbaddr;
    if (reset) begin
      wb_valid_0 <= 1'h0;
    end else begin
      if (_T_927) begin
        wb_valid_0 <= 1'h0;
      end else begin
        wb_valid_0 <= mem_valid_0;
      end
    end
    if (reset) begin
      wb_valid_1 <= 1'h0;
    end else begin
      if (_T_929) begin
        wb_valid_1 <= 1'h0;
      end else begin
        wb_valid_1 <= mem_valid_1;
      end
    end
    if (_T_866) begin
      wb_wbdata_0 <= io_mem_resp_bits_data;
    end else begin
      if (_T_867) begin
        wb_wbdata_0 <= csr_io_rw_rdata;
      end else begin
        wb_wbdata_0 <= mem_reg_wbdata_0;
      end
    end
    if (_T_885) begin
      wb_wbdata_1 <= io_mem_resp_bits_data;
    end else begin
      if (_T_886) begin
        wb_wbdata_1 <= csr_io_rw_rdata;
      end else begin
        wb_wbdata_1 <= mem_reg_wbdata_1;
      end
    end
    if (_T_600) begin
      mem_reg_wbdata_0 <= exe_wbdata_0;
    end
    if (_T_600) begin
      mem_reg_wbdata_1 <= exe_wbdata_1;
    end
    if (reset) begin
      mem_reg_jpnpc <= 32'h0;
    end else begin
      if (_T_600) begin
        mem_reg_jpnpc <= _T_810;
      end
    end
    if (_T_601) begin
      exe_btb_redirect <= io_front_pred_redirect;
    end
    if (_T_601) begin
      exe_btb_history <= io_front_pred_history;
    end
    if (_T_601) begin
      exe_btb_diff <= io_front_pred_diff;
    end
    if (_T_601) begin
      exe_btb_tgt <= io_front_pred_tgt;
    end
    if (_T_601) begin
      exe_branch <= io_front_branch;
    end
    if (_T_601) begin
      exe_call <= io_front_call;
    end
    if (_T_601) begin
      exe_retn <= io_front_retn;
    end
    if (reset) begin
      _T_759 <= 1'h1;
    end else begin
      if (_T_600) begin
        _T_759 <= 1'h1;
      end else begin
        if (exe_wire_retn) begin
          _T_759 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_767 <= 1'h1;
    end else begin
      if (_T_600) begin
        _T_767 <= 1'h1;
      end else begin
        if (exe_wire_call) begin
          _T_767 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_775 <= 1'h1;
    end else begin
      if (_T_600) begin
        _T_775 <= 1'h1;
      end else begin
        if (exe_bj_valid) begin
          _T_775 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_1127 <= 1'h1;
    end else begin
      if (_T_600) begin
        _T_1127 <= 1'h1;
      end else begin
        if (mispredict) begin
          _T_1127 <= 1'h0;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1198) begin
          $fwrite(32'h80000002,"Core: Cyc= %d PC(%x, %x, %x) [%c%c %c%c %c%c] %c%c %c%c Exe: DASM(%x)\n",io_cyc,io_front_pc_0,exe_0_pc,mem_0_pc,_T_1149,8'h30,8'h20,8'h30,_T_1157,8'h30,_T_1175,8'h30,_T_1179,8'h30,_T_1195); // @[BackEnd.scala 416:11:@8773.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1198) begin
          $fwrite(32'h80000002,"Core: Cyc= %d PC(%x, %x, %x) [%c%c %c%c %c%c] %c%c %c%c Exe: DASM(%x)\n",io_cyc,io_front_pc_1,exe_1_pc,mem_1_pc,_T_1201,8'h31,_T_1205,8'h31,_T_1209,8'h31,_T_1227,8'h31,_T_1179,8'h31,_T_1247); // @[BackEnd.scala 416:11:@8800.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid_0 & _T_1198) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_0_rf_wen,wb_0_wbaddr,regfile_io_wdata_0); // @[BackEnd.scala 435:13:@8806.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid_1 & _T_1198) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_1_rf_wen,wb_1_wbaddr,regfile_io_wdata_1); // @[BackEnd.scala 435:13:@8813.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_front_feedBack_valid & _T_1198) begin
          $fwrite(32'h80000002,"BranchJump: Cyc= %d kill %x pc %x tgt %x actual %x expect %x inst DASM(%x)\n",io_cyc,mispredict,io_front_fb_pc,io_front_feedBack_tgt,io_front_feedBack_redirect,exe_btb_redirect,_T_1257); // @[BackEnd.scala 445:11:@8821.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module fuxi( // @[:@8825.2]
  input         clock, // @[:@8826.4]
  input         reset, // @[:@8827.4]
  input         io_imem_addr_ready, // @[:@8828.4]
  output        io_imem_addr_valid, // @[:@8828.4]
  output [31:0] io_imem_addr_bits, // @[:@8828.4]
  input         io_imem_inst_0_valid, // @[:@8828.4]
  input  [31:0] io_imem_inst_0_bits, // @[:@8828.4]
  input         io_imem_inst_1_valid, // @[:@8828.4]
  input  [31:0] io_imem_inst_1_bits, // @[:@8828.4]
  output        io_dmem_req_valid, // @[:@8828.4]
  output [31:0] io_dmem_req_bits_addr, // @[:@8828.4]
  output [31:0] io_dmem_req_bits_data, // @[:@8828.4]
  output        io_dmem_req_bits_fcn, // @[:@8828.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:@8828.4]
  input         io_dmem_resp_valid, // @[:@8828.4]
  input  [31:0] io_dmem_resp_bits_data // @[:@8828.4]
);
  wire  frontEnd_clock; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_reset; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_cyc; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_mem_addr_ready; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_mem_addr_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_mem_addr_bits; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_mem_inst_0_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_mem_inst_0_bits; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_mem_inst_1_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_mem_inst_1_bits; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_xcpt_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_xcpt_bits; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_kill; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_forward_0; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_forward_1; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_inst_0_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_inst_0_bits; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_inst_1_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_inst_1_bits; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_pc_0; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_pc_1; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_split; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_pred_redirect; // @[Core.scala 37:24:@8830.4]
  wire [9:0] frontEnd_io_back_pred_history; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_pred_diff; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_pred_tgt; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_branch; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_call; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_retn; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_bj_sel_0; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_bj_sel_1; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_ras_pop; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_ras_push_valid; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_ras_push_bits; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_fb_pc; // @[Core.scala 37:24:@8830.4]
  wire [1:0] frontEnd_io_back_fb_type; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_feedBack_redirect; // @[Core.scala 37:24:@8830.4]
  wire [9:0] frontEnd_io_back_feedBack_history; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_feedBack_diff; // @[Core.scala 37:24:@8830.4]
  wire [31:0] frontEnd_io_back_feedBack_tgt; // @[Core.scala 37:24:@8830.4]
  wire  frontEnd_io_back_feedBack_valid; // @[Core.scala 37:24:@8830.4]
  wire  backEnd_clock; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_reset; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_mem_req_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_mem_req_bits_addr; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_mem_req_bits_data; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_mem_req_bits_fcn; // @[Core.scala 38:24:@8833.4]
  wire [2:0] backEnd_io_mem_req_bits_typ; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_mem_resp_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_mem_resp_bits_data; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_cyc; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_xcpt_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_xcpt_bits; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_kill; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_forward_0; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_forward_1; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_inst_0_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_inst_0_bits; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_inst_1_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_inst_1_bits; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_pc_0; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_pc_1; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_split; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_pred_redirect; // @[Core.scala 38:24:@8833.4]
  wire [9:0] backEnd_io_front_pred_history; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_pred_diff; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_pred_tgt; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_branch; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_call; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_retn; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_bj_sel_0; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_bj_sel_1; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_ras_pop; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_ras_push_valid; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_ras_push_bits; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_fb_pc; // @[Core.scala 38:24:@8833.4]
  wire [1:0] backEnd_io_front_fb_type; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_feedBack_redirect; // @[Core.scala 38:24:@8833.4]
  wire [9:0] backEnd_io_front_feedBack_history; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_feedBack_diff; // @[Core.scala 38:24:@8833.4]
  wire [31:0] backEnd_io_front_feedBack_tgt; // @[Core.scala 38:24:@8833.4]
  wire  backEnd_io_front_feedBack_valid; // @[Core.scala 38:24:@8833.4]
  FrontEnd frontEnd ( // @[Core.scala 37:24:@8830.4]
    .clock(frontEnd_clock),
    .reset(frontEnd_reset),
    .io_cyc(frontEnd_io_cyc),
    .io_mem_addr_ready(frontEnd_io_mem_addr_ready),
    .io_mem_addr_valid(frontEnd_io_mem_addr_valid),
    .io_mem_addr_bits(frontEnd_io_mem_addr_bits),
    .io_mem_inst_0_valid(frontEnd_io_mem_inst_0_valid),
    .io_mem_inst_0_bits(frontEnd_io_mem_inst_0_bits),
    .io_mem_inst_1_valid(frontEnd_io_mem_inst_1_valid),
    .io_mem_inst_1_bits(frontEnd_io_mem_inst_1_bits),
    .io_back_xcpt_valid(frontEnd_io_back_xcpt_valid),
    .io_back_xcpt_bits(frontEnd_io_back_xcpt_bits),
    .io_back_kill(frontEnd_io_back_kill),
    .io_back_forward_0(frontEnd_io_back_forward_0),
    .io_back_forward_1(frontEnd_io_back_forward_1),
    .io_back_inst_0_valid(frontEnd_io_back_inst_0_valid),
    .io_back_inst_0_bits(frontEnd_io_back_inst_0_bits),
    .io_back_inst_1_valid(frontEnd_io_back_inst_1_valid),
    .io_back_inst_1_bits(frontEnd_io_back_inst_1_bits),
    .io_back_pc_0(frontEnd_io_back_pc_0),
    .io_back_pc_1(frontEnd_io_back_pc_1),
    .io_back_split(frontEnd_io_back_split),
    .io_back_pred_redirect(frontEnd_io_back_pred_redirect),
    .io_back_pred_history(frontEnd_io_back_pred_history),
    .io_back_pred_diff(frontEnd_io_back_pred_diff),
    .io_back_pred_tgt(frontEnd_io_back_pred_tgt),
    .io_back_branch(frontEnd_io_back_branch),
    .io_back_call(frontEnd_io_back_call),
    .io_back_retn(frontEnd_io_back_retn),
    .io_back_bj_sel_0(frontEnd_io_back_bj_sel_0),
    .io_back_bj_sel_1(frontEnd_io_back_bj_sel_1),
    .io_back_ras_pop(frontEnd_io_back_ras_pop),
    .io_back_ras_push_valid(frontEnd_io_back_ras_push_valid),
    .io_back_ras_push_bits(frontEnd_io_back_ras_push_bits),
    .io_back_fb_pc(frontEnd_io_back_fb_pc),
    .io_back_fb_type(frontEnd_io_back_fb_type),
    .io_back_feedBack_redirect(frontEnd_io_back_feedBack_redirect),
    .io_back_feedBack_history(frontEnd_io_back_feedBack_history),
    .io_back_feedBack_diff(frontEnd_io_back_feedBack_diff),
    .io_back_feedBack_tgt(frontEnd_io_back_feedBack_tgt),
    .io_back_feedBack_valid(frontEnd_io_back_feedBack_valid)
  );
  BackEnd backEnd ( // @[Core.scala 38:24:@8833.4]
    .clock(backEnd_clock),
    .reset(backEnd_reset),
    .io_mem_req_valid(backEnd_io_mem_req_valid),
    .io_mem_req_bits_addr(backEnd_io_mem_req_bits_addr),
    .io_mem_req_bits_data(backEnd_io_mem_req_bits_data),
    .io_mem_req_bits_fcn(backEnd_io_mem_req_bits_fcn),
    .io_mem_req_bits_typ(backEnd_io_mem_req_bits_typ),
    .io_mem_resp_valid(backEnd_io_mem_resp_valid),
    .io_mem_resp_bits_data(backEnd_io_mem_resp_bits_data),
    .io_cyc(backEnd_io_cyc),
    .io_front_xcpt_valid(backEnd_io_front_xcpt_valid),
    .io_front_xcpt_bits(backEnd_io_front_xcpt_bits),
    .io_front_kill(backEnd_io_front_kill),
    .io_front_forward_0(backEnd_io_front_forward_0),
    .io_front_forward_1(backEnd_io_front_forward_1),
    .io_front_inst_0_valid(backEnd_io_front_inst_0_valid),
    .io_front_inst_0_bits(backEnd_io_front_inst_0_bits),
    .io_front_inst_1_valid(backEnd_io_front_inst_1_valid),
    .io_front_inst_1_bits(backEnd_io_front_inst_1_bits),
    .io_front_pc_0(backEnd_io_front_pc_0),
    .io_front_pc_1(backEnd_io_front_pc_1),
    .io_front_split(backEnd_io_front_split),
    .io_front_pred_redirect(backEnd_io_front_pred_redirect),
    .io_front_pred_history(backEnd_io_front_pred_history),
    .io_front_pred_diff(backEnd_io_front_pred_diff),
    .io_front_pred_tgt(backEnd_io_front_pred_tgt),
    .io_front_branch(backEnd_io_front_branch),
    .io_front_call(backEnd_io_front_call),
    .io_front_retn(backEnd_io_front_retn),
    .io_front_bj_sel_0(backEnd_io_front_bj_sel_0),
    .io_front_bj_sel_1(backEnd_io_front_bj_sel_1),
    .io_front_ras_pop(backEnd_io_front_ras_pop),
    .io_front_ras_push_valid(backEnd_io_front_ras_push_valid),
    .io_front_ras_push_bits(backEnd_io_front_ras_push_bits),
    .io_front_fb_pc(backEnd_io_front_fb_pc),
    .io_front_fb_type(backEnd_io_front_fb_type),
    .io_front_feedBack_redirect(backEnd_io_front_feedBack_redirect),
    .io_front_feedBack_history(backEnd_io_front_feedBack_history),
    .io_front_feedBack_diff(backEnd_io_front_feedBack_diff),
    .io_front_feedBack_tgt(backEnd_io_front_feedBack_tgt),
    .io_front_feedBack_valid(backEnd_io_front_feedBack_valid)
  );
  assign io_imem_addr_valid = frontEnd_io_mem_addr_valid; // @[Core.scala 39:19:@8841.4]
  assign io_imem_addr_bits = frontEnd_io_mem_addr_bits; // @[Core.scala 39:19:@8840.4]
  assign io_dmem_req_valid = backEnd_io_mem_req_valid; // @[Core.scala 40:19:@8849.4]
  assign io_dmem_req_bits_addr = backEnd_io_mem_req_bits_addr; // @[Core.scala 40:19:@8848.4]
  assign io_dmem_req_bits_data = backEnd_io_mem_req_bits_data; // @[Core.scala 40:19:@8847.4]
  assign io_dmem_req_bits_fcn = backEnd_io_mem_req_bits_fcn; // @[Core.scala 40:19:@8846.4]
  assign io_dmem_req_bits_typ = backEnd_io_mem_req_bits_typ; // @[Core.scala 40:19:@8845.4]
  assign frontEnd_clock = clock; // @[:@8831.4]
  assign frontEnd_reset = reset; // @[:@8832.4]
  assign frontEnd_io_cyc = backEnd_io_cyc; // @[Core.scala 43:20:@8882.4]
  assign frontEnd_io_mem_addr_ready = io_imem_addr_ready; // @[Core.scala 39:19:@8842.4]
  assign frontEnd_io_mem_inst_0_valid = io_imem_inst_0_valid; // @[Core.scala 39:19:@8837.4]
  assign frontEnd_io_mem_inst_0_bits = io_imem_inst_0_bits; // @[Core.scala 39:19:@8836.4]
  assign frontEnd_io_mem_inst_1_valid = io_imem_inst_1_valid; // @[Core.scala 39:19:@8839.4]
  assign frontEnd_io_mem_inst_1_bits = io_imem_inst_1_bits; // @[Core.scala 39:19:@8838.4]
  assign frontEnd_io_back_xcpt_valid = backEnd_io_front_xcpt_valid; // @[Core.scala 42:20:@8881.4]
  assign frontEnd_io_back_xcpt_bits = backEnd_io_front_xcpt_bits; // @[Core.scala 42:20:@8880.4]
  assign frontEnd_io_back_kill = backEnd_io_front_kill; // @[Core.scala 42:20:@8879.4]
  assign frontEnd_io_back_forward_0 = backEnd_io_front_forward_0; // @[Core.scala 42:20:@8877.4]
  assign frontEnd_io_back_forward_1 = backEnd_io_front_forward_1; // @[Core.scala 42:20:@8878.4]
  assign frontEnd_io_back_ras_pop = backEnd_io_front_ras_pop; // @[Core.scala 42:20:@8860.4]
  assign frontEnd_io_back_ras_push_valid = backEnd_io_front_ras_push_valid; // @[Core.scala 42:20:@8859.4]
  assign frontEnd_io_back_ras_push_bits = backEnd_io_front_ras_push_bits; // @[Core.scala 42:20:@8858.4]
  assign frontEnd_io_back_fb_pc = backEnd_io_front_fb_pc; // @[Core.scala 42:20:@8857.4]
  assign frontEnd_io_back_fb_type = backEnd_io_front_fb_type; // @[Core.scala 42:20:@8856.4]
  assign frontEnd_io_back_feedBack_redirect = backEnd_io_front_feedBack_redirect; // @[Core.scala 42:20:@8855.4]
  assign frontEnd_io_back_feedBack_history = backEnd_io_front_feedBack_history; // @[Core.scala 42:20:@8854.4]
  assign frontEnd_io_back_feedBack_diff = backEnd_io_front_feedBack_diff; // @[Core.scala 42:20:@8853.4]
  assign frontEnd_io_back_feedBack_tgt = backEnd_io_front_feedBack_tgt; // @[Core.scala 42:20:@8852.4]
  assign frontEnd_io_back_feedBack_valid = backEnd_io_front_feedBack_valid; // @[Core.scala 42:20:@8851.4]
  assign backEnd_clock = clock; // @[:@8834.4]
  assign backEnd_reset = reset; // @[:@8835.4]
  assign backEnd_io_mem_resp_valid = io_dmem_resp_valid; // @[Core.scala 40:19:@8844.4]
  assign backEnd_io_mem_resp_bits_data = io_dmem_resp_bits_data; // @[Core.scala 40:19:@8843.4]
  assign backEnd_io_front_inst_0_valid = frontEnd_io_back_inst_0_valid; // @[Core.scala 42:20:@8874.4]
  assign backEnd_io_front_inst_0_bits = frontEnd_io_back_inst_0_bits; // @[Core.scala 42:20:@8873.4]
  assign backEnd_io_front_inst_1_valid = frontEnd_io_back_inst_1_valid; // @[Core.scala 42:20:@8876.4]
  assign backEnd_io_front_inst_1_bits = frontEnd_io_back_inst_1_bits; // @[Core.scala 42:20:@8875.4]
  assign backEnd_io_front_pc_0 = frontEnd_io_back_pc_0; // @[Core.scala 42:20:@8871.4]
  assign backEnd_io_front_pc_1 = frontEnd_io_back_pc_1; // @[Core.scala 42:20:@8872.4]
  assign backEnd_io_front_split = frontEnd_io_back_split; // @[Core.scala 42:20:@8870.4]
  assign backEnd_io_front_pred_redirect = frontEnd_io_back_pred_redirect; // @[Core.scala 42:20:@8869.4]
  assign backEnd_io_front_pred_history = frontEnd_io_back_pred_history; // @[Core.scala 42:20:@8868.4]
  assign backEnd_io_front_pred_diff = frontEnd_io_back_pred_diff; // @[Core.scala 42:20:@8867.4]
  assign backEnd_io_front_pred_tgt = frontEnd_io_back_pred_tgt; // @[Core.scala 42:20:@8866.4]
  assign backEnd_io_front_branch = frontEnd_io_back_branch; // @[Core.scala 42:20:@8865.4]
  assign backEnd_io_front_call = frontEnd_io_back_call; // @[Core.scala 42:20:@8864.4]
  assign backEnd_io_front_retn = frontEnd_io_back_retn; // @[Core.scala 42:20:@8863.4]
  assign backEnd_io_front_bj_sel_0 = frontEnd_io_back_bj_sel_0; // @[Core.scala 42:20:@8861.4]
  assign backEnd_io_front_bj_sel_1 = frontEnd_io_back_bj_sel_1; // @[Core.scala 42:20:@8862.4]
endmodule