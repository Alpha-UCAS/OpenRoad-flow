module RAS( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input         io_push_valid, // @[:@6.4]
  input  [31:0] io_push_bits, // @[:@6.4]
  input         io_pop, // @[:@6.4]
  output [31:0] io_peek // @[:@6.4]
);
  reg [31:0] stack_0; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_0;
  reg [31:0] stack_1; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_1;
  reg [31:0] stack_2; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_2;
  reg [31:0] stack_3; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_3;
  reg [31:0] stack_4; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_4;
  reg [31:0] stack_5; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_5;
  reg [31:0] stack_6; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_6;
  reg [31:0] stack_7; // @[RAS.scala 15:18:@8.4]
  reg [31:0] _RAND_7;
  reg [2:0] pos; // @[RAS.scala 16:22:@9.4]
  reg [31:0] _RAND_8;
  reg [3:0] count; // @[RAS.scala 17:22:@10.4]
  reg [31:0] _RAND_9;
  wire  empty; // @[RAS.scala 18:27:@11.4]
  wire [3:0] _T_37; // @[RAS.scala 20:18:@13.4]
  wire [2:0] nextPos; // @[RAS.scala 20:18:@14.4]
  wire [31:0] _GEN_1; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_2; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_3; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_4; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_5; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_6; // @[RAS.scala 21:11:@16.4]
  wire [31:0] _GEN_8; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_9; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_10; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_11; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_12; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_13; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_14; // @[RAS.scala 25:18:@19.8]
  wire [31:0] _GEN_15; // @[RAS.scala 25:18:@19.8]
  wire  _T_42; // @[RAS.scala 27:19:@22.8]
  wire [4:0] _T_44; // @[RAS.scala 27:48:@24.10]
  wire [3:0] _T_45; // @[RAS.scala 27:48:@25.10]
  wire [3:0] _GEN_16; // @[RAS.scala 27:31:@23.8]
  wire [31:0] _GEN_17; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_18; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_19; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_20; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_21; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_22; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_23; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_24; // @[RAS.scala 28:22:@28.8]
  wire [31:0] _GEN_25; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_26; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_27; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_28; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_29; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_30; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_31; // @[RAS.scala 24:18:@18.6]
  wire [31:0] _GEN_32; // @[RAS.scala 24:18:@18.6]
  wire [3:0] _GEN_33; // @[RAS.scala 24:18:@18.6]
  wire [2:0] _GEN_34; // @[RAS.scala 24:18:@18.6]
  wire  _T_48; // @[RAS.scala 31:23:@33.6]
  wire  _T_49; // @[RAS.scala 31:21:@34.6]
  wire [4:0] _T_51; // @[RAS.scala 32:20:@36.8]
  wire [4:0] _T_52; // @[RAS.scala 32:20:@37.8]
  wire [3:0] _T_53; // @[RAS.scala 32:20:@38.8]
  wire [3:0] _T_55; // @[RAS.scala 33:16:@40.8]
  wire [3:0] _T_56; // @[RAS.scala 33:16:@41.8]
  wire [2:0] _T_57; // @[RAS.scala 33:16:@42.8]
  wire [3:0] _GEN_35; // @[RAS.scala 31:31:@35.6]
  wire [2:0] _GEN_36; // @[RAS.scala 31:31:@35.6]
  wire [3:0] _GEN_45; // @[RAS.scala 23:23:@17.4]
  wire [2:0] _GEN_46; // @[RAS.scala 23:23:@17.4]
  assign empty = count == 4'h0; // @[RAS.scala 18:27:@11.4]
  assign _T_37 = pos + 3'h1; // @[RAS.scala 20:18:@13.4]
  assign nextPos = pos + 3'h1; // @[RAS.scala 20:18:@14.4]
  assign _GEN_1 = 3'h1 == pos ? stack_1 : stack_0; // @[RAS.scala 21:11:@16.4]
  assign _GEN_2 = 3'h2 == pos ? stack_2 : _GEN_1; // @[RAS.scala 21:11:@16.4]
  assign _GEN_3 = 3'h3 == pos ? stack_3 : _GEN_2; // @[RAS.scala 21:11:@16.4]
  assign _GEN_4 = 3'h4 == pos ? stack_4 : _GEN_3; // @[RAS.scala 21:11:@16.4]
  assign _GEN_5 = 3'h5 == pos ? stack_5 : _GEN_4; // @[RAS.scala 21:11:@16.4]
  assign _GEN_6 = 3'h6 == pos ? stack_6 : _GEN_5; // @[RAS.scala 21:11:@16.4]
  assign _GEN_8 = 3'h0 == pos ? io_push_bits : stack_0; // @[RAS.scala 25:18:@19.8]
  assign _GEN_9 = 3'h1 == pos ? io_push_bits : stack_1; // @[RAS.scala 25:18:@19.8]
  assign _GEN_10 = 3'h2 == pos ? io_push_bits : stack_2; // @[RAS.scala 25:18:@19.8]
  assign _GEN_11 = 3'h3 == pos ? io_push_bits : stack_3; // @[RAS.scala 25:18:@19.8]
  assign _GEN_12 = 3'h4 == pos ? io_push_bits : stack_4; // @[RAS.scala 25:18:@19.8]
  assign _GEN_13 = 3'h5 == pos ? io_push_bits : stack_5; // @[RAS.scala 25:18:@19.8]
  assign _GEN_14 = 3'h6 == pos ? io_push_bits : stack_6; // @[RAS.scala 25:18:@19.8]
  assign _GEN_15 = 3'h7 == pos ? io_push_bits : stack_7; // @[RAS.scala 25:18:@19.8]
  assign _T_42 = count != 4'h8; // @[RAS.scala 27:19:@22.8]
  assign _T_44 = count + 4'h1; // @[RAS.scala 27:48:@24.10]
  assign _T_45 = count + 4'h1; // @[RAS.scala 27:48:@25.10]
  assign _GEN_16 = _T_42 ? _T_45 : count; // @[RAS.scala 27:31:@23.8]
  assign _GEN_17 = 3'h0 == nextPos ? io_push_bits : stack_0; // @[RAS.scala 28:22:@28.8]
  assign _GEN_18 = 3'h1 == nextPos ? io_push_bits : stack_1; // @[RAS.scala 28:22:@28.8]
  assign _GEN_19 = 3'h2 == nextPos ? io_push_bits : stack_2; // @[RAS.scala 28:22:@28.8]
  assign _GEN_20 = 3'h3 == nextPos ? io_push_bits : stack_3; // @[RAS.scala 28:22:@28.8]
  assign _GEN_21 = 3'h4 == nextPos ? io_push_bits : stack_4; // @[RAS.scala 28:22:@28.8]
  assign _GEN_22 = 3'h5 == nextPos ? io_push_bits : stack_5; // @[RAS.scala 28:22:@28.8]
  assign _GEN_23 = 3'h6 == nextPos ? io_push_bits : stack_6; // @[RAS.scala 28:22:@28.8]
  assign _GEN_24 = 3'h7 == nextPos ? io_push_bits : stack_7; // @[RAS.scala 28:22:@28.8]
  assign _GEN_25 = io_pop ? _GEN_8 : _GEN_17; // @[RAS.scala 24:18:@18.6]
  assign _GEN_26 = io_pop ? _GEN_9 : _GEN_18; // @[RAS.scala 24:18:@18.6]
  assign _GEN_27 = io_pop ? _GEN_10 : _GEN_19; // @[RAS.scala 24:18:@18.6]
  assign _GEN_28 = io_pop ? _GEN_11 : _GEN_20; // @[RAS.scala 24:18:@18.6]
  assign _GEN_29 = io_pop ? _GEN_12 : _GEN_21; // @[RAS.scala 24:18:@18.6]
  assign _GEN_30 = io_pop ? _GEN_13 : _GEN_22; // @[RAS.scala 24:18:@18.6]
  assign _GEN_31 = io_pop ? _GEN_14 : _GEN_23; // @[RAS.scala 24:18:@18.6]
  assign _GEN_32 = io_pop ? _GEN_15 : _GEN_24; // @[RAS.scala 24:18:@18.6]
  assign _GEN_33 = io_pop ? count : _GEN_16; // @[RAS.scala 24:18:@18.6]
  assign _GEN_34 = io_pop ? pos : nextPos; // @[RAS.scala 24:18:@18.6]
  assign _T_48 = empty == 1'h0; // @[RAS.scala 31:23:@33.6]
  assign _T_49 = io_pop & _T_48; // @[RAS.scala 31:21:@34.6]
  assign _T_51 = count - 4'h1; // @[RAS.scala 32:20:@36.8]
  assign _T_52 = $unsigned(_T_51); // @[RAS.scala 32:20:@37.8]
  assign _T_53 = _T_52[3:0]; // @[RAS.scala 32:20:@38.8]
  assign _T_55 = pos - 3'h1; // @[RAS.scala 33:16:@40.8]
  assign _T_56 = $unsigned(_T_55); // @[RAS.scala 33:16:@41.8]
  assign _T_57 = _T_56[2:0]; // @[RAS.scala 33:16:@42.8]
  assign _GEN_35 = _T_49 ? _T_53 : count; // @[RAS.scala 31:31:@35.6]
  assign _GEN_36 = _T_49 ? _T_57 : pos; // @[RAS.scala 31:31:@35.6]
  assign _GEN_45 = io_push_valid ? _GEN_33 : _GEN_35; // @[RAS.scala 23:23:@17.4]
  assign _GEN_46 = io_push_valid ? _GEN_34 : _GEN_36; // @[RAS.scala 23:23:@17.4]
  assign io_peek = 3'h7 == pos ? stack_7 : _GEN_6; // @[RAS.scala 21:11:@16.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  stack_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  stack_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  stack_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  stack_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  stack_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  stack_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  stack_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  stack_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  pos = _RAND_8[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  count = _RAND_9[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h0 == pos) begin
          stack_0 <= io_push_bits;
        end
      end else begin
        if (3'h0 == nextPos) begin
          stack_0 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h1 == pos) begin
          stack_1 <= io_push_bits;
        end
      end else begin
        if (3'h1 == nextPos) begin
          stack_1 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h2 == pos) begin
          stack_2 <= io_push_bits;
        end
      end else begin
        if (3'h2 == nextPos) begin
          stack_2 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h3 == pos) begin
          stack_3 <= io_push_bits;
        end
      end else begin
        if (3'h3 == nextPos) begin
          stack_3 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h4 == pos) begin
          stack_4 <= io_push_bits;
        end
      end else begin
        if (3'h4 == nextPos) begin
          stack_4 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h5 == pos) begin
          stack_5 <= io_push_bits;
        end
      end else begin
        if (3'h5 == nextPos) begin
          stack_5 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h6 == pos) begin
          stack_6 <= io_push_bits;
        end
      end else begin
        if (3'h6 == nextPos) begin
          stack_6 <= io_push_bits;
        end
      end
    end
    if (io_push_valid) begin
      if (io_pop) begin
        if (3'h7 == pos) begin
          stack_7 <= io_push_bits;
        end
      end else begin
        if (3'h7 == nextPos) begin
          stack_7 <= io_push_bits;
        end
      end
    end
    if (reset) begin
      pos <= 3'h0;
    end else begin
      if (io_push_valid) begin
        if (!(io_pop)) begin
          pos <= nextPos;
        end
      end else begin
        if (_T_49) begin
          pos <= _T_57;
        end
      end
    end
    if (reset) begin
      count <= 4'h0;
    end else begin
      if (io_push_valid) begin
        if (!(io_pop)) begin
          if (_T_42) begin
            count <= _T_45;
          end
        end
      end else begin
        if (_T_49) begin
          count <= _T_53;
        end
      end
    end
  end
endmodule
module BTB( // @[:@46.2]
  input         clock, // @[:@47.4]
  input         reset, // @[:@48.4]
  input  [31:0] io_if_pc, // @[:@49.4]
  output        io_predict_redirect, // @[:@49.4]
  output [9:0]  io_predict_history, // @[:@49.4]
  output        io_predict_diff, // @[:@49.4]
  output [31:0] io_predict_tgt, // @[:@49.4]
  input         io_branch, // @[:@49.4]
  input         io_forward, // @[:@49.4]
  input         io_ras_pop, // @[:@49.4]
  input         io_ras_push_valid, // @[:@49.4]
  input  [31:0] io_ras_push_bits, // @[:@49.4]
  input  [31:0] io_fb_pc, // @[:@49.4]
  input         io_fb_miss, // @[:@49.4]
  input  [1:0]  io_fb_type, // @[:@49.4]
  input         io_feedBack_redirect, // @[:@49.4]
  input  [9:0]  io_feedBack_history, // @[:@49.4]
  input         io_feedBack_diff, // @[:@49.4]
  input  [31:0] io_feedBack_tgt, // @[:@49.4]
  input         io_feedBack_valid, // @[:@49.4]
  input  [31:0] io_cyc // @[:@49.4]
);
  reg [1:0] bht [0:1023]; // @[BTB.scala 67:16:@52.4]
  reg [31:0] _RAND_0;
  wire [1:0] bht__T_1188_data; // @[BTB.scala 67:16:@52.4]
  wire [9:0] bht__T_1188_addr; // @[BTB.scala 67:16:@52.4]
  wire [1:0] bht__T_1774_data; // @[BTB.scala 67:16:@52.4]
  wire [9:0] bht__T_1774_addr; // @[BTB.scala 67:16:@52.4]
  wire [1:0] bht__T_2148_data; // @[BTB.scala 67:16:@52.4]
  wire [9:0] bht__T_2148_addr; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2148_mask; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2148_en; // @[BTB.scala 67:16:@52.4]
  wire [1:0] bht__T_2166_data; // @[BTB.scala 67:16:@52.4]
  wire [9:0] bht__T_2166_addr; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2166_mask; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2166_en; // @[BTB.scala 67:16:@52.4]
  wire [1:0] bht__T_2177_data; // @[BTB.scala 67:16:@52.4]
  wire [9:0] bht__T_2177_addr; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2177_mask; // @[BTB.scala 67:16:@52.4]
  wire  bht__T_2177_en; // @[BTB.scala 67:16:@52.4]
  reg  arb [0:1023]; // @[BTB.scala 68:16:@53.4]
  reg [31:0] _RAND_1;
  wire  arb__T_1187_data; // @[BTB.scala 68:16:@53.4]
  wire [9:0] arb__T_1187_addr; // @[BTB.scala 68:16:@53.4]
  wire  arb_gshare_sel_data; // @[BTB.scala 68:16:@53.4]
  wire [9:0] arb_gshare_sel_addr; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2185_data; // @[BTB.scala 68:16:@53.4]
  wire [9:0] arb__T_2185_addr; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2185_mask; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2185_en; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2187_data; // @[BTB.scala 68:16:@53.4]
  wire [9:0] arb__T_2187_addr; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2187_mask; // @[BTB.scala 68:16:@53.4]
  wire  arb__T_2187_en; // @[BTB.scala 68:16:@53.4]
  wire  RAS_clock; // @[BTB.scala 69:19:@54.4]
  wire  RAS_reset; // @[BTB.scala 69:19:@54.4]
  wire  RAS_io_push_valid; // @[BTB.scala 69:19:@54.4]
  wire [31:0] RAS_io_push_bits; // @[BTB.scala 69:19:@54.4]
  wire  RAS_io_pop; // @[BTB.scala 69:19:@54.4]
  wire [31:0] RAS_io_peek; // @[BTB.scala 69:19:@54.4]
  reg [9:0] gb_history; // @[BTB.scala 66:27:@51.4]
  reg [31:0] _RAND_2;
  reg  btb_valid_0; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_3;
  reg  btb_valid_1; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_4;
  reg  btb_valid_2; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_5;
  reg  btb_valid_3; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_6;
  reg  btb_valid_4; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_7;
  reg  btb_valid_5; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_8;
  reg  btb_valid_6; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_9;
  reg  btb_valid_7; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_10;
  reg  btb_valid_8; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_11;
  reg  btb_valid_9; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_12;
  reg  btb_valid_10; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_13;
  reg  btb_valid_11; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_14;
  reg  btb_valid_12; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_15;
  reg  btb_valid_13; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_16;
  reg  btb_valid_14; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_17;
  reg  btb_valid_15; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_18;
  reg  btb_valid_16; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_19;
  reg  btb_valid_17; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_20;
  reg  btb_valid_18; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_21;
  reg  btb_valid_19; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_22;
  reg  btb_valid_20; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_23;
  reg  btb_valid_21; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_24;
  reg  btb_valid_22; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_25;
  reg  btb_valid_23; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_26;
  reg  btb_valid_24; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_27;
  reg  btb_valid_25; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_28;
  reg  btb_valid_26; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_29;
  reg  btb_valid_27; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_30;
  reg  btb_valid_28; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_31;
  reg  btb_valid_29; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_32;
  reg  btb_valid_30; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_33;
  reg  btb_valid_31; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_34;
  reg  btb_valid_32; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_35;
  reg  btb_valid_33; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_36;
  reg  btb_valid_34; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_37;
  reg  btb_valid_35; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_38;
  reg  btb_valid_36; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_39;
  reg  btb_valid_37; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_40;
  reg  btb_valid_38; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_41;
  reg  btb_valid_39; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_42;
  reg  btb_valid_40; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_43;
  reg  btb_valid_41; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_44;
  reg  btb_valid_42; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_45;
  reg  btb_valid_43; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_46;
  reg  btb_valid_44; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_47;
  reg  btb_valid_45; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_48;
  reg  btb_valid_46; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_49;
  reg  btb_valid_47; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_50;
  reg  btb_valid_48; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_51;
  reg  btb_valid_49; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_52;
  reg  btb_valid_50; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_53;
  reg  btb_valid_51; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_54;
  reg  btb_valid_52; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_55;
  reg  btb_valid_53; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_56;
  reg  btb_valid_54; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_57;
  reg  btb_valid_55; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_58;
  reg  btb_valid_56; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_59;
  reg  btb_valid_57; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_60;
  reg  btb_valid_58; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_61;
  reg  btb_valid_59; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_62;
  reg  btb_valid_60; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_63;
  reg  btb_valid_61; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_64;
  reg  btb_valid_62; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_65;
  reg  btb_valid_63; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_66;
  reg [31:0] btb_pc_0; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_67;
  reg [31:0] btb_pc_1; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_68;
  reg [31:0] btb_pc_2; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_69;
  reg [31:0] btb_pc_3; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_70;
  reg [31:0] btb_pc_4; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_71;
  reg [31:0] btb_pc_5; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_72;
  reg [31:0] btb_pc_6; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_73;
  reg [31:0] btb_pc_7; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_74;
  reg [31:0] btb_pc_8; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_75;
  reg [31:0] btb_pc_9; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_76;
  reg [31:0] btb_pc_10; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_77;
  reg [31:0] btb_pc_11; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_78;
  reg [31:0] btb_pc_12; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_79;
  reg [31:0] btb_pc_13; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_80;
  reg [31:0] btb_pc_14; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_81;
  reg [31:0] btb_pc_15; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_82;
  reg [31:0] btb_pc_16; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_83;
  reg [31:0] btb_pc_17; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_84;
  reg [31:0] btb_pc_18; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_85;
  reg [31:0] btb_pc_19; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_86;
  reg [31:0] btb_pc_20; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_87;
  reg [31:0] btb_pc_21; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_88;
  reg [31:0] btb_pc_22; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_89;
  reg [31:0] btb_pc_23; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_90;
  reg [31:0] btb_pc_24; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_91;
  reg [31:0] btb_pc_25; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_92;
  reg [31:0] btb_pc_26; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_93;
  reg [31:0] btb_pc_27; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_94;
  reg [31:0] btb_pc_28; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_95;
  reg [31:0] btb_pc_29; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_96;
  reg [31:0] btb_pc_30; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_97;
  reg [31:0] btb_pc_31; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_98;
  reg [31:0] btb_pc_32; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_99;
  reg [31:0] btb_pc_33; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_100;
  reg [31:0] btb_pc_34; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_101;
  reg [31:0] btb_pc_35; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_102;
  reg [31:0] btb_pc_36; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_103;
  reg [31:0] btb_pc_37; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_104;
  reg [31:0] btb_pc_38; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_105;
  reg [31:0] btb_pc_39; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_106;
  reg [31:0] btb_pc_40; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_107;
  reg [31:0] btb_pc_41; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_108;
  reg [31:0] btb_pc_42; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_109;
  reg [31:0] btb_pc_43; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_110;
  reg [31:0] btb_pc_44; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_111;
  reg [31:0] btb_pc_45; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_112;
  reg [31:0] btb_pc_46; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_113;
  reg [31:0] btb_pc_47; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_114;
  reg [31:0] btb_pc_48; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_115;
  reg [31:0] btb_pc_49; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_116;
  reg [31:0] btb_pc_50; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_117;
  reg [31:0] btb_pc_51; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_118;
  reg [31:0] btb_pc_52; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_119;
  reg [31:0] btb_pc_53; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_120;
  reg [31:0] btb_pc_54; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_121;
  reg [31:0] btb_pc_55; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_122;
  reg [31:0] btb_pc_56; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_123;
  reg [31:0] btb_pc_57; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_124;
  reg [31:0] btb_pc_58; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_125;
  reg [31:0] btb_pc_59; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_126;
  reg [31:0] btb_pc_60; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_127;
  reg [31:0] btb_pc_61; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_128;
  reg [31:0] btb_pc_62; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_129;
  reg [31:0] btb_pc_63; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_130;
  reg [31:0] btb_tgt_0; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_131;
  reg [31:0] btb_tgt_1; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_132;
  reg [31:0] btb_tgt_2; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_133;
  reg [31:0] btb_tgt_3; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_134;
  reg [31:0] btb_tgt_4; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_135;
  reg [31:0] btb_tgt_5; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_136;
  reg [31:0] btb_tgt_6; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_137;
  reg [31:0] btb_tgt_7; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_138;
  reg [31:0] btb_tgt_8; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_139;
  reg [31:0] btb_tgt_9; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_140;
  reg [31:0] btb_tgt_10; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_141;
  reg [31:0] btb_tgt_11; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_142;
  reg [31:0] btb_tgt_12; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_143;
  reg [31:0] btb_tgt_13; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_144;
  reg [31:0] btb_tgt_14; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_145;
  reg [31:0] btb_tgt_15; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_146;
  reg [31:0] btb_tgt_16; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_147;
  reg [31:0] btb_tgt_17; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_148;
  reg [31:0] btb_tgt_18; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_149;
  reg [31:0] btb_tgt_19; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_150;
  reg [31:0] btb_tgt_20; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_151;
  reg [31:0] btb_tgt_21; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_152;
  reg [31:0] btb_tgt_22; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_153;
  reg [31:0] btb_tgt_23; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_154;
  reg [31:0] btb_tgt_24; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_155;
  reg [31:0] btb_tgt_25; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_156;
  reg [31:0] btb_tgt_26; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_157;
  reg [31:0] btb_tgt_27; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_158;
  reg [31:0] btb_tgt_28; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_159;
  reg [31:0] btb_tgt_29; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_160;
  reg [31:0] btb_tgt_30; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_161;
  reg [31:0] btb_tgt_31; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_162;
  reg [31:0] btb_tgt_32; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_163;
  reg [31:0] btb_tgt_33; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_164;
  reg [31:0] btb_tgt_34; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_165;
  reg [31:0] btb_tgt_35; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_166;
  reg [31:0] btb_tgt_36; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_167;
  reg [31:0] btb_tgt_37; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_168;
  reg [31:0] btb_tgt_38; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_169;
  reg [31:0] btb_tgt_39; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_170;
  reg [31:0] btb_tgt_40; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_171;
  reg [31:0] btb_tgt_41; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_172;
  reg [31:0] btb_tgt_42; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_173;
  reg [31:0] btb_tgt_43; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_174;
  reg [31:0] btb_tgt_44; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_175;
  reg [31:0] btb_tgt_45; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_176;
  reg [31:0] btb_tgt_46; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_177;
  reg [31:0] btb_tgt_47; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_178;
  reg [31:0] btb_tgt_48; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_179;
  reg [31:0] btb_tgt_49; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_180;
  reg [31:0] btb_tgt_50; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_181;
  reg [31:0] btb_tgt_51; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_182;
  reg [31:0] btb_tgt_52; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_183;
  reg [31:0] btb_tgt_53; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_184;
  reg [31:0] btb_tgt_54; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_185;
  reg [31:0] btb_tgt_55; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_186;
  reg [31:0] btb_tgt_56; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_187;
  reg [31:0] btb_tgt_57; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_188;
  reg [31:0] btb_tgt_58; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_189;
  reg [31:0] btb_tgt_59; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_190;
  reg [31:0] btb_tgt_60; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_191;
  reg [31:0] btb_tgt_61; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_192;
  reg [31:0] btb_tgt_62; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_193;
  reg [31:0] btb_tgt_63; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_194;
  reg [1:0] btb_bj_type_0; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_195;
  reg [1:0] btb_bj_type_1; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_196;
  reg [1:0] btb_bj_type_2; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_197;
  reg [1:0] btb_bj_type_3; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_198;
  reg [1:0] btb_bj_type_4; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_199;
  reg [1:0] btb_bj_type_5; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_200;
  reg [1:0] btb_bj_type_6; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_201;
  reg [1:0] btb_bj_type_7; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_202;
  reg [1:0] btb_bj_type_8; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_203;
  reg [1:0] btb_bj_type_9; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_204;
  reg [1:0] btb_bj_type_10; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_205;
  reg [1:0] btb_bj_type_11; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_206;
  reg [1:0] btb_bj_type_12; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_207;
  reg [1:0] btb_bj_type_13; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_208;
  reg [1:0] btb_bj_type_14; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_209;
  reg [1:0] btb_bj_type_15; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_210;
  reg [1:0] btb_bj_type_16; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_211;
  reg [1:0] btb_bj_type_17; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_212;
  reg [1:0] btb_bj_type_18; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_213;
  reg [1:0] btb_bj_type_19; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_214;
  reg [1:0] btb_bj_type_20; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_215;
  reg [1:0] btb_bj_type_21; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_216;
  reg [1:0] btb_bj_type_22; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_217;
  reg [1:0] btb_bj_type_23; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_218;
  reg [1:0] btb_bj_type_24; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_219;
  reg [1:0] btb_bj_type_25; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_220;
  reg [1:0] btb_bj_type_26; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_221;
  reg [1:0] btb_bj_type_27; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_222;
  reg [1:0] btb_bj_type_28; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_223;
  reg [1:0] btb_bj_type_29; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_224;
  reg [1:0] btb_bj_type_30; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_225;
  reg [1:0] btb_bj_type_31; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_226;
  reg [1:0] btb_bj_type_32; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_227;
  reg [1:0] btb_bj_type_33; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_228;
  reg [1:0] btb_bj_type_34; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_229;
  reg [1:0] btb_bj_type_35; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_230;
  reg [1:0] btb_bj_type_36; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_231;
  reg [1:0] btb_bj_type_37; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_232;
  reg [1:0] btb_bj_type_38; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_233;
  reg [1:0] btb_bj_type_39; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_234;
  reg [1:0] btb_bj_type_40; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_235;
  reg [1:0] btb_bj_type_41; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_236;
  reg [1:0] btb_bj_type_42; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_237;
  reg [1:0] btb_bj_type_43; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_238;
  reg [1:0] btb_bj_type_44; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_239;
  reg [1:0] btb_bj_type_45; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_240;
  reg [1:0] btb_bj_type_46; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_241;
  reg [1:0] btb_bj_type_47; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_242;
  reg [1:0] btb_bj_type_48; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_243;
  reg [1:0] btb_bj_type_49; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_244;
  reg [1:0] btb_bj_type_50; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_245;
  reg [1:0] btb_bj_type_51; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_246;
  reg [1:0] btb_bj_type_52; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_247;
  reg [1:0] btb_bj_type_53; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_248;
  reg [1:0] btb_bj_type_54; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_249;
  reg [1:0] btb_bj_type_55; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_250;
  reg [1:0] btb_bj_type_56; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_251;
  reg [1:0] btb_bj_type_57; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_252;
  reg [1:0] btb_bj_type_58; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_253;
  reg [1:0] btb_bj_type_59; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_254;
  reg [1:0] btb_bj_type_60; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_255;
  reg [1:0] btb_bj_type_61; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_256;
  reg [1:0] btb_bj_type_62; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_257;
  reg [1:0] btb_bj_type_63; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_258;
  reg [1:0] btb_h_count_0; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_259;
  reg [1:0] btb_h_count_1; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_260;
  reg [1:0] btb_h_count_2; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_261;
  reg [1:0] btb_h_count_3; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_262;
  reg [1:0] btb_h_count_4; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_263;
  reg [1:0] btb_h_count_5; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_264;
  reg [1:0] btb_h_count_6; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_265;
  reg [1:0] btb_h_count_7; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_266;
  reg [1:0] btb_h_count_8; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_267;
  reg [1:0] btb_h_count_9; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_268;
  reg [1:0] btb_h_count_10; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_269;
  reg [1:0] btb_h_count_11; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_270;
  reg [1:0] btb_h_count_12; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_271;
  reg [1:0] btb_h_count_13; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_272;
  reg [1:0] btb_h_count_14; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_273;
  reg [1:0] btb_h_count_15; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_274;
  reg [1:0] btb_h_count_16; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_275;
  reg [1:0] btb_h_count_17; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_276;
  reg [1:0] btb_h_count_18; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_277;
  reg [1:0] btb_h_count_19; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_278;
  reg [1:0] btb_h_count_20; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_279;
  reg [1:0] btb_h_count_21; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_280;
  reg [1:0] btb_h_count_22; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_281;
  reg [1:0] btb_h_count_23; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_282;
  reg [1:0] btb_h_count_24; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_283;
  reg [1:0] btb_h_count_25; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_284;
  reg [1:0] btb_h_count_26; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_285;
  reg [1:0] btb_h_count_27; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_286;
  reg [1:0] btb_h_count_28; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_287;
  reg [1:0] btb_h_count_29; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_288;
  reg [1:0] btb_h_count_30; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_289;
  reg [1:0] btb_h_count_31; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_290;
  reg [1:0] btb_h_count_32; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_291;
  reg [1:0] btb_h_count_33; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_292;
  reg [1:0] btb_h_count_34; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_293;
  reg [1:0] btb_h_count_35; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_294;
  reg [1:0] btb_h_count_36; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_295;
  reg [1:0] btb_h_count_37; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_296;
  reg [1:0] btb_h_count_38; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_297;
  reg [1:0] btb_h_count_39; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_298;
  reg [1:0] btb_h_count_40; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_299;
  reg [1:0] btb_h_count_41; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_300;
  reg [1:0] btb_h_count_42; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_301;
  reg [1:0] btb_h_count_43; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_302;
  reg [1:0] btb_h_count_44; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_303;
  reg [1:0] btb_h_count_45; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_304;
  reg [1:0] btb_h_count_46; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_305;
  reg [1:0] btb_h_count_47; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_306;
  reg [1:0] btb_h_count_48; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_307;
  reg [1:0] btb_h_count_49; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_308;
  reg [1:0] btb_h_count_50; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_309;
  reg [1:0] btb_h_count_51; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_310;
  reg [1:0] btb_h_count_52; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_311;
  reg [1:0] btb_h_count_53; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_312;
  reg [1:0] btb_h_count_54; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_313;
  reg [1:0] btb_h_count_55; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_314;
  reg [1:0] btb_h_count_56; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_315;
  reg [1:0] btb_h_count_57; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_316;
  reg [1:0] btb_h_count_58; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_317;
  reg [1:0] btb_h_count_59; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_318;
  reg [1:0] btb_h_count_60; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_319;
  reg [1:0] btb_h_count_61; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_320;
  reg [1:0] btb_h_count_62; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_321;
  reg [1:0] btb_h_count_63; // @[BTB.scala 72:20:@381.4]
  reg [31:0] _RAND_322;
  wire [32:0] _T_148; // @[BTB.scala 102:32:@383.4]
  wire [31:0] predict_cont_tgt; // @[BTB.scala 102:32:@384.4]
  wire  _T_150; // @[BTB.scala 103:42:@386.4]
  wire  _T_151; // @[BTB.scala 103:42:@387.4]
  wire  _T_152; // @[BTB.scala 103:42:@388.4]
  wire  _T_153; // @[BTB.scala 103:42:@389.4]
  wire  _T_154; // @[BTB.scala 103:42:@390.4]
  wire  _T_155; // @[BTB.scala 103:42:@391.4]
  wire  _T_156; // @[BTB.scala 103:42:@392.4]
  wire  _T_157; // @[BTB.scala 103:42:@393.4]
  wire  _T_158; // @[BTB.scala 103:42:@394.4]
  wire  _T_159; // @[BTB.scala 103:42:@395.4]
  wire  _T_160; // @[BTB.scala 103:42:@396.4]
  wire  _T_161; // @[BTB.scala 103:42:@397.4]
  wire  _T_162; // @[BTB.scala 103:42:@398.4]
  wire  _T_163; // @[BTB.scala 103:42:@399.4]
  wire  _T_164; // @[BTB.scala 103:42:@400.4]
  wire  _T_165; // @[BTB.scala 103:42:@401.4]
  wire  _T_166; // @[BTB.scala 103:42:@402.4]
  wire  _T_167; // @[BTB.scala 103:42:@403.4]
  wire  _T_168; // @[BTB.scala 103:42:@404.4]
  wire  _T_169; // @[BTB.scala 103:42:@405.4]
  wire  _T_170; // @[BTB.scala 103:42:@406.4]
  wire  _T_171; // @[BTB.scala 103:42:@407.4]
  wire  _T_172; // @[BTB.scala 103:42:@408.4]
  wire  _T_173; // @[BTB.scala 103:42:@409.4]
  wire  _T_174; // @[BTB.scala 103:42:@410.4]
  wire  _T_175; // @[BTB.scala 103:42:@411.4]
  wire  _T_176; // @[BTB.scala 103:42:@412.4]
  wire  _T_177; // @[BTB.scala 103:42:@413.4]
  wire  _T_178; // @[BTB.scala 103:42:@414.4]
  wire  _T_179; // @[BTB.scala 103:42:@415.4]
  wire  _T_180; // @[BTB.scala 103:42:@416.4]
  wire  _T_181; // @[BTB.scala 103:42:@417.4]
  wire  _T_182; // @[BTB.scala 103:42:@418.4]
  wire  _T_183; // @[BTB.scala 103:42:@419.4]
  wire  _T_184; // @[BTB.scala 103:42:@420.4]
  wire  _T_185; // @[BTB.scala 103:42:@421.4]
  wire  _T_186; // @[BTB.scala 103:42:@422.4]
  wire  _T_187; // @[BTB.scala 103:42:@423.4]
  wire  _T_188; // @[BTB.scala 103:42:@424.4]
  wire  _T_189; // @[BTB.scala 103:42:@425.4]
  wire  _T_190; // @[BTB.scala 103:42:@426.4]
  wire  _T_191; // @[BTB.scala 103:42:@427.4]
  wire  _T_192; // @[BTB.scala 103:42:@428.4]
  wire  _T_193; // @[BTB.scala 103:42:@429.4]
  wire  _T_194; // @[BTB.scala 103:42:@430.4]
  wire  _T_195; // @[BTB.scala 103:42:@431.4]
  wire  _T_196; // @[BTB.scala 103:42:@432.4]
  wire  _T_197; // @[BTB.scala 103:42:@433.4]
  wire  _T_198; // @[BTB.scala 103:42:@434.4]
  wire  _T_199; // @[BTB.scala 103:42:@435.4]
  wire  _T_200; // @[BTB.scala 103:42:@436.4]
  wire  _T_201; // @[BTB.scala 103:42:@437.4]
  wire  _T_202; // @[BTB.scala 103:42:@438.4]
  wire  _T_203; // @[BTB.scala 103:42:@439.4]
  wire  _T_204; // @[BTB.scala 103:42:@440.4]
  wire  _T_205; // @[BTB.scala 103:42:@441.4]
  wire  _T_206; // @[BTB.scala 103:42:@442.4]
  wire  _T_207; // @[BTB.scala 103:42:@443.4]
  wire  _T_208; // @[BTB.scala 103:42:@444.4]
  wire  _T_209; // @[BTB.scala 103:42:@445.4]
  wire  _T_210; // @[BTB.scala 103:42:@446.4]
  wire  _T_211; // @[BTB.scala 103:42:@447.4]
  wire  _T_212; // @[BTB.scala 103:42:@448.4]
  wire  _T_213; // @[BTB.scala 103:42:@449.4]
  wire [7:0] _T_290; // @[BTB.scala 103:57:@521.4]
  wire [15:0] _T_298; // @[BTB.scala 103:57:@529.4]
  wire [7:0] _T_305; // @[BTB.scala 103:57:@536.4]
  wire [31:0] _T_314; // @[BTB.scala 103:57:@545.4]
  wire [7:0] _T_321; // @[BTB.scala 103:57:@552.4]
  wire [15:0] _T_329; // @[BTB.scala 103:57:@560.4]
  wire [7:0] _T_336; // @[BTB.scala 103:57:@567.4]
  wire [31:0] _T_345; // @[BTB.scala 103:57:@576.4]
  wire [63:0] _T_346; // @[BTB.scala 103:57:@577.4]
  wire [7:0] _T_353; // @[BTB.scala 103:76:@584.4]
  wire [15:0] _T_361; // @[BTB.scala 103:76:@592.4]
  wire [7:0] _T_368; // @[BTB.scala 103:76:@599.4]
  wire [31:0] _T_377; // @[BTB.scala 103:76:@608.4]
  wire [7:0] _T_384; // @[BTB.scala 103:76:@615.4]
  wire [15:0] _T_392; // @[BTB.scala 103:76:@623.4]
  wire [7:0] _T_399; // @[BTB.scala 103:76:@630.4]
  wire [31:0] _T_408; // @[BTB.scala 103:76:@639.4]
  wire [63:0] _T_409; // @[BTB.scala 103:76:@640.4]
  wire [63:0] predict_lookup; // @[BTB.scala 103:64:@641.4]
  wire  _T_411; // @[Mux.scala 21:36:@643.4]
  wire  _T_412; // @[Mux.scala 21:36:@644.4]
  wire  _T_413; // @[Mux.scala 21:36:@645.4]
  wire  _T_414; // @[Mux.scala 21:36:@646.4]
  wire  _T_415; // @[Mux.scala 21:36:@647.4]
  wire  _T_416; // @[Mux.scala 21:36:@648.4]
  wire  _T_417; // @[Mux.scala 21:36:@649.4]
  wire  _T_418; // @[Mux.scala 21:36:@650.4]
  wire  _T_419; // @[Mux.scala 21:36:@651.4]
  wire  _T_420; // @[Mux.scala 21:36:@652.4]
  wire  _T_421; // @[Mux.scala 21:36:@653.4]
  wire  _T_422; // @[Mux.scala 21:36:@654.4]
  wire  _T_423; // @[Mux.scala 21:36:@655.4]
  wire  _T_424; // @[Mux.scala 21:36:@656.4]
  wire  _T_425; // @[Mux.scala 21:36:@657.4]
  wire  _T_426; // @[Mux.scala 21:36:@658.4]
  wire  _T_427; // @[Mux.scala 21:36:@659.4]
  wire  _T_428; // @[Mux.scala 21:36:@660.4]
  wire  _T_429; // @[Mux.scala 21:36:@661.4]
  wire  _T_430; // @[Mux.scala 21:36:@662.4]
  wire  _T_431; // @[Mux.scala 21:36:@663.4]
  wire  _T_432; // @[Mux.scala 21:36:@664.4]
  wire  _T_433; // @[Mux.scala 21:36:@665.4]
  wire  _T_434; // @[Mux.scala 21:36:@666.4]
  wire  _T_435; // @[Mux.scala 21:36:@667.4]
  wire  _T_436; // @[Mux.scala 21:36:@668.4]
  wire  _T_437; // @[Mux.scala 21:36:@669.4]
  wire  _T_438; // @[Mux.scala 21:36:@670.4]
  wire  _T_439; // @[Mux.scala 21:36:@671.4]
  wire  _T_440; // @[Mux.scala 21:36:@672.4]
  wire  _T_441; // @[Mux.scala 21:36:@673.4]
  wire  _T_442; // @[Mux.scala 21:36:@674.4]
  wire  _T_443; // @[Mux.scala 21:36:@675.4]
  wire  _T_444; // @[Mux.scala 21:36:@676.4]
  wire  _T_445; // @[Mux.scala 21:36:@677.4]
  wire  _T_446; // @[Mux.scala 21:36:@678.4]
  wire  _T_447; // @[Mux.scala 21:36:@679.4]
  wire  _T_448; // @[Mux.scala 21:36:@680.4]
  wire  _T_449; // @[Mux.scala 21:36:@681.4]
  wire  _T_450; // @[Mux.scala 21:36:@682.4]
  wire  _T_451; // @[Mux.scala 21:36:@683.4]
  wire  _T_452; // @[Mux.scala 21:36:@684.4]
  wire  _T_453; // @[Mux.scala 21:36:@685.4]
  wire  _T_454; // @[Mux.scala 21:36:@686.4]
  wire  _T_455; // @[Mux.scala 21:36:@687.4]
  wire  _T_456; // @[Mux.scala 21:36:@688.4]
  wire  _T_457; // @[Mux.scala 21:36:@689.4]
  wire  _T_458; // @[Mux.scala 21:36:@690.4]
  wire  _T_459; // @[Mux.scala 21:36:@691.4]
  wire  _T_460; // @[Mux.scala 21:36:@692.4]
  wire  _T_461; // @[Mux.scala 21:36:@693.4]
  wire  _T_462; // @[Mux.scala 21:36:@694.4]
  wire  _T_463; // @[Mux.scala 21:36:@695.4]
  wire  _T_464; // @[Mux.scala 21:36:@696.4]
  wire  _T_465; // @[Mux.scala 21:36:@697.4]
  wire  _T_466; // @[Mux.scala 21:36:@698.4]
  wire  _T_467; // @[Mux.scala 21:36:@699.4]
  wire  _T_468; // @[Mux.scala 21:36:@700.4]
  wire  _T_469; // @[Mux.scala 21:36:@701.4]
  wire  _T_470; // @[Mux.scala 21:36:@702.4]
  wire  _T_471; // @[Mux.scala 21:36:@703.4]
  wire  _T_472; // @[Mux.scala 21:36:@704.4]
  wire  _T_473; // @[Mux.scala 21:36:@705.4]
  wire  _T_474; // @[Mux.scala 21:36:@706.4]
  wire [31:0] _T_477; // @[Mux.scala 19:72:@707.4]
  wire [31:0] _T_479; // @[Mux.scala 19:72:@708.4]
  wire [31:0] _T_481; // @[Mux.scala 19:72:@709.4]
  wire [31:0] _T_483; // @[Mux.scala 19:72:@710.4]
  wire [31:0] _T_485; // @[Mux.scala 19:72:@711.4]
  wire [31:0] _T_487; // @[Mux.scala 19:72:@712.4]
  wire [31:0] _T_489; // @[Mux.scala 19:72:@713.4]
  wire [31:0] _T_491; // @[Mux.scala 19:72:@714.4]
  wire [31:0] _T_493; // @[Mux.scala 19:72:@715.4]
  wire [31:0] _T_495; // @[Mux.scala 19:72:@716.4]
  wire [31:0] _T_497; // @[Mux.scala 19:72:@717.4]
  wire [31:0] _T_499; // @[Mux.scala 19:72:@718.4]
  wire [31:0] _T_501; // @[Mux.scala 19:72:@719.4]
  wire [31:0] _T_503; // @[Mux.scala 19:72:@720.4]
  wire [31:0] _T_505; // @[Mux.scala 19:72:@721.4]
  wire [31:0] _T_507; // @[Mux.scala 19:72:@722.4]
  wire [31:0] _T_509; // @[Mux.scala 19:72:@723.4]
  wire [31:0] _T_511; // @[Mux.scala 19:72:@724.4]
  wire [31:0] _T_513; // @[Mux.scala 19:72:@725.4]
  wire [31:0] _T_515; // @[Mux.scala 19:72:@726.4]
  wire [31:0] _T_517; // @[Mux.scala 19:72:@727.4]
  wire [31:0] _T_519; // @[Mux.scala 19:72:@728.4]
  wire [31:0] _T_521; // @[Mux.scala 19:72:@729.4]
  wire [31:0] _T_523; // @[Mux.scala 19:72:@730.4]
  wire [31:0] _T_525; // @[Mux.scala 19:72:@731.4]
  wire [31:0] _T_527; // @[Mux.scala 19:72:@732.4]
  wire [31:0] _T_529; // @[Mux.scala 19:72:@733.4]
  wire [31:0] _T_531; // @[Mux.scala 19:72:@734.4]
  wire [31:0] _T_533; // @[Mux.scala 19:72:@735.4]
  wire [31:0] _T_535; // @[Mux.scala 19:72:@736.4]
  wire [31:0] _T_537; // @[Mux.scala 19:72:@737.4]
  wire [31:0] _T_539; // @[Mux.scala 19:72:@738.4]
  wire [31:0] _T_541; // @[Mux.scala 19:72:@739.4]
  wire [31:0] _T_543; // @[Mux.scala 19:72:@740.4]
  wire [31:0] _T_545; // @[Mux.scala 19:72:@741.4]
  wire [31:0] _T_547; // @[Mux.scala 19:72:@742.4]
  wire [31:0] _T_549; // @[Mux.scala 19:72:@743.4]
  wire [31:0] _T_551; // @[Mux.scala 19:72:@744.4]
  wire [31:0] _T_553; // @[Mux.scala 19:72:@745.4]
  wire [31:0] _T_555; // @[Mux.scala 19:72:@746.4]
  wire [31:0] _T_557; // @[Mux.scala 19:72:@747.4]
  wire [31:0] _T_559; // @[Mux.scala 19:72:@748.4]
  wire [31:0] _T_561; // @[Mux.scala 19:72:@749.4]
  wire [31:0] _T_563; // @[Mux.scala 19:72:@750.4]
  wire [31:0] _T_565; // @[Mux.scala 19:72:@751.4]
  wire [31:0] _T_567; // @[Mux.scala 19:72:@752.4]
  wire [31:0] _T_569; // @[Mux.scala 19:72:@753.4]
  wire [31:0] _T_571; // @[Mux.scala 19:72:@754.4]
  wire [31:0] _T_573; // @[Mux.scala 19:72:@755.4]
  wire [31:0] _T_575; // @[Mux.scala 19:72:@756.4]
  wire [31:0] _T_577; // @[Mux.scala 19:72:@757.4]
  wire [31:0] _T_579; // @[Mux.scala 19:72:@758.4]
  wire [31:0] _T_581; // @[Mux.scala 19:72:@759.4]
  wire [31:0] _T_583; // @[Mux.scala 19:72:@760.4]
  wire [31:0] _T_585; // @[Mux.scala 19:72:@761.4]
  wire [31:0] _T_587; // @[Mux.scala 19:72:@762.4]
  wire [31:0] _T_589; // @[Mux.scala 19:72:@763.4]
  wire [31:0] _T_591; // @[Mux.scala 19:72:@764.4]
  wire [31:0] _T_593; // @[Mux.scala 19:72:@765.4]
  wire [31:0] _T_595; // @[Mux.scala 19:72:@766.4]
  wire [31:0] _T_597; // @[Mux.scala 19:72:@767.4]
  wire [31:0] _T_599; // @[Mux.scala 19:72:@768.4]
  wire [31:0] _T_601; // @[Mux.scala 19:72:@769.4]
  wire [31:0] _T_603; // @[Mux.scala 19:72:@770.4]
  wire [31:0] _T_604; // @[Mux.scala 19:72:@771.4]
  wire [31:0] _T_605; // @[Mux.scala 19:72:@772.4]
  wire [31:0] _T_606; // @[Mux.scala 19:72:@773.4]
  wire [31:0] _T_607; // @[Mux.scala 19:72:@774.4]
  wire [31:0] _T_608; // @[Mux.scala 19:72:@775.4]
  wire [31:0] _T_609; // @[Mux.scala 19:72:@776.4]
  wire [31:0] _T_610; // @[Mux.scala 19:72:@777.4]
  wire [31:0] _T_611; // @[Mux.scala 19:72:@778.4]
  wire [31:0] _T_612; // @[Mux.scala 19:72:@779.4]
  wire [31:0] _T_613; // @[Mux.scala 19:72:@780.4]
  wire [31:0] _T_614; // @[Mux.scala 19:72:@781.4]
  wire [31:0] _T_615; // @[Mux.scala 19:72:@782.4]
  wire [31:0] _T_616; // @[Mux.scala 19:72:@783.4]
  wire [31:0] _T_617; // @[Mux.scala 19:72:@784.4]
  wire [31:0] _T_618; // @[Mux.scala 19:72:@785.4]
  wire [31:0] _T_619; // @[Mux.scala 19:72:@786.4]
  wire [31:0] _T_620; // @[Mux.scala 19:72:@787.4]
  wire [31:0] _T_621; // @[Mux.scala 19:72:@788.4]
  wire [31:0] _T_622; // @[Mux.scala 19:72:@789.4]
  wire [31:0] _T_623; // @[Mux.scala 19:72:@790.4]
  wire [31:0] _T_624; // @[Mux.scala 19:72:@791.4]
  wire [31:0] _T_625; // @[Mux.scala 19:72:@792.4]
  wire [31:0] _T_626; // @[Mux.scala 19:72:@793.4]
  wire [31:0] _T_627; // @[Mux.scala 19:72:@794.4]
  wire [31:0] _T_628; // @[Mux.scala 19:72:@795.4]
  wire [31:0] _T_629; // @[Mux.scala 19:72:@796.4]
  wire [31:0] _T_630; // @[Mux.scala 19:72:@797.4]
  wire [31:0] _T_631; // @[Mux.scala 19:72:@798.4]
  wire [31:0] _T_632; // @[Mux.scala 19:72:@799.4]
  wire [31:0] _T_633; // @[Mux.scala 19:72:@800.4]
  wire [31:0] _T_634; // @[Mux.scala 19:72:@801.4]
  wire [31:0] _T_635; // @[Mux.scala 19:72:@802.4]
  wire [31:0] _T_636; // @[Mux.scala 19:72:@803.4]
  wire [31:0] _T_637; // @[Mux.scala 19:72:@804.4]
  wire [31:0] _T_638; // @[Mux.scala 19:72:@805.4]
  wire [31:0] _T_639; // @[Mux.scala 19:72:@806.4]
  wire [31:0] _T_640; // @[Mux.scala 19:72:@807.4]
  wire [31:0] _T_641; // @[Mux.scala 19:72:@808.4]
  wire [31:0] _T_642; // @[Mux.scala 19:72:@809.4]
  wire [31:0] _T_643; // @[Mux.scala 19:72:@810.4]
  wire [31:0] _T_644; // @[Mux.scala 19:72:@811.4]
  wire [31:0] _T_645; // @[Mux.scala 19:72:@812.4]
  wire [31:0] _T_646; // @[Mux.scala 19:72:@813.4]
  wire [31:0] _T_647; // @[Mux.scala 19:72:@814.4]
  wire [31:0] _T_648; // @[Mux.scala 19:72:@815.4]
  wire [31:0] _T_649; // @[Mux.scala 19:72:@816.4]
  wire [31:0] _T_650; // @[Mux.scala 19:72:@817.4]
  wire [31:0] _T_651; // @[Mux.scala 19:72:@818.4]
  wire [31:0] _T_652; // @[Mux.scala 19:72:@819.4]
  wire [31:0] _T_653; // @[Mux.scala 19:72:@820.4]
  wire [31:0] _T_654; // @[Mux.scala 19:72:@821.4]
  wire [31:0] _T_655; // @[Mux.scala 19:72:@822.4]
  wire [31:0] _T_656; // @[Mux.scala 19:72:@823.4]
  wire [31:0] _T_657; // @[Mux.scala 19:72:@824.4]
  wire [31:0] _T_658; // @[Mux.scala 19:72:@825.4]
  wire [31:0] _T_659; // @[Mux.scala 19:72:@826.4]
  wire [31:0] _T_660; // @[Mux.scala 19:72:@827.4]
  wire [31:0] _T_661; // @[Mux.scala 19:72:@828.4]
  wire [31:0] _T_662; // @[Mux.scala 19:72:@829.4]
  wire [31:0] _T_663; // @[Mux.scala 19:72:@830.4]
  wire [31:0] _T_664; // @[Mux.scala 19:72:@831.4]
  wire [31:0] _T_665; // @[Mux.scala 19:72:@832.4]
  wire [31:0] predict_jump_tgt; // @[Mux.scala 19:72:@833.4]
  wire [1:0] _T_735; // @[Mux.scala 19:72:@901.4]
  wire [1:0] _T_737; // @[Mux.scala 19:72:@902.4]
  wire [1:0] _T_739; // @[Mux.scala 19:72:@903.4]
  wire [1:0] _T_741; // @[Mux.scala 19:72:@904.4]
  wire [1:0] _T_743; // @[Mux.scala 19:72:@905.4]
  wire [1:0] _T_745; // @[Mux.scala 19:72:@906.4]
  wire [1:0] _T_747; // @[Mux.scala 19:72:@907.4]
  wire [1:0] _T_749; // @[Mux.scala 19:72:@908.4]
  wire [1:0] _T_751; // @[Mux.scala 19:72:@909.4]
  wire [1:0] _T_753; // @[Mux.scala 19:72:@910.4]
  wire [1:0] _T_755; // @[Mux.scala 19:72:@911.4]
  wire [1:0] _T_757; // @[Mux.scala 19:72:@912.4]
  wire [1:0] _T_759; // @[Mux.scala 19:72:@913.4]
  wire [1:0] _T_761; // @[Mux.scala 19:72:@914.4]
  wire [1:0] _T_763; // @[Mux.scala 19:72:@915.4]
  wire [1:0] _T_765; // @[Mux.scala 19:72:@916.4]
  wire [1:0] _T_767; // @[Mux.scala 19:72:@917.4]
  wire [1:0] _T_769; // @[Mux.scala 19:72:@918.4]
  wire [1:0] _T_771; // @[Mux.scala 19:72:@919.4]
  wire [1:0] _T_773; // @[Mux.scala 19:72:@920.4]
  wire [1:0] _T_775; // @[Mux.scala 19:72:@921.4]
  wire [1:0] _T_777; // @[Mux.scala 19:72:@922.4]
  wire [1:0] _T_779; // @[Mux.scala 19:72:@923.4]
  wire [1:0] _T_781; // @[Mux.scala 19:72:@924.4]
  wire [1:0] _T_783; // @[Mux.scala 19:72:@925.4]
  wire [1:0] _T_785; // @[Mux.scala 19:72:@926.4]
  wire [1:0] _T_787; // @[Mux.scala 19:72:@927.4]
  wire [1:0] _T_789; // @[Mux.scala 19:72:@928.4]
  wire [1:0] _T_791; // @[Mux.scala 19:72:@929.4]
  wire [1:0] _T_793; // @[Mux.scala 19:72:@930.4]
  wire [1:0] _T_795; // @[Mux.scala 19:72:@931.4]
  wire [1:0] _T_797; // @[Mux.scala 19:72:@932.4]
  wire [1:0] _T_799; // @[Mux.scala 19:72:@933.4]
  wire [1:0] _T_801; // @[Mux.scala 19:72:@934.4]
  wire [1:0] _T_803; // @[Mux.scala 19:72:@935.4]
  wire [1:0] _T_805; // @[Mux.scala 19:72:@936.4]
  wire [1:0] _T_807; // @[Mux.scala 19:72:@937.4]
  wire [1:0] _T_809; // @[Mux.scala 19:72:@938.4]
  wire [1:0] _T_811; // @[Mux.scala 19:72:@939.4]
  wire [1:0] _T_813; // @[Mux.scala 19:72:@940.4]
  wire [1:0] _T_815; // @[Mux.scala 19:72:@941.4]
  wire [1:0] _T_817; // @[Mux.scala 19:72:@942.4]
  wire [1:0] _T_819; // @[Mux.scala 19:72:@943.4]
  wire [1:0] _T_821; // @[Mux.scala 19:72:@944.4]
  wire [1:0] _T_823; // @[Mux.scala 19:72:@945.4]
  wire [1:0] _T_825; // @[Mux.scala 19:72:@946.4]
  wire [1:0] _T_827; // @[Mux.scala 19:72:@947.4]
  wire [1:0] _T_829; // @[Mux.scala 19:72:@948.4]
  wire [1:0] _T_831; // @[Mux.scala 19:72:@949.4]
  wire [1:0] _T_833; // @[Mux.scala 19:72:@950.4]
  wire [1:0] _T_835; // @[Mux.scala 19:72:@951.4]
  wire [1:0] _T_837; // @[Mux.scala 19:72:@952.4]
  wire [1:0] _T_839; // @[Mux.scala 19:72:@953.4]
  wire [1:0] _T_841; // @[Mux.scala 19:72:@954.4]
  wire [1:0] _T_843; // @[Mux.scala 19:72:@955.4]
  wire [1:0] _T_845; // @[Mux.scala 19:72:@956.4]
  wire [1:0] _T_847; // @[Mux.scala 19:72:@957.4]
  wire [1:0] _T_849; // @[Mux.scala 19:72:@958.4]
  wire [1:0] _T_851; // @[Mux.scala 19:72:@959.4]
  wire [1:0] _T_853; // @[Mux.scala 19:72:@960.4]
  wire [1:0] _T_855; // @[Mux.scala 19:72:@961.4]
  wire [1:0] _T_857; // @[Mux.scala 19:72:@962.4]
  wire [1:0] _T_859; // @[Mux.scala 19:72:@963.4]
  wire [1:0] _T_861; // @[Mux.scala 19:72:@964.4]
  wire [1:0] _T_862; // @[Mux.scala 19:72:@965.4]
  wire [1:0] _T_863; // @[Mux.scala 19:72:@966.4]
  wire [1:0] _T_864; // @[Mux.scala 19:72:@967.4]
  wire [1:0] _T_865; // @[Mux.scala 19:72:@968.4]
  wire [1:0] _T_866; // @[Mux.scala 19:72:@969.4]
  wire [1:0] _T_867; // @[Mux.scala 19:72:@970.4]
  wire [1:0] _T_868; // @[Mux.scala 19:72:@971.4]
  wire [1:0] _T_869; // @[Mux.scala 19:72:@972.4]
  wire [1:0] _T_870; // @[Mux.scala 19:72:@973.4]
  wire [1:0] _T_871; // @[Mux.scala 19:72:@974.4]
  wire [1:0] _T_872; // @[Mux.scala 19:72:@975.4]
  wire [1:0] _T_873; // @[Mux.scala 19:72:@976.4]
  wire [1:0] _T_874; // @[Mux.scala 19:72:@977.4]
  wire [1:0] _T_875; // @[Mux.scala 19:72:@978.4]
  wire [1:0] _T_876; // @[Mux.scala 19:72:@979.4]
  wire [1:0] _T_877; // @[Mux.scala 19:72:@980.4]
  wire [1:0] _T_878; // @[Mux.scala 19:72:@981.4]
  wire [1:0] _T_879; // @[Mux.scala 19:72:@982.4]
  wire [1:0] _T_880; // @[Mux.scala 19:72:@983.4]
  wire [1:0] _T_881; // @[Mux.scala 19:72:@984.4]
  wire [1:0] _T_882; // @[Mux.scala 19:72:@985.4]
  wire [1:0] _T_883; // @[Mux.scala 19:72:@986.4]
  wire [1:0] _T_884; // @[Mux.scala 19:72:@987.4]
  wire [1:0] _T_885; // @[Mux.scala 19:72:@988.4]
  wire [1:0] _T_886; // @[Mux.scala 19:72:@989.4]
  wire [1:0] _T_887; // @[Mux.scala 19:72:@990.4]
  wire [1:0] _T_888; // @[Mux.scala 19:72:@991.4]
  wire [1:0] _T_889; // @[Mux.scala 19:72:@992.4]
  wire [1:0] _T_890; // @[Mux.scala 19:72:@993.4]
  wire [1:0] _T_891; // @[Mux.scala 19:72:@994.4]
  wire [1:0] _T_892; // @[Mux.scala 19:72:@995.4]
  wire [1:0] _T_893; // @[Mux.scala 19:72:@996.4]
  wire [1:0] _T_894; // @[Mux.scala 19:72:@997.4]
  wire [1:0] _T_895; // @[Mux.scala 19:72:@998.4]
  wire [1:0] _T_896; // @[Mux.scala 19:72:@999.4]
  wire [1:0] _T_897; // @[Mux.scala 19:72:@1000.4]
  wire [1:0] _T_898; // @[Mux.scala 19:72:@1001.4]
  wire [1:0] _T_899; // @[Mux.scala 19:72:@1002.4]
  wire [1:0] _T_900; // @[Mux.scala 19:72:@1003.4]
  wire [1:0] _T_901; // @[Mux.scala 19:72:@1004.4]
  wire [1:0] _T_902; // @[Mux.scala 19:72:@1005.4]
  wire [1:0] _T_903; // @[Mux.scala 19:72:@1006.4]
  wire [1:0] _T_904; // @[Mux.scala 19:72:@1007.4]
  wire [1:0] _T_905; // @[Mux.scala 19:72:@1008.4]
  wire [1:0] _T_906; // @[Mux.scala 19:72:@1009.4]
  wire [1:0] _T_907; // @[Mux.scala 19:72:@1010.4]
  wire [1:0] _T_908; // @[Mux.scala 19:72:@1011.4]
  wire [1:0] _T_909; // @[Mux.scala 19:72:@1012.4]
  wire [1:0] _T_910; // @[Mux.scala 19:72:@1013.4]
  wire [1:0] _T_911; // @[Mux.scala 19:72:@1014.4]
  wire [1:0] _T_912; // @[Mux.scala 19:72:@1015.4]
  wire [1:0] _T_913; // @[Mux.scala 19:72:@1016.4]
  wire [1:0] _T_914; // @[Mux.scala 19:72:@1017.4]
  wire [1:0] _T_915; // @[Mux.scala 19:72:@1018.4]
  wire [1:0] _T_916; // @[Mux.scala 19:72:@1019.4]
  wire [1:0] _T_917; // @[Mux.scala 19:72:@1020.4]
  wire [1:0] _T_918; // @[Mux.scala 19:72:@1021.4]
  wire [1:0] _T_919; // @[Mux.scala 19:72:@1022.4]
  wire [1:0] _T_920; // @[Mux.scala 19:72:@1023.4]
  wire [1:0] _T_921; // @[Mux.scala 19:72:@1024.4]
  wire [1:0] _T_922; // @[Mux.scala 19:72:@1025.4]
  wire [1:0] _T_923; // @[Mux.scala 19:72:@1026.4]
  wire [1:0] predict_bj_type; // @[Mux.scala 19:72:@1027.4]
  wire [1:0] _T_993; // @[Mux.scala 19:72:@1095.4]
  wire [1:0] _T_995; // @[Mux.scala 19:72:@1096.4]
  wire [1:0] _T_997; // @[Mux.scala 19:72:@1097.4]
  wire [1:0] _T_999; // @[Mux.scala 19:72:@1098.4]
  wire [1:0] _T_1001; // @[Mux.scala 19:72:@1099.4]
  wire [1:0] _T_1003; // @[Mux.scala 19:72:@1100.4]
  wire [1:0] _T_1005; // @[Mux.scala 19:72:@1101.4]
  wire [1:0] _T_1007; // @[Mux.scala 19:72:@1102.4]
  wire [1:0] _T_1009; // @[Mux.scala 19:72:@1103.4]
  wire [1:0] _T_1011; // @[Mux.scala 19:72:@1104.4]
  wire [1:0] _T_1013; // @[Mux.scala 19:72:@1105.4]
  wire [1:0] _T_1015; // @[Mux.scala 19:72:@1106.4]
  wire [1:0] _T_1017; // @[Mux.scala 19:72:@1107.4]
  wire [1:0] _T_1019; // @[Mux.scala 19:72:@1108.4]
  wire [1:0] _T_1021; // @[Mux.scala 19:72:@1109.4]
  wire [1:0] _T_1023; // @[Mux.scala 19:72:@1110.4]
  wire [1:0] _T_1025; // @[Mux.scala 19:72:@1111.4]
  wire [1:0] _T_1027; // @[Mux.scala 19:72:@1112.4]
  wire [1:0] _T_1029; // @[Mux.scala 19:72:@1113.4]
  wire [1:0] _T_1031; // @[Mux.scala 19:72:@1114.4]
  wire [1:0] _T_1033; // @[Mux.scala 19:72:@1115.4]
  wire [1:0] _T_1035; // @[Mux.scala 19:72:@1116.4]
  wire [1:0] _T_1037; // @[Mux.scala 19:72:@1117.4]
  wire [1:0] _T_1039; // @[Mux.scala 19:72:@1118.4]
  wire [1:0] _T_1041; // @[Mux.scala 19:72:@1119.4]
  wire [1:0] _T_1043; // @[Mux.scala 19:72:@1120.4]
  wire [1:0] _T_1045; // @[Mux.scala 19:72:@1121.4]
  wire [1:0] _T_1047; // @[Mux.scala 19:72:@1122.4]
  wire [1:0] _T_1049; // @[Mux.scala 19:72:@1123.4]
  wire [1:0] _T_1051; // @[Mux.scala 19:72:@1124.4]
  wire [1:0] _T_1053; // @[Mux.scala 19:72:@1125.4]
  wire [1:0] _T_1055; // @[Mux.scala 19:72:@1126.4]
  wire [1:0] _T_1057; // @[Mux.scala 19:72:@1127.4]
  wire [1:0] _T_1059; // @[Mux.scala 19:72:@1128.4]
  wire [1:0] _T_1061; // @[Mux.scala 19:72:@1129.4]
  wire [1:0] _T_1063; // @[Mux.scala 19:72:@1130.4]
  wire [1:0] _T_1065; // @[Mux.scala 19:72:@1131.4]
  wire [1:0] _T_1067; // @[Mux.scala 19:72:@1132.4]
  wire [1:0] _T_1069; // @[Mux.scala 19:72:@1133.4]
  wire [1:0] _T_1071; // @[Mux.scala 19:72:@1134.4]
  wire [1:0] _T_1073; // @[Mux.scala 19:72:@1135.4]
  wire [1:0] _T_1075; // @[Mux.scala 19:72:@1136.4]
  wire [1:0] _T_1077; // @[Mux.scala 19:72:@1137.4]
  wire [1:0] _T_1079; // @[Mux.scala 19:72:@1138.4]
  wire [1:0] _T_1081; // @[Mux.scala 19:72:@1139.4]
  wire [1:0] _T_1083; // @[Mux.scala 19:72:@1140.4]
  wire [1:0] _T_1085; // @[Mux.scala 19:72:@1141.4]
  wire [1:0] _T_1087; // @[Mux.scala 19:72:@1142.4]
  wire [1:0] _T_1089; // @[Mux.scala 19:72:@1143.4]
  wire [1:0] _T_1091; // @[Mux.scala 19:72:@1144.4]
  wire [1:0] _T_1093; // @[Mux.scala 19:72:@1145.4]
  wire [1:0] _T_1095; // @[Mux.scala 19:72:@1146.4]
  wire [1:0] _T_1097; // @[Mux.scala 19:72:@1147.4]
  wire [1:0] _T_1099; // @[Mux.scala 19:72:@1148.4]
  wire [1:0] _T_1101; // @[Mux.scala 19:72:@1149.4]
  wire [1:0] _T_1103; // @[Mux.scala 19:72:@1150.4]
  wire [1:0] _T_1105; // @[Mux.scala 19:72:@1151.4]
  wire [1:0] _T_1107; // @[Mux.scala 19:72:@1152.4]
  wire [1:0] _T_1109; // @[Mux.scala 19:72:@1153.4]
  wire [1:0] _T_1111; // @[Mux.scala 19:72:@1154.4]
  wire [1:0] _T_1113; // @[Mux.scala 19:72:@1155.4]
  wire [1:0] _T_1115; // @[Mux.scala 19:72:@1156.4]
  wire [1:0] _T_1117; // @[Mux.scala 19:72:@1157.4]
  wire [1:0] _T_1119; // @[Mux.scala 19:72:@1158.4]
  wire [1:0] _T_1120; // @[Mux.scala 19:72:@1159.4]
  wire [1:0] _T_1121; // @[Mux.scala 19:72:@1160.4]
  wire [1:0] _T_1122; // @[Mux.scala 19:72:@1161.4]
  wire [1:0] _T_1123; // @[Mux.scala 19:72:@1162.4]
  wire [1:0] _T_1124; // @[Mux.scala 19:72:@1163.4]
  wire [1:0] _T_1125; // @[Mux.scala 19:72:@1164.4]
  wire [1:0] _T_1126; // @[Mux.scala 19:72:@1165.4]
  wire [1:0] _T_1127; // @[Mux.scala 19:72:@1166.4]
  wire [1:0] _T_1128; // @[Mux.scala 19:72:@1167.4]
  wire [1:0] _T_1129; // @[Mux.scala 19:72:@1168.4]
  wire [1:0] _T_1130; // @[Mux.scala 19:72:@1169.4]
  wire [1:0] _T_1131; // @[Mux.scala 19:72:@1170.4]
  wire [1:0] _T_1132; // @[Mux.scala 19:72:@1171.4]
  wire [1:0] _T_1133; // @[Mux.scala 19:72:@1172.4]
  wire [1:0] _T_1134; // @[Mux.scala 19:72:@1173.4]
  wire [1:0] _T_1135; // @[Mux.scala 19:72:@1174.4]
  wire [1:0] _T_1136; // @[Mux.scala 19:72:@1175.4]
  wire [1:0] _T_1137; // @[Mux.scala 19:72:@1176.4]
  wire [1:0] _T_1138; // @[Mux.scala 19:72:@1177.4]
  wire [1:0] _T_1139; // @[Mux.scala 19:72:@1178.4]
  wire [1:0] _T_1140; // @[Mux.scala 19:72:@1179.4]
  wire [1:0] _T_1141; // @[Mux.scala 19:72:@1180.4]
  wire [1:0] _T_1142; // @[Mux.scala 19:72:@1181.4]
  wire [1:0] _T_1143; // @[Mux.scala 19:72:@1182.4]
  wire [1:0] _T_1144; // @[Mux.scala 19:72:@1183.4]
  wire [1:0] _T_1145; // @[Mux.scala 19:72:@1184.4]
  wire [1:0] _T_1146; // @[Mux.scala 19:72:@1185.4]
  wire [1:0] _T_1147; // @[Mux.scala 19:72:@1186.4]
  wire [1:0] _T_1148; // @[Mux.scala 19:72:@1187.4]
  wire [1:0] _T_1149; // @[Mux.scala 19:72:@1188.4]
  wire [1:0] _T_1150; // @[Mux.scala 19:72:@1189.4]
  wire [1:0] _T_1151; // @[Mux.scala 19:72:@1190.4]
  wire [1:0] _T_1152; // @[Mux.scala 19:72:@1191.4]
  wire [1:0] _T_1153; // @[Mux.scala 19:72:@1192.4]
  wire [1:0] _T_1154; // @[Mux.scala 19:72:@1193.4]
  wire [1:0] _T_1155; // @[Mux.scala 19:72:@1194.4]
  wire [1:0] _T_1156; // @[Mux.scala 19:72:@1195.4]
  wire [1:0] _T_1157; // @[Mux.scala 19:72:@1196.4]
  wire [1:0] _T_1158; // @[Mux.scala 19:72:@1197.4]
  wire [1:0] _T_1159; // @[Mux.scala 19:72:@1198.4]
  wire [1:0] _T_1160; // @[Mux.scala 19:72:@1199.4]
  wire [1:0] _T_1161; // @[Mux.scala 19:72:@1200.4]
  wire [1:0] _T_1162; // @[Mux.scala 19:72:@1201.4]
  wire [1:0] _T_1163; // @[Mux.scala 19:72:@1202.4]
  wire [1:0] _T_1164; // @[Mux.scala 19:72:@1203.4]
  wire [1:0] _T_1165; // @[Mux.scala 19:72:@1204.4]
  wire [1:0] _T_1166; // @[Mux.scala 19:72:@1205.4]
  wire [1:0] _T_1167; // @[Mux.scala 19:72:@1206.4]
  wire [1:0] _T_1168; // @[Mux.scala 19:72:@1207.4]
  wire [1:0] _T_1169; // @[Mux.scala 19:72:@1208.4]
  wire [1:0] _T_1170; // @[Mux.scala 19:72:@1209.4]
  wire [1:0] _T_1171; // @[Mux.scala 19:72:@1210.4]
  wire [1:0] _T_1172; // @[Mux.scala 19:72:@1211.4]
  wire [1:0] _T_1173; // @[Mux.scala 19:72:@1212.4]
  wire [1:0] _T_1174; // @[Mux.scala 19:72:@1213.4]
  wire [1:0] _T_1175; // @[Mux.scala 19:72:@1214.4]
  wire [1:0] _T_1176; // @[Mux.scala 19:72:@1215.4]
  wire [1:0] _T_1177; // @[Mux.scala 19:72:@1216.4]
  wire [1:0] _T_1178; // @[Mux.scala 19:72:@1217.4]
  wire [1:0] _T_1179; // @[Mux.scala 19:72:@1218.4]
  wire [1:0] _T_1180; // @[Mux.scala 19:72:@1219.4]
  wire [1:0] _T_1181; // @[Mux.scala 19:72:@1220.4]
  wire [1:0] predict_h_count; // @[Mux.scala 19:72:@1221.4]
  wire [9:0] _T_1186; // @[BTB.scala 107:46:@1226.4]
  wire [9:0] gshare_xor; // @[BTB.scala 107:36:@1227.4]
  reg  shift_reg; // @[BTB.scala 110:23:@1232.4]
  reg [31:0] _RAND_323;
  wire  shift_wire; // @[BTB.scala 111:30:@1233.4]
  wire  _T_1191; // @[BTB.scala 113:22:@1235.6]
  wire [8:0] _T_1192; // @[BTB.scala 114:44:@1237.8]
  wire [9:0] _T_1193; // @[Cat.scala 30:58:@1238.8]
  wire [9:0] _GEN_0; // @[BTB.scala 113:44:@1236.6]
  wire  _T_1195; // @[BTB.scala 90:30:@1247.8]
  wire  _T_1197; // @[BTB.scala 97:41:@1248.8]
  wire  _T_1198; // @[BTB.scala 97:30:@1249.8]
  wire  _T_1200; // @[BTB.scala 119:18:@1250.8]
  wire [8:0] _T_1201; // @[BTB.scala 121:35:@1253.10]
  wire [9:0] _T_1203; // @[Cat.scala 30:58:@1254.10]
  wire [1:0] predict_gshare; // @[BTB.scala 88:21:@382.4 BTB.scala 109:20:@1231.4]
  wire  _T_1210; // @[BTB.scala 95:41:@1263.12]
  wire  _T_1211; // @[BTB.scala 95:53:@1264.12]
  wire  predict_select; // @[BTB.scala 88:21:@382.4 BTB.scala 108:20:@1229.4]
  wire  _T_1212; // @[BTB.scala 95:26:@1265.12]
  wire [9:0] _T_1213; // @[Cat.scala 30:58:@1266.12]
  wire [9:0] _GEN_1; // @[BTB.scala 122:32:@1261.10]
  wire [9:0] _GEN_2; // @[BTB.scala 120:23:@1252.8]
  wire  _GEN_3; // @[BTB.scala 118:26:@1246.6]
  wire [9:0] _GEN_4; // @[BTB.scala 118:26:@1246.6]
  wire [9:0] _GEN_5; // @[BTB.scala 112:21:@1234.4]
  wire  _T_1217; // @[BTB.scala 98:44:@1271.4]
  wire  _T_1221; // @[BTB.scala 98:65:@1275.4]
  wire  _T_1222; // @[BTB.scala 98:32:@1276.4]
  wire  _T_1227; // @[BTB.scala 129:41:@1283.4]
  wire [31:0] _T_1237; // @[BTB.scala 130:8:@1291.4]
  reg  fb_reg_valid; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_324;
  reg  fb_reg_miss; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_325;
  reg  fb_reg_redirect; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_326;
  reg [1:0] fb_reg_btb_type; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_327;
  reg [31:0] fb_reg_pc; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_328;
  reg [31:0] fb_reg_tgt; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_329;
  reg  fb_reg_diff; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_330;
  reg [9:0] fb_reg_gshare; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_331;
  reg [5:0] fb_reg_lfsr; // @[BTB.scala 132:23:@1304.4]
  reg [31:0] _RAND_332;
  wire [9:0] _T_1247; // @[BTB.scala 167:57:@1313.4]
  wire [9:0] _T_1248; // @[BTB.scala 167:47:@1314.4]
  wire  _T_1249; // @[BTB.scala 146:22:@1316.4]
  wire  _T_1250; // @[BTB.scala 146:32:@1317.4]
  wire  _T_1251; // @[BTB.scala 146:26:@1318.4]
  wire [4:0] _T_1252; // @[BTB.scala 146:41:@1319.4]
  wire [5:0] _T_1253; // @[Cat.scala 30:58:@1320.4]
  wire  _T_1255; // @[BTB.scala 177:44:@1323.4]
  wire  _T_1256; // @[BTB.scala 177:44:@1324.4]
  wire  _T_1257; // @[BTB.scala 177:44:@1325.4]
  wire  _T_1258; // @[BTB.scala 177:44:@1326.4]
  wire  _T_1259; // @[BTB.scala 177:44:@1327.4]
  wire  _T_1260; // @[BTB.scala 177:44:@1328.4]
  wire  _T_1261; // @[BTB.scala 177:44:@1329.4]
  wire  _T_1262; // @[BTB.scala 177:44:@1330.4]
  wire  _T_1263; // @[BTB.scala 177:44:@1331.4]
  wire  _T_1264; // @[BTB.scala 177:44:@1332.4]
  wire  _T_1265; // @[BTB.scala 177:44:@1333.4]
  wire  _T_1266; // @[BTB.scala 177:44:@1334.4]
  wire  _T_1267; // @[BTB.scala 177:44:@1335.4]
  wire  _T_1268; // @[BTB.scala 177:44:@1336.4]
  wire  _T_1269; // @[BTB.scala 177:44:@1337.4]
  wire  _T_1270; // @[BTB.scala 177:44:@1338.4]
  wire  _T_1271; // @[BTB.scala 177:44:@1339.4]
  wire  _T_1272; // @[BTB.scala 177:44:@1340.4]
  wire  _T_1273; // @[BTB.scala 177:44:@1341.4]
  wire  _T_1274; // @[BTB.scala 177:44:@1342.4]
  wire  _T_1275; // @[BTB.scala 177:44:@1343.4]
  wire  _T_1276; // @[BTB.scala 177:44:@1344.4]
  wire  _T_1277; // @[BTB.scala 177:44:@1345.4]
  wire  _T_1278; // @[BTB.scala 177:44:@1346.4]
  wire  _T_1279; // @[BTB.scala 177:44:@1347.4]
  wire  _T_1280; // @[BTB.scala 177:44:@1348.4]
  wire  _T_1281; // @[BTB.scala 177:44:@1349.4]
  wire  _T_1282; // @[BTB.scala 177:44:@1350.4]
  wire  _T_1283; // @[BTB.scala 177:44:@1351.4]
  wire  _T_1284; // @[BTB.scala 177:44:@1352.4]
  wire  _T_1285; // @[BTB.scala 177:44:@1353.4]
  wire  _T_1286; // @[BTB.scala 177:44:@1354.4]
  wire  _T_1287; // @[BTB.scala 177:44:@1355.4]
  wire  _T_1288; // @[BTB.scala 177:44:@1356.4]
  wire  _T_1289; // @[BTB.scala 177:44:@1357.4]
  wire  _T_1290; // @[BTB.scala 177:44:@1358.4]
  wire  _T_1291; // @[BTB.scala 177:44:@1359.4]
  wire  _T_1292; // @[BTB.scala 177:44:@1360.4]
  wire  _T_1293; // @[BTB.scala 177:44:@1361.4]
  wire  _T_1294; // @[BTB.scala 177:44:@1362.4]
  wire  _T_1295; // @[BTB.scala 177:44:@1363.4]
  wire  _T_1296; // @[BTB.scala 177:44:@1364.4]
  wire  _T_1297; // @[BTB.scala 177:44:@1365.4]
  wire  _T_1298; // @[BTB.scala 177:44:@1366.4]
  wire  _T_1299; // @[BTB.scala 177:44:@1367.4]
  wire  _T_1300; // @[BTB.scala 177:44:@1368.4]
  wire  _T_1301; // @[BTB.scala 177:44:@1369.4]
  wire  _T_1302; // @[BTB.scala 177:44:@1370.4]
  wire  _T_1303; // @[BTB.scala 177:44:@1371.4]
  wire  _T_1304; // @[BTB.scala 177:44:@1372.4]
  wire  _T_1305; // @[BTB.scala 177:44:@1373.4]
  wire  _T_1306; // @[BTB.scala 177:44:@1374.4]
  wire  _T_1307; // @[BTB.scala 177:44:@1375.4]
  wire  _T_1308; // @[BTB.scala 177:44:@1376.4]
  wire  _T_1309; // @[BTB.scala 177:44:@1377.4]
  wire  _T_1310; // @[BTB.scala 177:44:@1378.4]
  wire  _T_1311; // @[BTB.scala 177:44:@1379.4]
  wire  _T_1312; // @[BTB.scala 177:44:@1380.4]
  wire  _T_1313; // @[BTB.scala 177:44:@1381.4]
  wire  _T_1314; // @[BTB.scala 177:44:@1382.4]
  wire  _T_1315; // @[BTB.scala 177:44:@1383.4]
  wire  _T_1316; // @[BTB.scala 177:44:@1384.4]
  wire  _T_1317; // @[BTB.scala 177:44:@1385.4]
  wire  _T_1318; // @[BTB.scala 177:44:@1386.4]
  wire [7:0] _T_1395; // @[BTB.scala 177:60:@1458.4]
  wire [15:0] _T_1403; // @[BTB.scala 177:60:@1466.4]
  wire [7:0] _T_1410; // @[BTB.scala 177:60:@1473.4]
  wire [31:0] _T_1419; // @[BTB.scala 177:60:@1482.4]
  wire [7:0] _T_1426; // @[BTB.scala 177:60:@1489.4]
  wire [15:0] _T_1434; // @[BTB.scala 177:60:@1497.4]
  wire [7:0] _T_1441; // @[BTB.scala 177:60:@1504.4]
  wire [31:0] _T_1450; // @[BTB.scala 177:60:@1513.4]
  wire [63:0] _T_1451; // @[BTB.scala 177:60:@1514.4]
  wire [63:0] feedback_lookup; // @[BTB.scala 177:67:@1578.4]
  wire  _T_1516; // @[Mux.scala 21:36:@1580.4]
  wire  _T_1517; // @[Mux.scala 21:36:@1581.4]
  wire  _T_1518; // @[Mux.scala 21:36:@1582.4]
  wire  _T_1519; // @[Mux.scala 21:36:@1583.4]
  wire  _T_1520; // @[Mux.scala 21:36:@1584.4]
  wire  _T_1521; // @[Mux.scala 21:36:@1585.4]
  wire  _T_1522; // @[Mux.scala 21:36:@1586.4]
  wire  _T_1523; // @[Mux.scala 21:36:@1587.4]
  wire  _T_1524; // @[Mux.scala 21:36:@1588.4]
  wire  _T_1525; // @[Mux.scala 21:36:@1589.4]
  wire  _T_1526; // @[Mux.scala 21:36:@1590.4]
  wire  _T_1527; // @[Mux.scala 21:36:@1591.4]
  wire  _T_1528; // @[Mux.scala 21:36:@1592.4]
  wire  _T_1529; // @[Mux.scala 21:36:@1593.4]
  wire  _T_1530; // @[Mux.scala 21:36:@1594.4]
  wire  _T_1531; // @[Mux.scala 21:36:@1595.4]
  wire  _T_1532; // @[Mux.scala 21:36:@1596.4]
  wire  _T_1533; // @[Mux.scala 21:36:@1597.4]
  wire  _T_1534; // @[Mux.scala 21:36:@1598.4]
  wire  _T_1535; // @[Mux.scala 21:36:@1599.4]
  wire  _T_1536; // @[Mux.scala 21:36:@1600.4]
  wire  _T_1537; // @[Mux.scala 21:36:@1601.4]
  wire  _T_1538; // @[Mux.scala 21:36:@1602.4]
  wire  _T_1539; // @[Mux.scala 21:36:@1603.4]
  wire  _T_1540; // @[Mux.scala 21:36:@1604.4]
  wire  _T_1541; // @[Mux.scala 21:36:@1605.4]
  wire  _T_1542; // @[Mux.scala 21:36:@1606.4]
  wire  _T_1543; // @[Mux.scala 21:36:@1607.4]
  wire  _T_1544; // @[Mux.scala 21:36:@1608.4]
  wire  _T_1545; // @[Mux.scala 21:36:@1609.4]
  wire  _T_1546; // @[Mux.scala 21:36:@1610.4]
  wire  _T_1547; // @[Mux.scala 21:36:@1611.4]
  wire  _T_1548; // @[Mux.scala 21:36:@1612.4]
  wire  _T_1549; // @[Mux.scala 21:36:@1613.4]
  wire  _T_1550; // @[Mux.scala 21:36:@1614.4]
  wire  _T_1551; // @[Mux.scala 21:36:@1615.4]
  wire  _T_1552; // @[Mux.scala 21:36:@1616.4]
  wire  _T_1553; // @[Mux.scala 21:36:@1617.4]
  wire  _T_1554; // @[Mux.scala 21:36:@1618.4]
  wire  _T_1555; // @[Mux.scala 21:36:@1619.4]
  wire  _T_1556; // @[Mux.scala 21:36:@1620.4]
  wire  _T_1557; // @[Mux.scala 21:36:@1621.4]
  wire  _T_1558; // @[Mux.scala 21:36:@1622.4]
  wire  _T_1559; // @[Mux.scala 21:36:@1623.4]
  wire  _T_1560; // @[Mux.scala 21:36:@1624.4]
  wire  _T_1561; // @[Mux.scala 21:36:@1625.4]
  wire  _T_1562; // @[Mux.scala 21:36:@1626.4]
  wire  _T_1563; // @[Mux.scala 21:36:@1627.4]
  wire  _T_1564; // @[Mux.scala 21:36:@1628.4]
  wire  _T_1565; // @[Mux.scala 21:36:@1629.4]
  wire  _T_1566; // @[Mux.scala 21:36:@1630.4]
  wire  _T_1567; // @[Mux.scala 21:36:@1631.4]
  wire  _T_1568; // @[Mux.scala 21:36:@1632.4]
  wire  _T_1569; // @[Mux.scala 21:36:@1633.4]
  wire  _T_1570; // @[Mux.scala 21:36:@1634.4]
  wire  _T_1571; // @[Mux.scala 21:36:@1635.4]
  wire  _T_1572; // @[Mux.scala 21:36:@1636.4]
  wire  _T_1573; // @[Mux.scala 21:36:@1637.4]
  wire  _T_1574; // @[Mux.scala 21:36:@1638.4]
  wire  _T_1575; // @[Mux.scala 21:36:@1639.4]
  wire  _T_1576; // @[Mux.scala 21:36:@1640.4]
  wire  _T_1577; // @[Mux.scala 21:36:@1641.4]
  wire  _T_1578; // @[Mux.scala 21:36:@1642.4]
  wire  _T_1579; // @[Mux.scala 21:36:@1643.4]
  wire [1:0] _T_1582; // @[Mux.scala 19:72:@1644.4]
  wire [1:0] _T_1584; // @[Mux.scala 19:72:@1645.4]
  wire [1:0] _T_1586; // @[Mux.scala 19:72:@1646.4]
  wire [1:0] _T_1588; // @[Mux.scala 19:72:@1647.4]
  wire [1:0] _T_1590; // @[Mux.scala 19:72:@1648.4]
  wire [1:0] _T_1592; // @[Mux.scala 19:72:@1649.4]
  wire [1:0] _T_1594; // @[Mux.scala 19:72:@1650.4]
  wire [1:0] _T_1596; // @[Mux.scala 19:72:@1651.4]
  wire [1:0] _T_1598; // @[Mux.scala 19:72:@1652.4]
  wire [1:0] _T_1600; // @[Mux.scala 19:72:@1653.4]
  wire [1:0] _T_1602; // @[Mux.scala 19:72:@1654.4]
  wire [1:0] _T_1604; // @[Mux.scala 19:72:@1655.4]
  wire [1:0] _T_1606; // @[Mux.scala 19:72:@1656.4]
  wire [1:0] _T_1608; // @[Mux.scala 19:72:@1657.4]
  wire [1:0] _T_1610; // @[Mux.scala 19:72:@1658.4]
  wire [1:0] _T_1612; // @[Mux.scala 19:72:@1659.4]
  wire [1:0] _T_1614; // @[Mux.scala 19:72:@1660.4]
  wire [1:0] _T_1616; // @[Mux.scala 19:72:@1661.4]
  wire [1:0] _T_1618; // @[Mux.scala 19:72:@1662.4]
  wire [1:0] _T_1620; // @[Mux.scala 19:72:@1663.4]
  wire [1:0] _T_1622; // @[Mux.scala 19:72:@1664.4]
  wire [1:0] _T_1624; // @[Mux.scala 19:72:@1665.4]
  wire [1:0] _T_1626; // @[Mux.scala 19:72:@1666.4]
  wire [1:0] _T_1628; // @[Mux.scala 19:72:@1667.4]
  wire [1:0] _T_1630; // @[Mux.scala 19:72:@1668.4]
  wire [1:0] _T_1632; // @[Mux.scala 19:72:@1669.4]
  wire [1:0] _T_1634; // @[Mux.scala 19:72:@1670.4]
  wire [1:0] _T_1636; // @[Mux.scala 19:72:@1671.4]
  wire [1:0] _T_1638; // @[Mux.scala 19:72:@1672.4]
  wire [1:0] _T_1640; // @[Mux.scala 19:72:@1673.4]
  wire [1:0] _T_1642; // @[Mux.scala 19:72:@1674.4]
  wire [1:0] _T_1644; // @[Mux.scala 19:72:@1675.4]
  wire [1:0] _T_1646; // @[Mux.scala 19:72:@1676.4]
  wire [1:0] _T_1648; // @[Mux.scala 19:72:@1677.4]
  wire [1:0] _T_1650; // @[Mux.scala 19:72:@1678.4]
  wire [1:0] _T_1652; // @[Mux.scala 19:72:@1679.4]
  wire [1:0] _T_1654; // @[Mux.scala 19:72:@1680.4]
  wire [1:0] _T_1656; // @[Mux.scala 19:72:@1681.4]
  wire [1:0] _T_1658; // @[Mux.scala 19:72:@1682.4]
  wire [1:0] _T_1660; // @[Mux.scala 19:72:@1683.4]
  wire [1:0] _T_1662; // @[Mux.scala 19:72:@1684.4]
  wire [1:0] _T_1664; // @[Mux.scala 19:72:@1685.4]
  wire [1:0] _T_1666; // @[Mux.scala 19:72:@1686.4]
  wire [1:0] _T_1668; // @[Mux.scala 19:72:@1687.4]
  wire [1:0] _T_1670; // @[Mux.scala 19:72:@1688.4]
  wire [1:0] _T_1672; // @[Mux.scala 19:72:@1689.4]
  wire [1:0] _T_1674; // @[Mux.scala 19:72:@1690.4]
  wire [1:0] _T_1676; // @[Mux.scala 19:72:@1691.4]
  wire [1:0] _T_1678; // @[Mux.scala 19:72:@1692.4]
  wire [1:0] _T_1680; // @[Mux.scala 19:72:@1693.4]
  wire [1:0] _T_1682; // @[Mux.scala 19:72:@1694.4]
  wire [1:0] _T_1684; // @[Mux.scala 19:72:@1695.4]
  wire [1:0] _T_1686; // @[Mux.scala 19:72:@1696.4]
  wire [1:0] _T_1688; // @[Mux.scala 19:72:@1697.4]
  wire [1:0] _T_1690; // @[Mux.scala 19:72:@1698.4]
  wire [1:0] _T_1692; // @[Mux.scala 19:72:@1699.4]
  wire [1:0] _T_1694; // @[Mux.scala 19:72:@1700.4]
  wire [1:0] _T_1696; // @[Mux.scala 19:72:@1701.4]
  wire [1:0] _T_1698; // @[Mux.scala 19:72:@1702.4]
  wire [1:0] _T_1700; // @[Mux.scala 19:72:@1703.4]
  wire [1:0] _T_1702; // @[Mux.scala 19:72:@1704.4]
  wire [1:0] _T_1704; // @[Mux.scala 19:72:@1705.4]
  wire [1:0] _T_1706; // @[Mux.scala 19:72:@1706.4]
  wire [1:0] _T_1708; // @[Mux.scala 19:72:@1707.4]
  wire [1:0] _T_1709; // @[Mux.scala 19:72:@1708.4]
  wire [1:0] _T_1710; // @[Mux.scala 19:72:@1709.4]
  wire [1:0] _T_1711; // @[Mux.scala 19:72:@1710.4]
  wire [1:0] _T_1712; // @[Mux.scala 19:72:@1711.4]
  wire [1:0] _T_1713; // @[Mux.scala 19:72:@1712.4]
  wire [1:0] _T_1714; // @[Mux.scala 19:72:@1713.4]
  wire [1:0] _T_1715; // @[Mux.scala 19:72:@1714.4]
  wire [1:0] _T_1716; // @[Mux.scala 19:72:@1715.4]
  wire [1:0] _T_1717; // @[Mux.scala 19:72:@1716.4]
  wire [1:0] _T_1718; // @[Mux.scala 19:72:@1717.4]
  wire [1:0] _T_1719; // @[Mux.scala 19:72:@1718.4]
  wire [1:0] _T_1720; // @[Mux.scala 19:72:@1719.4]
  wire [1:0] _T_1721; // @[Mux.scala 19:72:@1720.4]
  wire [1:0] _T_1722; // @[Mux.scala 19:72:@1721.4]
  wire [1:0] _T_1723; // @[Mux.scala 19:72:@1722.4]
  wire [1:0] _T_1724; // @[Mux.scala 19:72:@1723.4]
  wire [1:0] _T_1725; // @[Mux.scala 19:72:@1724.4]
  wire [1:0] _T_1726; // @[Mux.scala 19:72:@1725.4]
  wire [1:0] _T_1727; // @[Mux.scala 19:72:@1726.4]
  wire [1:0] _T_1728; // @[Mux.scala 19:72:@1727.4]
  wire [1:0] _T_1729; // @[Mux.scala 19:72:@1728.4]
  wire [1:0] _T_1730; // @[Mux.scala 19:72:@1729.4]
  wire [1:0] _T_1731; // @[Mux.scala 19:72:@1730.4]
  wire [1:0] _T_1732; // @[Mux.scala 19:72:@1731.4]
  wire [1:0] _T_1733; // @[Mux.scala 19:72:@1732.4]
  wire [1:0] _T_1734; // @[Mux.scala 19:72:@1733.4]
  wire [1:0] _T_1735; // @[Mux.scala 19:72:@1734.4]
  wire [1:0] _T_1736; // @[Mux.scala 19:72:@1735.4]
  wire [1:0] _T_1737; // @[Mux.scala 19:72:@1736.4]
  wire [1:0] _T_1738; // @[Mux.scala 19:72:@1737.4]
  wire [1:0] _T_1739; // @[Mux.scala 19:72:@1738.4]
  wire [1:0] _T_1740; // @[Mux.scala 19:72:@1739.4]
  wire [1:0] _T_1741; // @[Mux.scala 19:72:@1740.4]
  wire [1:0] _T_1742; // @[Mux.scala 19:72:@1741.4]
  wire [1:0] _T_1743; // @[Mux.scala 19:72:@1742.4]
  wire [1:0] _T_1744; // @[Mux.scala 19:72:@1743.4]
  wire [1:0] _T_1745; // @[Mux.scala 19:72:@1744.4]
  wire [1:0] _T_1746; // @[Mux.scala 19:72:@1745.4]
  wire [1:0] _T_1747; // @[Mux.scala 19:72:@1746.4]
  wire [1:0] _T_1748; // @[Mux.scala 19:72:@1747.4]
  wire [1:0] _T_1749; // @[Mux.scala 19:72:@1748.4]
  wire [1:0] _T_1750; // @[Mux.scala 19:72:@1749.4]
  wire [1:0] _T_1751; // @[Mux.scala 19:72:@1750.4]
  wire [1:0] _T_1752; // @[Mux.scala 19:72:@1751.4]
  wire [1:0] _T_1753; // @[Mux.scala 19:72:@1752.4]
  wire [1:0] _T_1754; // @[Mux.scala 19:72:@1753.4]
  wire [1:0] _T_1755; // @[Mux.scala 19:72:@1754.4]
  wire [1:0] _T_1756; // @[Mux.scala 19:72:@1755.4]
  wire [1:0] _T_1757; // @[Mux.scala 19:72:@1756.4]
  wire [1:0] _T_1758; // @[Mux.scala 19:72:@1757.4]
  wire [1:0] _T_1759; // @[Mux.scala 19:72:@1758.4]
  wire [1:0] _T_1760; // @[Mux.scala 19:72:@1759.4]
  wire [1:0] _T_1761; // @[Mux.scala 19:72:@1760.4]
  wire [1:0] _T_1762; // @[Mux.scala 19:72:@1761.4]
  wire [1:0] _T_1763; // @[Mux.scala 19:72:@1762.4]
  wire [1:0] _T_1764; // @[Mux.scala 19:72:@1763.4]
  wire [1:0] _T_1765; // @[Mux.scala 19:72:@1764.4]
  wire [1:0] _T_1766; // @[Mux.scala 19:72:@1765.4]
  wire [1:0] _T_1767; // @[Mux.scala 19:72:@1766.4]
  wire [1:0] _T_1768; // @[Mux.scala 19:72:@1767.4]
  wire [1:0] _T_1769; // @[Mux.scala 19:72:@1768.4]
  wire [1:0] _T_1770; // @[Mux.scala 19:72:@1769.4]
  wire [1:0] feedback_h_count; // @[Mux.scala 19:72:@1770.4]
  wire  _T_1776; // @[BTB.scala 172:30:@1776.4]
  wire [31:0] _T_1777; // @[OneHot.scala 26:18:@1777.4]
  wire [31:0] _T_1778; // @[OneHot.scala 27:18:@1778.4]
  wire  _T_1780; // @[OneHot.scala 28:14:@1779.4]
  wire [31:0] _T_1781; // @[OneHot.scala 28:28:@1780.4]
  wire [15:0] _T_1782; // @[OneHot.scala 26:18:@1781.4]
  wire [15:0] _T_1783; // @[OneHot.scala 27:18:@1782.4]
  wire  _T_1785; // @[OneHot.scala 28:14:@1783.4]
  wire [15:0] _T_1786; // @[OneHot.scala 28:28:@1784.4]
  wire [7:0] _T_1787; // @[OneHot.scala 26:18:@1785.4]
  wire [7:0] _T_1788; // @[OneHot.scala 27:18:@1786.4]
  wire  _T_1790; // @[OneHot.scala 28:14:@1787.4]
  wire [7:0] _T_1791; // @[OneHot.scala 28:28:@1788.4]
  wire [3:0] _T_1792; // @[OneHot.scala 26:18:@1789.4]
  wire [3:0] _T_1793; // @[OneHot.scala 27:18:@1790.4]
  wire  _T_1795; // @[OneHot.scala 28:14:@1791.4]
  wire [3:0] _T_1796; // @[OneHot.scala 28:28:@1792.4]
  wire [1:0] _T_1797; // @[OneHot.scala 26:18:@1793.4]
  wire [1:0] _T_1798; // @[OneHot.scala 27:18:@1794.4]
  wire  _T_1800; // @[OneHot.scala 28:14:@1795.4]
  wire [1:0] _T_1801; // @[OneHot.scala 28:28:@1796.4]
  wire  _T_1802; // @[CircuitMath.scala 30:8:@1797.4]
  wire [5:0] _T_1807; // @[Cat.scala 30:58:@1802.4]
  wire [63:0] _T_1871; // @[BTB.scala 181:26:@1866.4]
  wire  _T_1873; // @[BTB.scala 181:26:@1867.4]
  wire  _T_1938; // @[OneHot.scala 39:40:@1932.4]
  wire  _T_1939; // @[OneHot.scala 39:40:@1933.4]
  wire  _T_1940; // @[OneHot.scala 39:40:@1934.4]
  wire  _T_1941; // @[OneHot.scala 39:40:@1935.4]
  wire  _T_1942; // @[OneHot.scala 39:40:@1936.4]
  wire  _T_1943; // @[OneHot.scala 39:40:@1937.4]
  wire  _T_1944; // @[OneHot.scala 39:40:@1938.4]
  wire  _T_1945; // @[OneHot.scala 39:40:@1939.4]
  wire  _T_1946; // @[OneHot.scala 39:40:@1940.4]
  wire  _T_1947; // @[OneHot.scala 39:40:@1941.4]
  wire  _T_1948; // @[OneHot.scala 39:40:@1942.4]
  wire  _T_1949; // @[OneHot.scala 39:40:@1943.4]
  wire  _T_1950; // @[OneHot.scala 39:40:@1944.4]
  wire  _T_1951; // @[OneHot.scala 39:40:@1945.4]
  wire  _T_1952; // @[OneHot.scala 39:40:@1946.4]
  wire  _T_1953; // @[OneHot.scala 39:40:@1947.4]
  wire  _T_1954; // @[OneHot.scala 39:40:@1948.4]
  wire  _T_1955; // @[OneHot.scala 39:40:@1949.4]
  wire  _T_1956; // @[OneHot.scala 39:40:@1950.4]
  wire  _T_1957; // @[OneHot.scala 39:40:@1951.4]
  wire  _T_1958; // @[OneHot.scala 39:40:@1952.4]
  wire  _T_1959; // @[OneHot.scala 39:40:@1953.4]
  wire  _T_1960; // @[OneHot.scala 39:40:@1954.4]
  wire  _T_1961; // @[OneHot.scala 39:40:@1955.4]
  wire  _T_1962; // @[OneHot.scala 39:40:@1956.4]
  wire  _T_1963; // @[OneHot.scala 39:40:@1957.4]
  wire  _T_1964; // @[OneHot.scala 39:40:@1958.4]
  wire  _T_1965; // @[OneHot.scala 39:40:@1959.4]
  wire  _T_1966; // @[OneHot.scala 39:40:@1960.4]
  wire  _T_1967; // @[OneHot.scala 39:40:@1961.4]
  wire  _T_1968; // @[OneHot.scala 39:40:@1962.4]
  wire  _T_1969; // @[OneHot.scala 39:40:@1963.4]
  wire  _T_1970; // @[OneHot.scala 39:40:@1964.4]
  wire  _T_1971; // @[OneHot.scala 39:40:@1965.4]
  wire  _T_1972; // @[OneHot.scala 39:40:@1966.4]
  wire  _T_1973; // @[OneHot.scala 39:40:@1967.4]
  wire  _T_1974; // @[OneHot.scala 39:40:@1968.4]
  wire  _T_1975; // @[OneHot.scala 39:40:@1969.4]
  wire  _T_1976; // @[OneHot.scala 39:40:@1970.4]
  wire  _T_1977; // @[OneHot.scala 39:40:@1971.4]
  wire  _T_1978; // @[OneHot.scala 39:40:@1972.4]
  wire  _T_1979; // @[OneHot.scala 39:40:@1973.4]
  wire  _T_1980; // @[OneHot.scala 39:40:@1974.4]
  wire  _T_1981; // @[OneHot.scala 39:40:@1975.4]
  wire  _T_1982; // @[OneHot.scala 39:40:@1976.4]
  wire  _T_1983; // @[OneHot.scala 39:40:@1977.4]
  wire  _T_1984; // @[OneHot.scala 39:40:@1978.4]
  wire  _T_1985; // @[OneHot.scala 39:40:@1979.4]
  wire  _T_1986; // @[OneHot.scala 39:40:@1980.4]
  wire  _T_1987; // @[OneHot.scala 39:40:@1981.4]
  wire  _T_1988; // @[OneHot.scala 39:40:@1982.4]
  wire  _T_1989; // @[OneHot.scala 39:40:@1983.4]
  wire  _T_1990; // @[OneHot.scala 39:40:@1984.4]
  wire  _T_1991; // @[OneHot.scala 39:40:@1985.4]
  wire  _T_1992; // @[OneHot.scala 39:40:@1986.4]
  wire  _T_1993; // @[OneHot.scala 39:40:@1987.4]
  wire  _T_1994; // @[OneHot.scala 39:40:@1988.4]
  wire  _T_1995; // @[OneHot.scala 39:40:@1989.4]
  wire  _T_1996; // @[OneHot.scala 39:40:@1990.4]
  wire  _T_1997; // @[OneHot.scala 39:40:@1991.4]
  wire  _T_1998; // @[OneHot.scala 39:40:@1992.4]
  wire  _T_1999; // @[OneHot.scala 39:40:@1993.4]
  wire  _T_2000; // @[OneHot.scala 39:40:@1994.4]
  wire [5:0] _T_2066; // @[Mux.scala 31:69:@1996.4]
  wire [5:0] _T_2067; // @[Mux.scala 31:69:@1997.4]
  wire [5:0] _T_2068; // @[Mux.scala 31:69:@1998.4]
  wire [5:0] _T_2069; // @[Mux.scala 31:69:@1999.4]
  wire [5:0] _T_2070; // @[Mux.scala 31:69:@2000.4]
  wire [5:0] _T_2071; // @[Mux.scala 31:69:@2001.4]
  wire [5:0] _T_2072; // @[Mux.scala 31:69:@2002.4]
  wire [5:0] _T_2073; // @[Mux.scala 31:69:@2003.4]
  wire [5:0] _T_2074; // @[Mux.scala 31:69:@2004.4]
  wire [5:0] _T_2075; // @[Mux.scala 31:69:@2005.4]
  wire [5:0] _T_2076; // @[Mux.scala 31:69:@2006.4]
  wire [5:0] _T_2077; // @[Mux.scala 31:69:@2007.4]
  wire [5:0] _T_2078; // @[Mux.scala 31:69:@2008.4]
  wire [5:0] _T_2079; // @[Mux.scala 31:69:@2009.4]
  wire [5:0] _T_2080; // @[Mux.scala 31:69:@2010.4]
  wire [5:0] _T_2081; // @[Mux.scala 31:69:@2011.4]
  wire [5:0] _T_2082; // @[Mux.scala 31:69:@2012.4]
  wire [5:0] _T_2083; // @[Mux.scala 31:69:@2013.4]
  wire [5:0] _T_2084; // @[Mux.scala 31:69:@2014.4]
  wire [5:0] _T_2085; // @[Mux.scala 31:69:@2015.4]
  wire [5:0] _T_2086; // @[Mux.scala 31:69:@2016.4]
  wire [5:0] _T_2087; // @[Mux.scala 31:69:@2017.4]
  wire [5:0] _T_2088; // @[Mux.scala 31:69:@2018.4]
  wire [5:0] _T_2089; // @[Mux.scala 31:69:@2019.4]
  wire [5:0] _T_2090; // @[Mux.scala 31:69:@2020.4]
  wire [5:0] _T_2091; // @[Mux.scala 31:69:@2021.4]
  wire [5:0] _T_2092; // @[Mux.scala 31:69:@2022.4]
  wire [5:0] _T_2093; // @[Mux.scala 31:69:@2023.4]
  wire [5:0] _T_2094; // @[Mux.scala 31:69:@2024.4]
  wire [5:0] _T_2095; // @[Mux.scala 31:69:@2025.4]
  wire [5:0] _T_2096; // @[Mux.scala 31:69:@2026.4]
  wire [5:0] _T_2097; // @[Mux.scala 31:69:@2027.4]
  wire [5:0] _T_2098; // @[Mux.scala 31:69:@2028.4]
  wire [5:0] _T_2099; // @[Mux.scala 31:69:@2029.4]
  wire [5:0] _T_2100; // @[Mux.scala 31:69:@2030.4]
  wire [5:0] _T_2101; // @[Mux.scala 31:69:@2031.4]
  wire [5:0] _T_2102; // @[Mux.scala 31:69:@2032.4]
  wire [5:0] _T_2103; // @[Mux.scala 31:69:@2033.4]
  wire [5:0] _T_2104; // @[Mux.scala 31:69:@2034.4]
  wire [5:0] _T_2105; // @[Mux.scala 31:69:@2035.4]
  wire [5:0] _T_2106; // @[Mux.scala 31:69:@2036.4]
  wire [5:0] _T_2107; // @[Mux.scala 31:69:@2037.4]
  wire [5:0] _T_2108; // @[Mux.scala 31:69:@2038.4]
  wire [5:0] _T_2109; // @[Mux.scala 31:69:@2039.4]
  wire [5:0] _T_2110; // @[Mux.scala 31:69:@2040.4]
  wire [5:0] _T_2111; // @[Mux.scala 31:69:@2041.4]
  wire [5:0] _T_2112; // @[Mux.scala 31:69:@2042.4]
  wire [5:0] _T_2113; // @[Mux.scala 31:69:@2043.4]
  wire [5:0] _T_2114; // @[Mux.scala 31:69:@2044.4]
  wire [5:0] _T_2115; // @[Mux.scala 31:69:@2045.4]
  wire [5:0] _T_2116; // @[Mux.scala 31:69:@2046.4]
  wire [5:0] _T_2117; // @[Mux.scala 31:69:@2047.4]
  wire [5:0] _T_2118; // @[Mux.scala 31:69:@2048.4]
  wire [5:0] _T_2119; // @[Mux.scala 31:69:@2049.4]
  wire [5:0] _T_2120; // @[Mux.scala 31:69:@2050.4]
  wire [5:0] _T_2121; // @[Mux.scala 31:69:@2051.4]
  wire [5:0] _T_2122; // @[Mux.scala 31:69:@2052.4]
  wire [5:0] _T_2123; // @[Mux.scala 31:69:@2053.4]
  wire [5:0] _T_2124; // @[Mux.scala 31:69:@2054.4]
  wire [5:0] _T_2125; // @[Mux.scala 31:69:@2055.4]
  wire [5:0] _T_2126; // @[Mux.scala 31:69:@2056.4]
  wire [5:0] _T_2127; // @[Mux.scala 31:69:@2057.4]
  wire [5:0] _T_2128; // @[Mux.scala 31:69:@2058.4]
  wire [5:0] _T_2129; // @[BTB.scala 181:8:@2059.4]
  wire [5:0] feedback_idx; // @[BTB.scala 180:22:@2060.4]
  wire  _GEN_7; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_8; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_9; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_10; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_11; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_12; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_13; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_14; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_15; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_16; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_17; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_18; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_19; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_20; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_21; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_22; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_23; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_24; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_25; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_26; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_27; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_28; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_29; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_30; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_31; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_32; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_33; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_34; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_35; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_36; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_37; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_38; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_39; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_40; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_41; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_42; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_43; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_44; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_45; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_46; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_47; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_48; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_49; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_50; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_51; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_52; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_53; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_54; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_55; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_56; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_57; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_58; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_59; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_60; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_61; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_62; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_63; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_64; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_65; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_66; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_67; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_68; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_69; // @[BTB.scala 185:32:@2064.8]
  wire  _GEN_70; // @[BTB.scala 185:32:@2064.8]
  wire  _T_2135; // @[BTB.scala 187:51:@2069.10]
  wire  _GEN_71; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_72; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_73; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_74; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_75; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_76; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_77; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_78; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_79; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_80; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_81; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_82; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_83; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_84; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_85; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_86; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_87; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_88; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_89; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_90; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_91; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_92; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_93; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_94; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_95; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_96; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_97; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_98; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_99; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_100; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_101; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_102; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_103; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_104; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_105; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_106; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_107; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_108; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_109; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_110; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_111; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_112; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_113; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_114; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_115; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_116; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_117; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_118; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_119; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_120; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_121; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_122; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_123; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_124; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_125; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_126; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_127; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_128; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_129; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_130; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_131; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_132; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_133; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_134; // @[BTB.scala 187:32:@2070.10]
  wire  _GEN_135; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_136; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_137; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_138; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_139; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_140; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_141; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_142; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_143; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_144; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_145; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_146; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_147; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_148; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_149; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_150; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_151; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_152; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_153; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_154; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_155; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_156; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_157; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_158; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_159; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_160; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_161; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_162; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_163; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_164; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_165; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_166; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_167; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_168; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_169; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_170; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_171; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_172; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_173; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_174; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_175; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_176; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_177; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_178; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_179; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_180; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_181; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_182; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_183; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_184; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_185; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_186; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_187; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_188; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_189; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_190; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_191; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_192; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_193; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_194; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_195; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_196; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_197; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_198; // @[BTB.scala 186:32:@2068.8]
  wire  _GEN_199; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_200; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_201; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_202; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_203; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_204; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_205; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_206; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_207; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_208; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_209; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_210; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_211; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_212; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_213; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_214; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_215; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_216; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_217; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_218; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_219; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_220; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_221; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_222; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_223; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_224; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_225; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_226; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_227; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_228; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_229; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_230; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_231; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_232; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_233; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_234; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_235; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_236; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_237; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_238; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_239; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_240; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_241; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_242; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_243; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_244; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_245; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_246; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_247; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_248; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_249; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_250; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_251; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_252; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_253; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_254; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_255; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_256; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_257; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_258; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_259; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_260; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_261; // @[BTB.scala 184:28:@2063.6]
  wire  _GEN_262; // @[BTB.scala 184:28:@2063.6]
  wire [31:0] _GEN_263; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_264; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_265; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_266; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_267; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_268; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_269; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_270; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_271; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_272; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_273; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_274; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_275; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_276; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_277; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_278; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_279; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_280; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_281; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_282; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_283; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_284; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_285; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_286; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_287; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_288; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_289; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_290; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_291; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_292; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_293; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_294; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_295; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_296; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_297; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_298; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_299; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_300; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_301; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_302; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_303; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_304; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_305; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_306; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_307; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_308; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_309; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_310; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_311; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_312; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_313; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_314; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_315; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_316; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_317; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_318; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_319; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_320; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_321; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_322; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_323; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_324; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_325; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_326; // @[BTB.scala 190:33:@2073.8]
  wire [31:0] _GEN_327; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_328; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_329; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_330; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_331; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_332; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_333; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_334; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_335; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_336; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_337; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_338; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_339; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_340; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_341; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_342; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_343; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_344; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_345; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_346; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_347; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_348; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_349; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_350; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_351; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_352; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_353; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_354; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_355; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_356; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_357; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_358; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_359; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_360; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_361; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_362; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_363; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_364; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_365; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_366; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_367; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_368; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_369; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_370; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_371; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_372; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_373; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_374; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_375; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_376; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_377; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_378; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_379; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_380; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_381; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_382; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_383; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_384; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_385; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_386; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_387; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_388; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_389; // @[BTB.scala 191:33:@2074.8]
  wire [31:0] _GEN_390; // @[BTB.scala 191:33:@2074.8]
  wire [1:0] _GEN_391; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_392; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_393; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_394; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_395; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_396; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_397; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_398; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_399; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_400; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_401; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_402; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_403; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_404; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_405; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_406; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_407; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_408; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_409; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_410; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_411; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_412; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_413; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_414; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_415; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_416; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_417; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_418; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_419; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_420; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_421; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_422; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_423; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_424; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_425; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_426; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_427; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_428; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_429; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_430; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_431; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_432; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_433; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_434; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_435; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_436; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_437; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_438; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_439; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_440; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_441; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_442; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_443; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_444; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_445; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_446; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_447; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_448; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_449; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_450; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_451; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_452; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_453; // @[BTB.scala 192:33:@2075.8]
  wire [1:0] _GEN_454; // @[BTB.scala 192:33:@2075.8]
  wire [31:0] _GEN_455; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_456; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_457; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_458; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_459; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_460; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_461; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_462; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_463; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_464; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_465; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_466; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_467; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_468; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_469; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_470; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_471; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_472; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_473; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_474; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_475; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_476; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_477; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_478; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_479; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_480; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_481; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_482; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_483; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_484; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_485; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_486; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_487; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_488; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_489; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_490; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_491; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_492; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_493; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_494; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_495; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_496; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_497; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_498; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_499; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_500; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_501; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_502; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_503; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_504; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_505; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_506; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_507; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_508; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_509; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_510; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_511; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_512; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_513; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_514; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_515; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_516; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_517; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_518; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_519; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_520; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_521; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_522; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_523; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_524; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_525; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_526; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_527; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_528; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_529; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_530; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_531; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_532; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_533; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_534; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_535; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_536; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_537; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_538; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_539; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_540; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_541; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_542; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_543; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_544; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_545; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_546; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_547; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_548; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_549; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_550; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_551; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_552; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_553; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_554; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_555; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_556; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_557; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_558; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_559; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_560; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_561; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_562; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_563; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_564; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_565; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_566; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_567; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_568; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_569; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_570; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_571; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_572; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_573; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_574; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_575; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_576; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_577; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_578; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_579; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_580; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_581; // @[BTB.scala 189:28:@2072.6]
  wire [31:0] _GEN_582; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_583; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_584; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_585; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_586; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_587; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_588; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_589; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_590; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_591; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_592; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_593; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_594; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_595; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_596; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_597; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_598; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_599; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_600; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_601; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_602; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_603; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_604; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_605; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_606; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_607; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_608; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_609; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_610; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_611; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_612; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_613; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_614; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_615; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_616; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_617; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_618; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_619; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_620; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_621; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_622; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_623; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_624; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_625; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_626; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_627; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_628; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_629; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_630; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_631; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_632; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_633; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_634; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_635; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_636; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_637; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_638; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_639; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_640; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_641; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_642; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_643; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_644; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_645; // @[BTB.scala 189:28:@2072.6]
  wire [1:0] _GEN_646; // @[BTB.scala 189:28:@2072.6]
  wire  _T_2141; // @[BTB.scala 62:38:@2082.12]
  wire  _T_2142; // @[BTB.scala 62:45:@2083.12]
  wire  _T_2143; // @[BTB.scala 62:54:@2084.12]
  wire  _T_2145; // @[BTB.scala 62:52:@2085.12]
  wire  _T_2146; // @[BTB.scala 62:49:@2086.12]
  wire [1:0] _T_2147; // @[Cat.scala 30:58:@2087.12]
  wire [1:0] _GEN_647; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_648; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_649; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_650; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_651; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_652; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_653; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_654; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_655; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_656; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_657; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_658; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_659; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_660; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_661; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_662; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_663; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_664; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_665; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_666; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_667; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_668; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_669; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_670; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_671; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_672; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_673; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_674; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_675; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_676; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_677; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_678; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_679; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_680; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_681; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_682; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_683; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_684; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_685; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_686; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_687; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_688; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_689; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_690; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_691; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_692; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_693; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_694; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_695; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_696; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_697; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_698; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_699; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_700; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_701; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_702; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_703; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_704; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_705; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_706; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_707; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_708; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_709; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] _GEN_710; // @[BTB.scala 198:37:@2088.12]
  wire [1:0] feedback_gshare; // @[BTB.scala 170:22:@1322.4 BTB.scala 179:20:@1775.4]
  wire  _T_2150; // @[BTB.scala 62:38:@2090.12]
  wire  _T_2151; // @[BTB.scala 62:45:@2091.12]
  wire  _T_2152; // @[BTB.scala 62:54:@2092.12]
  wire  _T_2154; // @[BTB.scala 62:52:@2093.12]
  wire  _T_2155; // @[BTB.scala 62:49:@2094.12]
  wire [1:0] _T_2157; // @[BTB.scala 64:38:@2099.12]
  wire  _T_2159; // @[BTB.scala 64:38:@2100.12]
  wire  _T_2164; // @[BTB.scala 64:49:@2104.12]
  wire [1:0] _T_2165; // @[Cat.scala 30:58:@2105.12]
  wire [1:0] _GEN_711; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_712; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_713; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_714; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_715; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_716; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_717; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_718; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_719; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_720; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_721; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_722; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_723; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_724; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_725; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_726; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_727; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_728; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_729; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_730; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_731; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_732; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_733; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_734; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_735; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_736; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_737; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_738; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_739; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_740; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_741; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_742; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_743; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_744; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_745; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_746; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_747; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_748; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_749; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_750; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_751; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_752; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_753; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_754; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_755; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_756; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_757; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_758; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_759; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_760; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_761; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_762; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_763; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_764; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_765; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_766; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_767; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_768; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_769; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_770; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_771; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_772; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_773; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _GEN_774; // @[BTB.scala 201:37:@2106.12]
  wire [1:0] _T_2167; // @[BTB.scala 64:38:@2108.12]
  wire  _T_2169; // @[BTB.scala 64:38:@2109.12]
  wire  _T_2174; // @[BTB.scala 64:49:@2113.12]
  wire [1:0] _GEN_775; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_776; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_777; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_778; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_779; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_780; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_781; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_782; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_783; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_784; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_785; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_786; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_787; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_788; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_789; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_790; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_791; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_792; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_793; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_794; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_795; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_796; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_797; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_798; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_799; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_800; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_801; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_802; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_803; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_804; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_805; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_806; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_807; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_808; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_809; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_810; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_811; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_812; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_813; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_814; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_815; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_816; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_817; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_818; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_819; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_820; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_821; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_822; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_823; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_824; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_825; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_826; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_827; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_828; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_829; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_830; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_831; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_832; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_833; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_834; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_835; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_836; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_837; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_838; // @[BTB.scala 197:32:@2081.10]
  wire  _GEN_846; // @[BTB.scala 197:32:@2081.10]
  wire [1:0] _GEN_849; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_850; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_851; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_852; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_853; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_854; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_855; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_856; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_857; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_858; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_859; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_860; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_861; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_862; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_863; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_864; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_865; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_866; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_867; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_868; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_869; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_870; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_871; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_872; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_873; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_874; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_875; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_876; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_877; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_878; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_879; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_880; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_881; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_882; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_883; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_884; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_885; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_886; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_887; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_888; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_889; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_890; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_891; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_892; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_893; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_894; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_895; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_896; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_897; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_898; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_899; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_900; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_901; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_902; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_903; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_904; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_905; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_906; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_907; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_908; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_909; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_910; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_911; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_912; // @[BTB.scala 205:35:@2120.12]
  wire [1:0] _GEN_913; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_914; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_915; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_916; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_917; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_918; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_919; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_920; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_921; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_922; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_923; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_924; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_925; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_926; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_927; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_928; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_929; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_930; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_931; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_932; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_933; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_934; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_935; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_936; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_937; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_938; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_939; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_940; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_941; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_942; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_943; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_944; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_945; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_946; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_947; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_948; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_949; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_950; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_951; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_952; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_953; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_954; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_955; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_956; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_957; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_958; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_959; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_960; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_961; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_962; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_963; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_964; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_965; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_966; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_967; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_968; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_969; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_970; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_971; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_972; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_973; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_974; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_975; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_976; // @[BTB.scala 204:35:@2119.10]
  wire [1:0] _GEN_978; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_979; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_980; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_981; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_982; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_983; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_984; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_985; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_986; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_987; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_988; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_989; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_990; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_991; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_992; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_993; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_994; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_995; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_996; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_997; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_998; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_999; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1000; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1001; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1002; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1003; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1004; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1005; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1006; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1007; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1008; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1009; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1010; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1011; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1012; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1013; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1014; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1015; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1016; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1017; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1018; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1019; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1020; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1021; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1022; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1023; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1024; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1025; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1026; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1027; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1028; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1029; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1030; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1031; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1032; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1033; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1034; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1035; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1036; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1037; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1038; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1039; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1040; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1041; // @[BTB.scala 196:29:@2080.8]
  wire  _GEN_1044; // @[BTB.scala 196:29:@2080.8]
  wire  _GEN_1049; // @[BTB.scala 196:29:@2080.8]
  wire  _GEN_1054; // @[BTB.scala 196:29:@2080.8]
  wire [1:0] _GEN_1057; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1058; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1059; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1060; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1061; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1062; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1063; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1064; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1065; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1066; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1067; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1068; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1069; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1070; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1071; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1072; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1073; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1074; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1075; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1076; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1077; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1078; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1079; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1080; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1081; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1082; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1083; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1084; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1085; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1086; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1087; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1088; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1089; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1090; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1091; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1092; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1093; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1094; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1095; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1096; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1097; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1098; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1099; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1100; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1101; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1102; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1103; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1104; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1105; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1106; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1107; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1108; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1109; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1110; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1111; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1112; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1113; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1114; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1115; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1116; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1117; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1118; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1119; // @[BTB.scala 195:49:@2078.6]
  wire [1:0] _GEN_1120; // @[BTB.scala 195:49:@2078.6]
  wire  _GEN_1123; // @[BTB.scala 195:49:@2078.6]
  wire  _GEN_1128; // @[BTB.scala 195:49:@2078.6]
  wire  _GEN_1133; // @[BTB.scala 195:49:@2078.6]
  wire  _GEN_1136; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1137; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1138; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1139; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1140; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1141; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1142; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1143; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1144; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1145; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1146; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1147; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1148; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1149; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1150; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1151; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1152; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1153; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1154; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1155; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1156; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1157; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1158; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1159; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1160; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1161; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1162; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1163; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1164; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1165; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1166; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1167; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1168; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1169; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1170; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1171; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1172; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1173; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1174; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1175; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1176; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1177; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1178; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1179; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1180; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1181; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1182; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1183; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1184; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1185; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1186; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1187; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1188; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1189; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1190; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1191; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1192; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1193; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1194; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1195; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1196; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1197; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1198; // @[BTB.scala 183:23:@2062.4]
  wire  _GEN_1199; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1200; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1201; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1202; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1203; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1204; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1205; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1206; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1207; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1208; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1209; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1210; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1211; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1212; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1213; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1214; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1215; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1216; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1217; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1218; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1219; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1220; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1221; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1222; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1223; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1224; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1225; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1226; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1227; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1228; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1229; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1230; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1231; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1232; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1233; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1234; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1235; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1236; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1237; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1238; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1239; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1240; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1241; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1242; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1243; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1244; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1245; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1246; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1247; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1248; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1249; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1250; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1251; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1252; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1253; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1254; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1255; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1256; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1257; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1258; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1259; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1260; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1261; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1262; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1263; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1264; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1265; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1266; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1267; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1268; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1269; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1270; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1271; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1272; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1273; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1274; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1275; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1276; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1277; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1278; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1279; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1280; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1281; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1282; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1283; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1284; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1285; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1286; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1287; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1288; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1289; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1290; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1291; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1292; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1293; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1294; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1295; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1296; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1297; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1298; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1299; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1300; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1301; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1302; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1303; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1304; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1305; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1306; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1307; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1308; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1309; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1310; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1311; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1312; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1313; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1314; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1315; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1316; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1317; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1318; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1319; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1320; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1321; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1322; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1323; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1324; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1325; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1326; // @[BTB.scala 183:23:@2062.4]
  wire [31:0] _GEN_1327; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1328; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1329; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1330; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1331; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1332; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1333; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1334; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1335; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1336; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1337; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1338; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1339; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1340; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1341; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1342; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1343; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1344; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1345; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1346; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1347; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1348; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1349; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1350; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1351; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1352; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1353; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1354; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1355; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1356; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1357; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1358; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1359; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1360; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1361; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1362; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1363; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1364; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1365; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1366; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1367; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1368; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1369; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1370; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1371; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1372; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1373; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1374; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1375; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1376; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1377; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1378; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1379; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1380; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1381; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1382; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1383; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1384; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1385; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1386; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1387; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1388; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1389; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1390; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1391; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1392; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1393; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1394; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1395; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1396; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1397; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1398; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1399; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1400; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1401; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1402; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1403; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1404; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1405; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1406; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1407; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1408; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1409; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1410; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1411; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1412; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1413; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1414; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1415; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1416; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1417; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1418; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1419; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1420; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1421; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1422; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1423; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1424; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1425; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1426; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1427; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1428; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1429; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1430; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1431; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1432; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1433; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1434; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1435; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1436; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1437; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1438; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1439; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1440; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1441; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1442; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1443; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1444; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1445; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1446; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1447; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1448; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1449; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1450; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1451; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1452; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1453; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1454; // @[BTB.scala 183:23:@2062.4]
  wire [1:0] _GEN_1455; // @[BTB.scala 183:23:@2062.4]
  wire  _T_2181; // @[BTB.scala 212:21:@2128.4]
  wire  _T_2183; // @[BTB.scala 213:26:@2130.6]
  wire  _T_2184; // @[BTB.scala 213:23:@2131.6]
  wire  _GEN_1477; // @[BTB.scala 213:39:@2132.6]
  wire [31:0] _T_2191; // @[OneHot.scala 26:18:@2143.6]
  wire [31:0] _T_2192; // @[OneHot.scala 27:18:@2144.6]
  wire  _T_2194; // @[OneHot.scala 28:14:@2145.6]
  wire [31:0] _T_2195; // @[OneHot.scala 28:28:@2146.6]
  wire [15:0] _T_2196; // @[OneHot.scala 26:18:@2147.6]
  wire [15:0] _T_2197; // @[OneHot.scala 27:18:@2148.6]
  wire  _T_2199; // @[OneHot.scala 28:14:@2149.6]
  wire [15:0] _T_2200; // @[OneHot.scala 28:28:@2150.6]
  wire [7:0] _T_2201; // @[OneHot.scala 26:18:@2151.6]
  wire [7:0] _T_2202; // @[OneHot.scala 27:18:@2152.6]
  wire  _T_2204; // @[OneHot.scala 28:14:@2153.6]
  wire [7:0] _T_2205; // @[OneHot.scala 28:28:@2154.6]
  wire [3:0] _T_2206; // @[OneHot.scala 26:18:@2155.6]
  wire [3:0] _T_2207; // @[OneHot.scala 27:18:@2156.6]
  wire  _T_2209; // @[OneHot.scala 28:14:@2157.6]
  wire [3:0] _T_2210; // @[OneHot.scala 28:28:@2158.6]
  wire [1:0] _T_2211; // @[OneHot.scala 26:18:@2159.6]
  wire [1:0] _T_2212; // @[OneHot.scala 27:18:@2160.6]
  wire  _T_2214; // @[OneHot.scala 28:14:@2161.6]
  wire [1:0] _T_2215; // @[OneHot.scala 28:28:@2162.6]
  wire  _T_2216; // @[CircuitMath.scala 30:8:@2163.6]
  wire [5:0] _T_2221; // @[Cat.scala 30:58:@2168.6]
  wire  _T_2224; // @[BTB.scala 221:11:@2170.6]
  wire  _T_2225; // @[BTB.scala 231:47:@2174.6]
  wire  _T_2229; // @[BTB.scala 231:47:@2180.6]
  wire  _T_2233; // @[BTB.scala 231:47:@2186.6]
  wire  _T_2237; // @[BTB.scala 231:47:@2192.6]
  wire  _T_2241; // @[BTB.scala 231:47:@2198.6]
  wire  _T_2245; // @[BTB.scala 231:47:@2204.6]
  wire  _T_2249; // @[BTB.scala 231:47:@2210.6]
  wire  _T_2253; // @[BTB.scala 231:47:@2216.6]
  wire  _T_2257; // @[BTB.scala 231:47:@2222.6]
  wire  _T_2261; // @[BTB.scala 232:26:@2228.6]
  RAS RAS ( // @[BTB.scala 69:19:@54.4]
    .clock(RAS_clock),
    .reset(RAS_reset),
    .io_push_valid(RAS_io_push_valid),
    .io_push_bits(RAS_io_push_bits),
    .io_pop(RAS_io_pop),
    .io_peek(RAS_io_peek)
  );
  assign bht__T_1188_addr = gb_history ^ _T_1186;
  assign bht__T_1188_data = bht[bht__T_1188_addr]; // @[BTB.scala 67:16:@52.4]
  assign bht__T_1774_addr = fb_reg_gshare;
  assign bht__T_1774_data = bht[bht__T_1774_addr]; // @[BTB.scala 67:16:@52.4]
  assign bht__T_2148_data = {_T_2150,_T_2155};
  assign bht__T_2148_addr = fb_reg_gshare;
  assign bht__T_2148_mask = 1'h1;
  assign bht__T_2148_en = fb_reg_valid ? _GEN_1123 : 1'h0;
  assign bht__T_2166_data = {_T_2169,_T_2174};
  assign bht__T_2166_addr = fb_reg_gshare;
  assign bht__T_2166_mask = 1'h1;
  assign bht__T_2166_en = fb_reg_valid ? _GEN_1128 : 1'h0;
  assign bht__T_2177_data = 2'h2;
  assign bht__T_2177_addr = fb_reg_gshare;
  assign bht__T_2177_mask = 1'h1;
  assign bht__T_2177_en = fb_reg_valid ? _GEN_1133 : 1'h0;
  assign arb__T_1187_addr = gb_history ^ _T_1186;
  assign arb__T_1187_data = arb[arb__T_1187_addr]; // @[BTB.scala 68:16:@53.4]
  assign arb_gshare_sel_addr = fb_reg_gshare;
  assign arb_gshare_sel_data = arb[arb_gshare_sel_addr]; // @[BTB.scala 68:16:@53.4]
  assign arb__T_2185_data = 1'h1;
  assign arb__T_2185_addr = fb_reg_gshare;
  assign arb__T_2185_mask = 1'h1;
  assign arb__T_2185_en = _T_2181 ? _T_2184 : 1'h0;
  assign arb__T_2187_data = 1'h0;
  assign arb__T_2187_addr = fb_reg_gshare;
  assign arb__T_2187_mask = 1'h1;
  assign arb__T_2187_en = _T_2181 ? _GEN_1477 : 1'h0;
  assign _T_148 = io_if_pc + 32'h4; // @[BTB.scala 102:32:@383.4]
  assign predict_cont_tgt = io_if_pc + 32'h4; // @[BTB.scala 102:32:@384.4]
  assign _T_150 = btb_pc_0 == io_if_pc; // @[BTB.scala 103:42:@386.4]
  assign _T_151 = btb_pc_1 == io_if_pc; // @[BTB.scala 103:42:@387.4]
  assign _T_152 = btb_pc_2 == io_if_pc; // @[BTB.scala 103:42:@388.4]
  assign _T_153 = btb_pc_3 == io_if_pc; // @[BTB.scala 103:42:@389.4]
  assign _T_154 = btb_pc_4 == io_if_pc; // @[BTB.scala 103:42:@390.4]
  assign _T_155 = btb_pc_5 == io_if_pc; // @[BTB.scala 103:42:@391.4]
  assign _T_156 = btb_pc_6 == io_if_pc; // @[BTB.scala 103:42:@392.4]
  assign _T_157 = btb_pc_7 == io_if_pc; // @[BTB.scala 103:42:@393.4]
  assign _T_158 = btb_pc_8 == io_if_pc; // @[BTB.scala 103:42:@394.4]
  assign _T_159 = btb_pc_9 == io_if_pc; // @[BTB.scala 103:42:@395.4]
  assign _T_160 = btb_pc_10 == io_if_pc; // @[BTB.scala 103:42:@396.4]
  assign _T_161 = btb_pc_11 == io_if_pc; // @[BTB.scala 103:42:@397.4]
  assign _T_162 = btb_pc_12 == io_if_pc; // @[BTB.scala 103:42:@398.4]
  assign _T_163 = btb_pc_13 == io_if_pc; // @[BTB.scala 103:42:@399.4]
  assign _T_164 = btb_pc_14 == io_if_pc; // @[BTB.scala 103:42:@400.4]
  assign _T_165 = btb_pc_15 == io_if_pc; // @[BTB.scala 103:42:@401.4]
  assign _T_166 = btb_pc_16 == io_if_pc; // @[BTB.scala 103:42:@402.4]
  assign _T_167 = btb_pc_17 == io_if_pc; // @[BTB.scala 103:42:@403.4]
  assign _T_168 = btb_pc_18 == io_if_pc; // @[BTB.scala 103:42:@404.4]
  assign _T_169 = btb_pc_19 == io_if_pc; // @[BTB.scala 103:42:@405.4]
  assign _T_170 = btb_pc_20 == io_if_pc; // @[BTB.scala 103:42:@406.4]
  assign _T_171 = btb_pc_21 == io_if_pc; // @[BTB.scala 103:42:@407.4]
  assign _T_172 = btb_pc_22 == io_if_pc; // @[BTB.scala 103:42:@408.4]
  assign _T_173 = btb_pc_23 == io_if_pc; // @[BTB.scala 103:42:@409.4]
  assign _T_174 = btb_pc_24 == io_if_pc; // @[BTB.scala 103:42:@410.4]
  assign _T_175 = btb_pc_25 == io_if_pc; // @[BTB.scala 103:42:@411.4]
  assign _T_176 = btb_pc_26 == io_if_pc; // @[BTB.scala 103:42:@412.4]
  assign _T_177 = btb_pc_27 == io_if_pc; // @[BTB.scala 103:42:@413.4]
  assign _T_178 = btb_pc_28 == io_if_pc; // @[BTB.scala 103:42:@414.4]
  assign _T_179 = btb_pc_29 == io_if_pc; // @[BTB.scala 103:42:@415.4]
  assign _T_180 = btb_pc_30 == io_if_pc; // @[BTB.scala 103:42:@416.4]
  assign _T_181 = btb_pc_31 == io_if_pc; // @[BTB.scala 103:42:@417.4]
  assign _T_182 = btb_pc_32 == io_if_pc; // @[BTB.scala 103:42:@418.4]
  assign _T_183 = btb_pc_33 == io_if_pc; // @[BTB.scala 103:42:@419.4]
  assign _T_184 = btb_pc_34 == io_if_pc; // @[BTB.scala 103:42:@420.4]
  assign _T_185 = btb_pc_35 == io_if_pc; // @[BTB.scala 103:42:@421.4]
  assign _T_186 = btb_pc_36 == io_if_pc; // @[BTB.scala 103:42:@422.4]
  assign _T_187 = btb_pc_37 == io_if_pc; // @[BTB.scala 103:42:@423.4]
  assign _T_188 = btb_pc_38 == io_if_pc; // @[BTB.scala 103:42:@424.4]
  assign _T_189 = btb_pc_39 == io_if_pc; // @[BTB.scala 103:42:@425.4]
  assign _T_190 = btb_pc_40 == io_if_pc; // @[BTB.scala 103:42:@426.4]
  assign _T_191 = btb_pc_41 == io_if_pc; // @[BTB.scala 103:42:@427.4]
  assign _T_192 = btb_pc_42 == io_if_pc; // @[BTB.scala 103:42:@428.4]
  assign _T_193 = btb_pc_43 == io_if_pc; // @[BTB.scala 103:42:@429.4]
  assign _T_194 = btb_pc_44 == io_if_pc; // @[BTB.scala 103:42:@430.4]
  assign _T_195 = btb_pc_45 == io_if_pc; // @[BTB.scala 103:42:@431.4]
  assign _T_196 = btb_pc_46 == io_if_pc; // @[BTB.scala 103:42:@432.4]
  assign _T_197 = btb_pc_47 == io_if_pc; // @[BTB.scala 103:42:@433.4]
  assign _T_198 = btb_pc_48 == io_if_pc; // @[BTB.scala 103:42:@434.4]
  assign _T_199 = btb_pc_49 == io_if_pc; // @[BTB.scala 103:42:@435.4]
  assign _T_200 = btb_pc_50 == io_if_pc; // @[BTB.scala 103:42:@436.4]
  assign _T_201 = btb_pc_51 == io_if_pc; // @[BTB.scala 103:42:@437.4]
  assign _T_202 = btb_pc_52 == io_if_pc; // @[BTB.scala 103:42:@438.4]
  assign _T_203 = btb_pc_53 == io_if_pc; // @[BTB.scala 103:42:@439.4]
  assign _T_204 = btb_pc_54 == io_if_pc; // @[BTB.scala 103:42:@440.4]
  assign _T_205 = btb_pc_55 == io_if_pc; // @[BTB.scala 103:42:@441.4]
  assign _T_206 = btb_pc_56 == io_if_pc; // @[BTB.scala 103:42:@442.4]
  assign _T_207 = btb_pc_57 == io_if_pc; // @[BTB.scala 103:42:@443.4]
  assign _T_208 = btb_pc_58 == io_if_pc; // @[BTB.scala 103:42:@444.4]
  assign _T_209 = btb_pc_59 == io_if_pc; // @[BTB.scala 103:42:@445.4]
  assign _T_210 = btb_pc_60 == io_if_pc; // @[BTB.scala 103:42:@446.4]
  assign _T_211 = btb_pc_61 == io_if_pc; // @[BTB.scala 103:42:@447.4]
  assign _T_212 = btb_pc_62 == io_if_pc; // @[BTB.scala 103:42:@448.4]
  assign _T_213 = btb_pc_63 == io_if_pc; // @[BTB.scala 103:42:@449.4]
  assign _T_290 = {_T_157,_T_156,_T_155,_T_154,_T_153,_T_152,_T_151,_T_150}; // @[BTB.scala 103:57:@521.4]
  assign _T_298 = {_T_165,_T_164,_T_163,_T_162,_T_161,_T_160,_T_159,_T_158,_T_290}; // @[BTB.scala 103:57:@529.4]
  assign _T_305 = {_T_173,_T_172,_T_171,_T_170,_T_169,_T_168,_T_167,_T_166}; // @[BTB.scala 103:57:@536.4]
  assign _T_314 = {_T_181,_T_180,_T_179,_T_178,_T_177,_T_176,_T_175,_T_174,_T_305,_T_298}; // @[BTB.scala 103:57:@545.4]
  assign _T_321 = {_T_189,_T_188,_T_187,_T_186,_T_185,_T_184,_T_183,_T_182}; // @[BTB.scala 103:57:@552.4]
  assign _T_329 = {_T_197,_T_196,_T_195,_T_194,_T_193,_T_192,_T_191,_T_190,_T_321}; // @[BTB.scala 103:57:@560.4]
  assign _T_336 = {_T_205,_T_204,_T_203,_T_202,_T_201,_T_200,_T_199,_T_198}; // @[BTB.scala 103:57:@567.4]
  assign _T_345 = {_T_213,_T_212,_T_211,_T_210,_T_209,_T_208,_T_207,_T_206,_T_336,_T_329}; // @[BTB.scala 103:57:@576.4]
  assign _T_346 = {_T_345,_T_314}; // @[BTB.scala 103:57:@577.4]
  assign _T_353 = {btb_valid_7,btb_valid_6,btb_valid_5,btb_valid_4,btb_valid_3,btb_valid_2,btb_valid_1,btb_valid_0}; // @[BTB.scala 103:76:@584.4]
  assign _T_361 = {btb_valid_15,btb_valid_14,btb_valid_13,btb_valid_12,btb_valid_11,btb_valid_10,btb_valid_9,btb_valid_8,_T_353}; // @[BTB.scala 103:76:@592.4]
  assign _T_368 = {btb_valid_23,btb_valid_22,btb_valid_21,btb_valid_20,btb_valid_19,btb_valid_18,btb_valid_17,btb_valid_16}; // @[BTB.scala 103:76:@599.4]
  assign _T_377 = {btb_valid_31,btb_valid_30,btb_valid_29,btb_valid_28,btb_valid_27,btb_valid_26,btb_valid_25,btb_valid_24,_T_368,_T_361}; // @[BTB.scala 103:76:@608.4]
  assign _T_384 = {btb_valid_39,btb_valid_38,btb_valid_37,btb_valid_36,btb_valid_35,btb_valid_34,btb_valid_33,btb_valid_32}; // @[BTB.scala 103:76:@615.4]
  assign _T_392 = {btb_valid_47,btb_valid_46,btb_valid_45,btb_valid_44,btb_valid_43,btb_valid_42,btb_valid_41,btb_valid_40,_T_384}; // @[BTB.scala 103:76:@623.4]
  assign _T_399 = {btb_valid_55,btb_valid_54,btb_valid_53,btb_valid_52,btb_valid_51,btb_valid_50,btb_valid_49,btb_valid_48}; // @[BTB.scala 103:76:@630.4]
  assign _T_408 = {btb_valid_63,btb_valid_62,btb_valid_61,btb_valid_60,btb_valid_59,btb_valid_58,btb_valid_57,btb_valid_56,_T_399,_T_392}; // @[BTB.scala 103:76:@639.4]
  assign _T_409 = {_T_408,_T_377}; // @[BTB.scala 103:76:@640.4]
  assign predict_lookup = _T_346 & _T_409; // @[BTB.scala 103:64:@641.4]
  assign _T_411 = predict_lookup[0]; // @[Mux.scala 21:36:@643.4]
  assign _T_412 = predict_lookup[1]; // @[Mux.scala 21:36:@644.4]
  assign _T_413 = predict_lookup[2]; // @[Mux.scala 21:36:@645.4]
  assign _T_414 = predict_lookup[3]; // @[Mux.scala 21:36:@646.4]
  assign _T_415 = predict_lookup[4]; // @[Mux.scala 21:36:@647.4]
  assign _T_416 = predict_lookup[5]; // @[Mux.scala 21:36:@648.4]
  assign _T_417 = predict_lookup[6]; // @[Mux.scala 21:36:@649.4]
  assign _T_418 = predict_lookup[7]; // @[Mux.scala 21:36:@650.4]
  assign _T_419 = predict_lookup[8]; // @[Mux.scala 21:36:@651.4]
  assign _T_420 = predict_lookup[9]; // @[Mux.scala 21:36:@652.4]
  assign _T_421 = predict_lookup[10]; // @[Mux.scala 21:36:@653.4]
  assign _T_422 = predict_lookup[11]; // @[Mux.scala 21:36:@654.4]
  assign _T_423 = predict_lookup[12]; // @[Mux.scala 21:36:@655.4]
  assign _T_424 = predict_lookup[13]; // @[Mux.scala 21:36:@656.4]
  assign _T_425 = predict_lookup[14]; // @[Mux.scala 21:36:@657.4]
  assign _T_426 = predict_lookup[15]; // @[Mux.scala 21:36:@658.4]
  assign _T_427 = predict_lookup[16]; // @[Mux.scala 21:36:@659.4]
  assign _T_428 = predict_lookup[17]; // @[Mux.scala 21:36:@660.4]
  assign _T_429 = predict_lookup[18]; // @[Mux.scala 21:36:@661.4]
  assign _T_430 = predict_lookup[19]; // @[Mux.scala 21:36:@662.4]
  assign _T_431 = predict_lookup[20]; // @[Mux.scala 21:36:@663.4]
  assign _T_432 = predict_lookup[21]; // @[Mux.scala 21:36:@664.4]
  assign _T_433 = predict_lookup[22]; // @[Mux.scala 21:36:@665.4]
  assign _T_434 = predict_lookup[23]; // @[Mux.scala 21:36:@666.4]
  assign _T_435 = predict_lookup[24]; // @[Mux.scala 21:36:@667.4]
  assign _T_436 = predict_lookup[25]; // @[Mux.scala 21:36:@668.4]
  assign _T_437 = predict_lookup[26]; // @[Mux.scala 21:36:@669.4]
  assign _T_438 = predict_lookup[27]; // @[Mux.scala 21:36:@670.4]
  assign _T_439 = predict_lookup[28]; // @[Mux.scala 21:36:@671.4]
  assign _T_440 = predict_lookup[29]; // @[Mux.scala 21:36:@672.4]
  assign _T_441 = predict_lookup[30]; // @[Mux.scala 21:36:@673.4]
  assign _T_442 = predict_lookup[31]; // @[Mux.scala 21:36:@674.4]
  assign _T_443 = predict_lookup[32]; // @[Mux.scala 21:36:@675.4]
  assign _T_444 = predict_lookup[33]; // @[Mux.scala 21:36:@676.4]
  assign _T_445 = predict_lookup[34]; // @[Mux.scala 21:36:@677.4]
  assign _T_446 = predict_lookup[35]; // @[Mux.scala 21:36:@678.4]
  assign _T_447 = predict_lookup[36]; // @[Mux.scala 21:36:@679.4]
  assign _T_448 = predict_lookup[37]; // @[Mux.scala 21:36:@680.4]
  assign _T_449 = predict_lookup[38]; // @[Mux.scala 21:36:@681.4]
  assign _T_450 = predict_lookup[39]; // @[Mux.scala 21:36:@682.4]
  assign _T_451 = predict_lookup[40]; // @[Mux.scala 21:36:@683.4]
  assign _T_452 = predict_lookup[41]; // @[Mux.scala 21:36:@684.4]
  assign _T_453 = predict_lookup[42]; // @[Mux.scala 21:36:@685.4]
  assign _T_454 = predict_lookup[43]; // @[Mux.scala 21:36:@686.4]
  assign _T_455 = predict_lookup[44]; // @[Mux.scala 21:36:@687.4]
  assign _T_456 = predict_lookup[45]; // @[Mux.scala 21:36:@688.4]
  assign _T_457 = predict_lookup[46]; // @[Mux.scala 21:36:@689.4]
  assign _T_458 = predict_lookup[47]; // @[Mux.scala 21:36:@690.4]
  assign _T_459 = predict_lookup[48]; // @[Mux.scala 21:36:@691.4]
  assign _T_460 = predict_lookup[49]; // @[Mux.scala 21:36:@692.4]
  assign _T_461 = predict_lookup[50]; // @[Mux.scala 21:36:@693.4]
  assign _T_462 = predict_lookup[51]; // @[Mux.scala 21:36:@694.4]
  assign _T_463 = predict_lookup[52]; // @[Mux.scala 21:36:@695.4]
  assign _T_464 = predict_lookup[53]; // @[Mux.scala 21:36:@696.4]
  assign _T_465 = predict_lookup[54]; // @[Mux.scala 21:36:@697.4]
  assign _T_466 = predict_lookup[55]; // @[Mux.scala 21:36:@698.4]
  assign _T_467 = predict_lookup[56]; // @[Mux.scala 21:36:@699.4]
  assign _T_468 = predict_lookup[57]; // @[Mux.scala 21:36:@700.4]
  assign _T_469 = predict_lookup[58]; // @[Mux.scala 21:36:@701.4]
  assign _T_470 = predict_lookup[59]; // @[Mux.scala 21:36:@702.4]
  assign _T_471 = predict_lookup[60]; // @[Mux.scala 21:36:@703.4]
  assign _T_472 = predict_lookup[61]; // @[Mux.scala 21:36:@704.4]
  assign _T_473 = predict_lookup[62]; // @[Mux.scala 21:36:@705.4]
  assign _T_474 = predict_lookup[63]; // @[Mux.scala 21:36:@706.4]
  assign _T_477 = _T_411 ? btb_tgt_0 : 32'h0; // @[Mux.scala 19:72:@707.4]
  assign _T_479 = _T_412 ? btb_tgt_1 : 32'h0; // @[Mux.scala 19:72:@708.4]
  assign _T_481 = _T_413 ? btb_tgt_2 : 32'h0; // @[Mux.scala 19:72:@709.4]
  assign _T_483 = _T_414 ? btb_tgt_3 : 32'h0; // @[Mux.scala 19:72:@710.4]
  assign _T_485 = _T_415 ? btb_tgt_4 : 32'h0; // @[Mux.scala 19:72:@711.4]
  assign _T_487 = _T_416 ? btb_tgt_5 : 32'h0; // @[Mux.scala 19:72:@712.4]
  assign _T_489 = _T_417 ? btb_tgt_6 : 32'h0; // @[Mux.scala 19:72:@713.4]
  assign _T_491 = _T_418 ? btb_tgt_7 : 32'h0; // @[Mux.scala 19:72:@714.4]
  assign _T_493 = _T_419 ? btb_tgt_8 : 32'h0; // @[Mux.scala 19:72:@715.4]
  assign _T_495 = _T_420 ? btb_tgt_9 : 32'h0; // @[Mux.scala 19:72:@716.4]
  assign _T_497 = _T_421 ? btb_tgt_10 : 32'h0; // @[Mux.scala 19:72:@717.4]
  assign _T_499 = _T_422 ? btb_tgt_11 : 32'h0; // @[Mux.scala 19:72:@718.4]
  assign _T_501 = _T_423 ? btb_tgt_12 : 32'h0; // @[Mux.scala 19:72:@719.4]
  assign _T_503 = _T_424 ? btb_tgt_13 : 32'h0; // @[Mux.scala 19:72:@720.4]
  assign _T_505 = _T_425 ? btb_tgt_14 : 32'h0; // @[Mux.scala 19:72:@721.4]
  assign _T_507 = _T_426 ? btb_tgt_15 : 32'h0; // @[Mux.scala 19:72:@722.4]
  assign _T_509 = _T_427 ? btb_tgt_16 : 32'h0; // @[Mux.scala 19:72:@723.4]
  assign _T_511 = _T_428 ? btb_tgt_17 : 32'h0; // @[Mux.scala 19:72:@724.4]
  assign _T_513 = _T_429 ? btb_tgt_18 : 32'h0; // @[Mux.scala 19:72:@725.4]
  assign _T_515 = _T_430 ? btb_tgt_19 : 32'h0; // @[Mux.scala 19:72:@726.4]
  assign _T_517 = _T_431 ? btb_tgt_20 : 32'h0; // @[Mux.scala 19:72:@727.4]
  assign _T_519 = _T_432 ? btb_tgt_21 : 32'h0; // @[Mux.scala 19:72:@728.4]
  assign _T_521 = _T_433 ? btb_tgt_22 : 32'h0; // @[Mux.scala 19:72:@729.4]
  assign _T_523 = _T_434 ? btb_tgt_23 : 32'h0; // @[Mux.scala 19:72:@730.4]
  assign _T_525 = _T_435 ? btb_tgt_24 : 32'h0; // @[Mux.scala 19:72:@731.4]
  assign _T_527 = _T_436 ? btb_tgt_25 : 32'h0; // @[Mux.scala 19:72:@732.4]
  assign _T_529 = _T_437 ? btb_tgt_26 : 32'h0; // @[Mux.scala 19:72:@733.4]
  assign _T_531 = _T_438 ? btb_tgt_27 : 32'h0; // @[Mux.scala 19:72:@734.4]
  assign _T_533 = _T_439 ? btb_tgt_28 : 32'h0; // @[Mux.scala 19:72:@735.4]
  assign _T_535 = _T_440 ? btb_tgt_29 : 32'h0; // @[Mux.scala 19:72:@736.4]
  assign _T_537 = _T_441 ? btb_tgt_30 : 32'h0; // @[Mux.scala 19:72:@737.4]
  assign _T_539 = _T_442 ? btb_tgt_31 : 32'h0; // @[Mux.scala 19:72:@738.4]
  assign _T_541 = _T_443 ? btb_tgt_32 : 32'h0; // @[Mux.scala 19:72:@739.4]
  assign _T_543 = _T_444 ? btb_tgt_33 : 32'h0; // @[Mux.scala 19:72:@740.4]
  assign _T_545 = _T_445 ? btb_tgt_34 : 32'h0; // @[Mux.scala 19:72:@741.4]
  assign _T_547 = _T_446 ? btb_tgt_35 : 32'h0; // @[Mux.scala 19:72:@742.4]
  assign _T_549 = _T_447 ? btb_tgt_36 : 32'h0; // @[Mux.scala 19:72:@743.4]
  assign _T_551 = _T_448 ? btb_tgt_37 : 32'h0; // @[Mux.scala 19:72:@744.4]
  assign _T_553 = _T_449 ? btb_tgt_38 : 32'h0; // @[Mux.scala 19:72:@745.4]
  assign _T_555 = _T_450 ? btb_tgt_39 : 32'h0; // @[Mux.scala 19:72:@746.4]
  assign _T_557 = _T_451 ? btb_tgt_40 : 32'h0; // @[Mux.scala 19:72:@747.4]
  assign _T_559 = _T_452 ? btb_tgt_41 : 32'h0; // @[Mux.scala 19:72:@748.4]
  assign _T_561 = _T_453 ? btb_tgt_42 : 32'h0; // @[Mux.scala 19:72:@749.4]
  assign _T_563 = _T_454 ? btb_tgt_43 : 32'h0; // @[Mux.scala 19:72:@750.4]
  assign _T_565 = _T_455 ? btb_tgt_44 : 32'h0; // @[Mux.scala 19:72:@751.4]
  assign _T_567 = _T_456 ? btb_tgt_45 : 32'h0; // @[Mux.scala 19:72:@752.4]
  assign _T_569 = _T_457 ? btb_tgt_46 : 32'h0; // @[Mux.scala 19:72:@753.4]
  assign _T_571 = _T_458 ? btb_tgt_47 : 32'h0; // @[Mux.scala 19:72:@754.4]
  assign _T_573 = _T_459 ? btb_tgt_48 : 32'h0; // @[Mux.scala 19:72:@755.4]
  assign _T_575 = _T_460 ? btb_tgt_49 : 32'h0; // @[Mux.scala 19:72:@756.4]
  assign _T_577 = _T_461 ? btb_tgt_50 : 32'h0; // @[Mux.scala 19:72:@757.4]
  assign _T_579 = _T_462 ? btb_tgt_51 : 32'h0; // @[Mux.scala 19:72:@758.4]
  assign _T_581 = _T_463 ? btb_tgt_52 : 32'h0; // @[Mux.scala 19:72:@759.4]
  assign _T_583 = _T_464 ? btb_tgt_53 : 32'h0; // @[Mux.scala 19:72:@760.4]
  assign _T_585 = _T_465 ? btb_tgt_54 : 32'h0; // @[Mux.scala 19:72:@761.4]
  assign _T_587 = _T_466 ? btb_tgt_55 : 32'h0; // @[Mux.scala 19:72:@762.4]
  assign _T_589 = _T_467 ? btb_tgt_56 : 32'h0; // @[Mux.scala 19:72:@763.4]
  assign _T_591 = _T_468 ? btb_tgt_57 : 32'h0; // @[Mux.scala 19:72:@764.4]
  assign _T_593 = _T_469 ? btb_tgt_58 : 32'h0; // @[Mux.scala 19:72:@765.4]
  assign _T_595 = _T_470 ? btb_tgt_59 : 32'h0; // @[Mux.scala 19:72:@766.4]
  assign _T_597 = _T_471 ? btb_tgt_60 : 32'h0; // @[Mux.scala 19:72:@767.4]
  assign _T_599 = _T_472 ? btb_tgt_61 : 32'h0; // @[Mux.scala 19:72:@768.4]
  assign _T_601 = _T_473 ? btb_tgt_62 : 32'h0; // @[Mux.scala 19:72:@769.4]
  assign _T_603 = _T_474 ? btb_tgt_63 : 32'h0; // @[Mux.scala 19:72:@770.4]
  assign _T_604 = _T_477 | _T_479; // @[Mux.scala 19:72:@771.4]
  assign _T_605 = _T_604 | _T_481; // @[Mux.scala 19:72:@772.4]
  assign _T_606 = _T_605 | _T_483; // @[Mux.scala 19:72:@773.4]
  assign _T_607 = _T_606 | _T_485; // @[Mux.scala 19:72:@774.4]
  assign _T_608 = _T_607 | _T_487; // @[Mux.scala 19:72:@775.4]
  assign _T_609 = _T_608 | _T_489; // @[Mux.scala 19:72:@776.4]
  assign _T_610 = _T_609 | _T_491; // @[Mux.scala 19:72:@777.4]
  assign _T_611 = _T_610 | _T_493; // @[Mux.scala 19:72:@778.4]
  assign _T_612 = _T_611 | _T_495; // @[Mux.scala 19:72:@779.4]
  assign _T_613 = _T_612 | _T_497; // @[Mux.scala 19:72:@780.4]
  assign _T_614 = _T_613 | _T_499; // @[Mux.scala 19:72:@781.4]
  assign _T_615 = _T_614 | _T_501; // @[Mux.scala 19:72:@782.4]
  assign _T_616 = _T_615 | _T_503; // @[Mux.scala 19:72:@783.4]
  assign _T_617 = _T_616 | _T_505; // @[Mux.scala 19:72:@784.4]
  assign _T_618 = _T_617 | _T_507; // @[Mux.scala 19:72:@785.4]
  assign _T_619 = _T_618 | _T_509; // @[Mux.scala 19:72:@786.4]
  assign _T_620 = _T_619 | _T_511; // @[Mux.scala 19:72:@787.4]
  assign _T_621 = _T_620 | _T_513; // @[Mux.scala 19:72:@788.4]
  assign _T_622 = _T_621 | _T_515; // @[Mux.scala 19:72:@789.4]
  assign _T_623 = _T_622 | _T_517; // @[Mux.scala 19:72:@790.4]
  assign _T_624 = _T_623 | _T_519; // @[Mux.scala 19:72:@791.4]
  assign _T_625 = _T_624 | _T_521; // @[Mux.scala 19:72:@792.4]
  assign _T_626 = _T_625 | _T_523; // @[Mux.scala 19:72:@793.4]
  assign _T_627 = _T_626 | _T_525; // @[Mux.scala 19:72:@794.4]
  assign _T_628 = _T_627 | _T_527; // @[Mux.scala 19:72:@795.4]
  assign _T_629 = _T_628 | _T_529; // @[Mux.scala 19:72:@796.4]
  assign _T_630 = _T_629 | _T_531; // @[Mux.scala 19:72:@797.4]
  assign _T_631 = _T_630 | _T_533; // @[Mux.scala 19:72:@798.4]
  assign _T_632 = _T_631 | _T_535; // @[Mux.scala 19:72:@799.4]
  assign _T_633 = _T_632 | _T_537; // @[Mux.scala 19:72:@800.4]
  assign _T_634 = _T_633 | _T_539; // @[Mux.scala 19:72:@801.4]
  assign _T_635 = _T_634 | _T_541; // @[Mux.scala 19:72:@802.4]
  assign _T_636 = _T_635 | _T_543; // @[Mux.scala 19:72:@803.4]
  assign _T_637 = _T_636 | _T_545; // @[Mux.scala 19:72:@804.4]
  assign _T_638 = _T_637 | _T_547; // @[Mux.scala 19:72:@805.4]
  assign _T_639 = _T_638 | _T_549; // @[Mux.scala 19:72:@806.4]
  assign _T_640 = _T_639 | _T_551; // @[Mux.scala 19:72:@807.4]
  assign _T_641 = _T_640 | _T_553; // @[Mux.scala 19:72:@808.4]
  assign _T_642 = _T_641 | _T_555; // @[Mux.scala 19:72:@809.4]
  assign _T_643 = _T_642 | _T_557; // @[Mux.scala 19:72:@810.4]
  assign _T_644 = _T_643 | _T_559; // @[Mux.scala 19:72:@811.4]
  assign _T_645 = _T_644 | _T_561; // @[Mux.scala 19:72:@812.4]
  assign _T_646 = _T_645 | _T_563; // @[Mux.scala 19:72:@813.4]
  assign _T_647 = _T_646 | _T_565; // @[Mux.scala 19:72:@814.4]
  assign _T_648 = _T_647 | _T_567; // @[Mux.scala 19:72:@815.4]
  assign _T_649 = _T_648 | _T_569; // @[Mux.scala 19:72:@816.4]
  assign _T_650 = _T_649 | _T_571; // @[Mux.scala 19:72:@817.4]
  assign _T_651 = _T_650 | _T_573; // @[Mux.scala 19:72:@818.4]
  assign _T_652 = _T_651 | _T_575; // @[Mux.scala 19:72:@819.4]
  assign _T_653 = _T_652 | _T_577; // @[Mux.scala 19:72:@820.4]
  assign _T_654 = _T_653 | _T_579; // @[Mux.scala 19:72:@821.4]
  assign _T_655 = _T_654 | _T_581; // @[Mux.scala 19:72:@822.4]
  assign _T_656 = _T_655 | _T_583; // @[Mux.scala 19:72:@823.4]
  assign _T_657 = _T_656 | _T_585; // @[Mux.scala 19:72:@824.4]
  assign _T_658 = _T_657 | _T_587; // @[Mux.scala 19:72:@825.4]
  assign _T_659 = _T_658 | _T_589; // @[Mux.scala 19:72:@826.4]
  assign _T_660 = _T_659 | _T_591; // @[Mux.scala 19:72:@827.4]
  assign _T_661 = _T_660 | _T_593; // @[Mux.scala 19:72:@828.4]
  assign _T_662 = _T_661 | _T_595; // @[Mux.scala 19:72:@829.4]
  assign _T_663 = _T_662 | _T_597; // @[Mux.scala 19:72:@830.4]
  assign _T_664 = _T_663 | _T_599; // @[Mux.scala 19:72:@831.4]
  assign _T_665 = _T_664 | _T_601; // @[Mux.scala 19:72:@832.4]
  assign predict_jump_tgt = _T_665 | _T_603; // @[Mux.scala 19:72:@833.4]
  assign _T_735 = _T_411 ? btb_bj_type_0 : 2'h0; // @[Mux.scala 19:72:@901.4]
  assign _T_737 = _T_412 ? btb_bj_type_1 : 2'h0; // @[Mux.scala 19:72:@902.4]
  assign _T_739 = _T_413 ? btb_bj_type_2 : 2'h0; // @[Mux.scala 19:72:@903.4]
  assign _T_741 = _T_414 ? btb_bj_type_3 : 2'h0; // @[Mux.scala 19:72:@904.4]
  assign _T_743 = _T_415 ? btb_bj_type_4 : 2'h0; // @[Mux.scala 19:72:@905.4]
  assign _T_745 = _T_416 ? btb_bj_type_5 : 2'h0; // @[Mux.scala 19:72:@906.4]
  assign _T_747 = _T_417 ? btb_bj_type_6 : 2'h0; // @[Mux.scala 19:72:@907.4]
  assign _T_749 = _T_418 ? btb_bj_type_7 : 2'h0; // @[Mux.scala 19:72:@908.4]
  assign _T_751 = _T_419 ? btb_bj_type_8 : 2'h0; // @[Mux.scala 19:72:@909.4]
  assign _T_753 = _T_420 ? btb_bj_type_9 : 2'h0; // @[Mux.scala 19:72:@910.4]
  assign _T_755 = _T_421 ? btb_bj_type_10 : 2'h0; // @[Mux.scala 19:72:@911.4]
  assign _T_757 = _T_422 ? btb_bj_type_11 : 2'h0; // @[Mux.scala 19:72:@912.4]
  assign _T_759 = _T_423 ? btb_bj_type_12 : 2'h0; // @[Mux.scala 19:72:@913.4]
  assign _T_761 = _T_424 ? btb_bj_type_13 : 2'h0; // @[Mux.scala 19:72:@914.4]
  assign _T_763 = _T_425 ? btb_bj_type_14 : 2'h0; // @[Mux.scala 19:72:@915.4]
  assign _T_765 = _T_426 ? btb_bj_type_15 : 2'h0; // @[Mux.scala 19:72:@916.4]
  assign _T_767 = _T_427 ? btb_bj_type_16 : 2'h0; // @[Mux.scala 19:72:@917.4]
  assign _T_769 = _T_428 ? btb_bj_type_17 : 2'h0; // @[Mux.scala 19:72:@918.4]
  assign _T_771 = _T_429 ? btb_bj_type_18 : 2'h0; // @[Mux.scala 19:72:@919.4]
  assign _T_773 = _T_430 ? btb_bj_type_19 : 2'h0; // @[Mux.scala 19:72:@920.4]
  assign _T_775 = _T_431 ? btb_bj_type_20 : 2'h0; // @[Mux.scala 19:72:@921.4]
  assign _T_777 = _T_432 ? btb_bj_type_21 : 2'h0; // @[Mux.scala 19:72:@922.4]
  assign _T_779 = _T_433 ? btb_bj_type_22 : 2'h0; // @[Mux.scala 19:72:@923.4]
  assign _T_781 = _T_434 ? btb_bj_type_23 : 2'h0; // @[Mux.scala 19:72:@924.4]
  assign _T_783 = _T_435 ? btb_bj_type_24 : 2'h0; // @[Mux.scala 19:72:@925.4]
  assign _T_785 = _T_436 ? btb_bj_type_25 : 2'h0; // @[Mux.scala 19:72:@926.4]
  assign _T_787 = _T_437 ? btb_bj_type_26 : 2'h0; // @[Mux.scala 19:72:@927.4]
  assign _T_789 = _T_438 ? btb_bj_type_27 : 2'h0; // @[Mux.scala 19:72:@928.4]
  assign _T_791 = _T_439 ? btb_bj_type_28 : 2'h0; // @[Mux.scala 19:72:@929.4]
  assign _T_793 = _T_440 ? btb_bj_type_29 : 2'h0; // @[Mux.scala 19:72:@930.4]
  assign _T_795 = _T_441 ? btb_bj_type_30 : 2'h0; // @[Mux.scala 19:72:@931.4]
  assign _T_797 = _T_442 ? btb_bj_type_31 : 2'h0; // @[Mux.scala 19:72:@932.4]
  assign _T_799 = _T_443 ? btb_bj_type_32 : 2'h0; // @[Mux.scala 19:72:@933.4]
  assign _T_801 = _T_444 ? btb_bj_type_33 : 2'h0; // @[Mux.scala 19:72:@934.4]
  assign _T_803 = _T_445 ? btb_bj_type_34 : 2'h0; // @[Mux.scala 19:72:@935.4]
  assign _T_805 = _T_446 ? btb_bj_type_35 : 2'h0; // @[Mux.scala 19:72:@936.4]
  assign _T_807 = _T_447 ? btb_bj_type_36 : 2'h0; // @[Mux.scala 19:72:@937.4]
  assign _T_809 = _T_448 ? btb_bj_type_37 : 2'h0; // @[Mux.scala 19:72:@938.4]
  assign _T_811 = _T_449 ? btb_bj_type_38 : 2'h0; // @[Mux.scala 19:72:@939.4]
  assign _T_813 = _T_450 ? btb_bj_type_39 : 2'h0; // @[Mux.scala 19:72:@940.4]
  assign _T_815 = _T_451 ? btb_bj_type_40 : 2'h0; // @[Mux.scala 19:72:@941.4]
  assign _T_817 = _T_452 ? btb_bj_type_41 : 2'h0; // @[Mux.scala 19:72:@942.4]
  assign _T_819 = _T_453 ? btb_bj_type_42 : 2'h0; // @[Mux.scala 19:72:@943.4]
  assign _T_821 = _T_454 ? btb_bj_type_43 : 2'h0; // @[Mux.scala 19:72:@944.4]
  assign _T_823 = _T_455 ? btb_bj_type_44 : 2'h0; // @[Mux.scala 19:72:@945.4]
  assign _T_825 = _T_456 ? btb_bj_type_45 : 2'h0; // @[Mux.scala 19:72:@946.4]
  assign _T_827 = _T_457 ? btb_bj_type_46 : 2'h0; // @[Mux.scala 19:72:@947.4]
  assign _T_829 = _T_458 ? btb_bj_type_47 : 2'h0; // @[Mux.scala 19:72:@948.4]
  assign _T_831 = _T_459 ? btb_bj_type_48 : 2'h0; // @[Mux.scala 19:72:@949.4]
  assign _T_833 = _T_460 ? btb_bj_type_49 : 2'h0; // @[Mux.scala 19:72:@950.4]
  assign _T_835 = _T_461 ? btb_bj_type_50 : 2'h0; // @[Mux.scala 19:72:@951.4]
  assign _T_837 = _T_462 ? btb_bj_type_51 : 2'h0; // @[Mux.scala 19:72:@952.4]
  assign _T_839 = _T_463 ? btb_bj_type_52 : 2'h0; // @[Mux.scala 19:72:@953.4]
  assign _T_841 = _T_464 ? btb_bj_type_53 : 2'h0; // @[Mux.scala 19:72:@954.4]
  assign _T_843 = _T_465 ? btb_bj_type_54 : 2'h0; // @[Mux.scala 19:72:@955.4]
  assign _T_845 = _T_466 ? btb_bj_type_55 : 2'h0; // @[Mux.scala 19:72:@956.4]
  assign _T_847 = _T_467 ? btb_bj_type_56 : 2'h0; // @[Mux.scala 19:72:@957.4]
  assign _T_849 = _T_468 ? btb_bj_type_57 : 2'h0; // @[Mux.scala 19:72:@958.4]
  assign _T_851 = _T_469 ? btb_bj_type_58 : 2'h0; // @[Mux.scala 19:72:@959.4]
  assign _T_853 = _T_470 ? btb_bj_type_59 : 2'h0; // @[Mux.scala 19:72:@960.4]
  assign _T_855 = _T_471 ? btb_bj_type_60 : 2'h0; // @[Mux.scala 19:72:@961.4]
  assign _T_857 = _T_472 ? btb_bj_type_61 : 2'h0; // @[Mux.scala 19:72:@962.4]
  assign _T_859 = _T_473 ? btb_bj_type_62 : 2'h0; // @[Mux.scala 19:72:@963.4]
  assign _T_861 = _T_474 ? btb_bj_type_63 : 2'h0; // @[Mux.scala 19:72:@964.4]
  assign _T_862 = _T_735 | _T_737; // @[Mux.scala 19:72:@965.4]
  assign _T_863 = _T_862 | _T_739; // @[Mux.scala 19:72:@966.4]
  assign _T_864 = _T_863 | _T_741; // @[Mux.scala 19:72:@967.4]
  assign _T_865 = _T_864 | _T_743; // @[Mux.scala 19:72:@968.4]
  assign _T_866 = _T_865 | _T_745; // @[Mux.scala 19:72:@969.4]
  assign _T_867 = _T_866 | _T_747; // @[Mux.scala 19:72:@970.4]
  assign _T_868 = _T_867 | _T_749; // @[Mux.scala 19:72:@971.4]
  assign _T_869 = _T_868 | _T_751; // @[Mux.scala 19:72:@972.4]
  assign _T_870 = _T_869 | _T_753; // @[Mux.scala 19:72:@973.4]
  assign _T_871 = _T_870 | _T_755; // @[Mux.scala 19:72:@974.4]
  assign _T_872 = _T_871 | _T_757; // @[Mux.scala 19:72:@975.4]
  assign _T_873 = _T_872 | _T_759; // @[Mux.scala 19:72:@976.4]
  assign _T_874 = _T_873 | _T_761; // @[Mux.scala 19:72:@977.4]
  assign _T_875 = _T_874 | _T_763; // @[Mux.scala 19:72:@978.4]
  assign _T_876 = _T_875 | _T_765; // @[Mux.scala 19:72:@979.4]
  assign _T_877 = _T_876 | _T_767; // @[Mux.scala 19:72:@980.4]
  assign _T_878 = _T_877 | _T_769; // @[Mux.scala 19:72:@981.4]
  assign _T_879 = _T_878 | _T_771; // @[Mux.scala 19:72:@982.4]
  assign _T_880 = _T_879 | _T_773; // @[Mux.scala 19:72:@983.4]
  assign _T_881 = _T_880 | _T_775; // @[Mux.scala 19:72:@984.4]
  assign _T_882 = _T_881 | _T_777; // @[Mux.scala 19:72:@985.4]
  assign _T_883 = _T_882 | _T_779; // @[Mux.scala 19:72:@986.4]
  assign _T_884 = _T_883 | _T_781; // @[Mux.scala 19:72:@987.4]
  assign _T_885 = _T_884 | _T_783; // @[Mux.scala 19:72:@988.4]
  assign _T_886 = _T_885 | _T_785; // @[Mux.scala 19:72:@989.4]
  assign _T_887 = _T_886 | _T_787; // @[Mux.scala 19:72:@990.4]
  assign _T_888 = _T_887 | _T_789; // @[Mux.scala 19:72:@991.4]
  assign _T_889 = _T_888 | _T_791; // @[Mux.scala 19:72:@992.4]
  assign _T_890 = _T_889 | _T_793; // @[Mux.scala 19:72:@993.4]
  assign _T_891 = _T_890 | _T_795; // @[Mux.scala 19:72:@994.4]
  assign _T_892 = _T_891 | _T_797; // @[Mux.scala 19:72:@995.4]
  assign _T_893 = _T_892 | _T_799; // @[Mux.scala 19:72:@996.4]
  assign _T_894 = _T_893 | _T_801; // @[Mux.scala 19:72:@997.4]
  assign _T_895 = _T_894 | _T_803; // @[Mux.scala 19:72:@998.4]
  assign _T_896 = _T_895 | _T_805; // @[Mux.scala 19:72:@999.4]
  assign _T_897 = _T_896 | _T_807; // @[Mux.scala 19:72:@1000.4]
  assign _T_898 = _T_897 | _T_809; // @[Mux.scala 19:72:@1001.4]
  assign _T_899 = _T_898 | _T_811; // @[Mux.scala 19:72:@1002.4]
  assign _T_900 = _T_899 | _T_813; // @[Mux.scala 19:72:@1003.4]
  assign _T_901 = _T_900 | _T_815; // @[Mux.scala 19:72:@1004.4]
  assign _T_902 = _T_901 | _T_817; // @[Mux.scala 19:72:@1005.4]
  assign _T_903 = _T_902 | _T_819; // @[Mux.scala 19:72:@1006.4]
  assign _T_904 = _T_903 | _T_821; // @[Mux.scala 19:72:@1007.4]
  assign _T_905 = _T_904 | _T_823; // @[Mux.scala 19:72:@1008.4]
  assign _T_906 = _T_905 | _T_825; // @[Mux.scala 19:72:@1009.4]
  assign _T_907 = _T_906 | _T_827; // @[Mux.scala 19:72:@1010.4]
  assign _T_908 = _T_907 | _T_829; // @[Mux.scala 19:72:@1011.4]
  assign _T_909 = _T_908 | _T_831; // @[Mux.scala 19:72:@1012.4]
  assign _T_910 = _T_909 | _T_833; // @[Mux.scala 19:72:@1013.4]
  assign _T_911 = _T_910 | _T_835; // @[Mux.scala 19:72:@1014.4]
  assign _T_912 = _T_911 | _T_837; // @[Mux.scala 19:72:@1015.4]
  assign _T_913 = _T_912 | _T_839; // @[Mux.scala 19:72:@1016.4]
  assign _T_914 = _T_913 | _T_841; // @[Mux.scala 19:72:@1017.4]
  assign _T_915 = _T_914 | _T_843; // @[Mux.scala 19:72:@1018.4]
  assign _T_916 = _T_915 | _T_845; // @[Mux.scala 19:72:@1019.4]
  assign _T_917 = _T_916 | _T_847; // @[Mux.scala 19:72:@1020.4]
  assign _T_918 = _T_917 | _T_849; // @[Mux.scala 19:72:@1021.4]
  assign _T_919 = _T_918 | _T_851; // @[Mux.scala 19:72:@1022.4]
  assign _T_920 = _T_919 | _T_853; // @[Mux.scala 19:72:@1023.4]
  assign _T_921 = _T_920 | _T_855; // @[Mux.scala 19:72:@1024.4]
  assign _T_922 = _T_921 | _T_857; // @[Mux.scala 19:72:@1025.4]
  assign _T_923 = _T_922 | _T_859; // @[Mux.scala 19:72:@1026.4]
  assign predict_bj_type = _T_923 | _T_861; // @[Mux.scala 19:72:@1027.4]
  assign _T_993 = _T_411 ? btb_h_count_0 : 2'h0; // @[Mux.scala 19:72:@1095.4]
  assign _T_995 = _T_412 ? btb_h_count_1 : 2'h0; // @[Mux.scala 19:72:@1096.4]
  assign _T_997 = _T_413 ? btb_h_count_2 : 2'h0; // @[Mux.scala 19:72:@1097.4]
  assign _T_999 = _T_414 ? btb_h_count_3 : 2'h0; // @[Mux.scala 19:72:@1098.4]
  assign _T_1001 = _T_415 ? btb_h_count_4 : 2'h0; // @[Mux.scala 19:72:@1099.4]
  assign _T_1003 = _T_416 ? btb_h_count_5 : 2'h0; // @[Mux.scala 19:72:@1100.4]
  assign _T_1005 = _T_417 ? btb_h_count_6 : 2'h0; // @[Mux.scala 19:72:@1101.4]
  assign _T_1007 = _T_418 ? btb_h_count_7 : 2'h0; // @[Mux.scala 19:72:@1102.4]
  assign _T_1009 = _T_419 ? btb_h_count_8 : 2'h0; // @[Mux.scala 19:72:@1103.4]
  assign _T_1011 = _T_420 ? btb_h_count_9 : 2'h0; // @[Mux.scala 19:72:@1104.4]
  assign _T_1013 = _T_421 ? btb_h_count_10 : 2'h0; // @[Mux.scala 19:72:@1105.4]
  assign _T_1015 = _T_422 ? btb_h_count_11 : 2'h0; // @[Mux.scala 19:72:@1106.4]
  assign _T_1017 = _T_423 ? btb_h_count_12 : 2'h0; // @[Mux.scala 19:72:@1107.4]
  assign _T_1019 = _T_424 ? btb_h_count_13 : 2'h0; // @[Mux.scala 19:72:@1108.4]
  assign _T_1021 = _T_425 ? btb_h_count_14 : 2'h0; // @[Mux.scala 19:72:@1109.4]
  assign _T_1023 = _T_426 ? btb_h_count_15 : 2'h0; // @[Mux.scala 19:72:@1110.4]
  assign _T_1025 = _T_427 ? btb_h_count_16 : 2'h0; // @[Mux.scala 19:72:@1111.4]
  assign _T_1027 = _T_428 ? btb_h_count_17 : 2'h0; // @[Mux.scala 19:72:@1112.4]
  assign _T_1029 = _T_429 ? btb_h_count_18 : 2'h0; // @[Mux.scala 19:72:@1113.4]
  assign _T_1031 = _T_430 ? btb_h_count_19 : 2'h0; // @[Mux.scala 19:72:@1114.4]
  assign _T_1033 = _T_431 ? btb_h_count_20 : 2'h0; // @[Mux.scala 19:72:@1115.4]
  assign _T_1035 = _T_432 ? btb_h_count_21 : 2'h0; // @[Mux.scala 19:72:@1116.4]
  assign _T_1037 = _T_433 ? btb_h_count_22 : 2'h0; // @[Mux.scala 19:72:@1117.4]
  assign _T_1039 = _T_434 ? btb_h_count_23 : 2'h0; // @[Mux.scala 19:72:@1118.4]
  assign _T_1041 = _T_435 ? btb_h_count_24 : 2'h0; // @[Mux.scala 19:72:@1119.4]
  assign _T_1043 = _T_436 ? btb_h_count_25 : 2'h0; // @[Mux.scala 19:72:@1120.4]
  assign _T_1045 = _T_437 ? btb_h_count_26 : 2'h0; // @[Mux.scala 19:72:@1121.4]
  assign _T_1047 = _T_438 ? btb_h_count_27 : 2'h0; // @[Mux.scala 19:72:@1122.4]
  assign _T_1049 = _T_439 ? btb_h_count_28 : 2'h0; // @[Mux.scala 19:72:@1123.4]
  assign _T_1051 = _T_440 ? btb_h_count_29 : 2'h0; // @[Mux.scala 19:72:@1124.4]
  assign _T_1053 = _T_441 ? btb_h_count_30 : 2'h0; // @[Mux.scala 19:72:@1125.4]
  assign _T_1055 = _T_442 ? btb_h_count_31 : 2'h0; // @[Mux.scala 19:72:@1126.4]
  assign _T_1057 = _T_443 ? btb_h_count_32 : 2'h0; // @[Mux.scala 19:72:@1127.4]
  assign _T_1059 = _T_444 ? btb_h_count_33 : 2'h0; // @[Mux.scala 19:72:@1128.4]
  assign _T_1061 = _T_445 ? btb_h_count_34 : 2'h0; // @[Mux.scala 19:72:@1129.4]
  assign _T_1063 = _T_446 ? btb_h_count_35 : 2'h0; // @[Mux.scala 19:72:@1130.4]
  assign _T_1065 = _T_447 ? btb_h_count_36 : 2'h0; // @[Mux.scala 19:72:@1131.4]
  assign _T_1067 = _T_448 ? btb_h_count_37 : 2'h0; // @[Mux.scala 19:72:@1132.4]
  assign _T_1069 = _T_449 ? btb_h_count_38 : 2'h0; // @[Mux.scala 19:72:@1133.4]
  assign _T_1071 = _T_450 ? btb_h_count_39 : 2'h0; // @[Mux.scala 19:72:@1134.4]
  assign _T_1073 = _T_451 ? btb_h_count_40 : 2'h0; // @[Mux.scala 19:72:@1135.4]
  assign _T_1075 = _T_452 ? btb_h_count_41 : 2'h0; // @[Mux.scala 19:72:@1136.4]
  assign _T_1077 = _T_453 ? btb_h_count_42 : 2'h0; // @[Mux.scala 19:72:@1137.4]
  assign _T_1079 = _T_454 ? btb_h_count_43 : 2'h0; // @[Mux.scala 19:72:@1138.4]
  assign _T_1081 = _T_455 ? btb_h_count_44 : 2'h0; // @[Mux.scala 19:72:@1139.4]
  assign _T_1083 = _T_456 ? btb_h_count_45 : 2'h0; // @[Mux.scala 19:72:@1140.4]
  assign _T_1085 = _T_457 ? btb_h_count_46 : 2'h0; // @[Mux.scala 19:72:@1141.4]
  assign _T_1087 = _T_458 ? btb_h_count_47 : 2'h0; // @[Mux.scala 19:72:@1142.4]
  assign _T_1089 = _T_459 ? btb_h_count_48 : 2'h0; // @[Mux.scala 19:72:@1143.4]
  assign _T_1091 = _T_460 ? btb_h_count_49 : 2'h0; // @[Mux.scala 19:72:@1144.4]
  assign _T_1093 = _T_461 ? btb_h_count_50 : 2'h0; // @[Mux.scala 19:72:@1145.4]
  assign _T_1095 = _T_462 ? btb_h_count_51 : 2'h0; // @[Mux.scala 19:72:@1146.4]
  assign _T_1097 = _T_463 ? btb_h_count_52 : 2'h0; // @[Mux.scala 19:72:@1147.4]
  assign _T_1099 = _T_464 ? btb_h_count_53 : 2'h0; // @[Mux.scala 19:72:@1148.4]
  assign _T_1101 = _T_465 ? btb_h_count_54 : 2'h0; // @[Mux.scala 19:72:@1149.4]
  assign _T_1103 = _T_466 ? btb_h_count_55 : 2'h0; // @[Mux.scala 19:72:@1150.4]
  assign _T_1105 = _T_467 ? btb_h_count_56 : 2'h0; // @[Mux.scala 19:72:@1151.4]
  assign _T_1107 = _T_468 ? btb_h_count_57 : 2'h0; // @[Mux.scala 19:72:@1152.4]
  assign _T_1109 = _T_469 ? btb_h_count_58 : 2'h0; // @[Mux.scala 19:72:@1153.4]
  assign _T_1111 = _T_470 ? btb_h_count_59 : 2'h0; // @[Mux.scala 19:72:@1154.4]
  assign _T_1113 = _T_471 ? btb_h_count_60 : 2'h0; // @[Mux.scala 19:72:@1155.4]
  assign _T_1115 = _T_472 ? btb_h_count_61 : 2'h0; // @[Mux.scala 19:72:@1156.4]
  assign _T_1117 = _T_473 ? btb_h_count_62 : 2'h0; // @[Mux.scala 19:72:@1157.4]
  assign _T_1119 = _T_474 ? btb_h_count_63 : 2'h0; // @[Mux.scala 19:72:@1158.4]
  assign _T_1120 = _T_993 | _T_995; // @[Mux.scala 19:72:@1159.4]
  assign _T_1121 = _T_1120 | _T_997; // @[Mux.scala 19:72:@1160.4]
  assign _T_1122 = _T_1121 | _T_999; // @[Mux.scala 19:72:@1161.4]
  assign _T_1123 = _T_1122 | _T_1001; // @[Mux.scala 19:72:@1162.4]
  assign _T_1124 = _T_1123 | _T_1003; // @[Mux.scala 19:72:@1163.4]
  assign _T_1125 = _T_1124 | _T_1005; // @[Mux.scala 19:72:@1164.4]
  assign _T_1126 = _T_1125 | _T_1007; // @[Mux.scala 19:72:@1165.4]
  assign _T_1127 = _T_1126 | _T_1009; // @[Mux.scala 19:72:@1166.4]
  assign _T_1128 = _T_1127 | _T_1011; // @[Mux.scala 19:72:@1167.4]
  assign _T_1129 = _T_1128 | _T_1013; // @[Mux.scala 19:72:@1168.4]
  assign _T_1130 = _T_1129 | _T_1015; // @[Mux.scala 19:72:@1169.4]
  assign _T_1131 = _T_1130 | _T_1017; // @[Mux.scala 19:72:@1170.4]
  assign _T_1132 = _T_1131 | _T_1019; // @[Mux.scala 19:72:@1171.4]
  assign _T_1133 = _T_1132 | _T_1021; // @[Mux.scala 19:72:@1172.4]
  assign _T_1134 = _T_1133 | _T_1023; // @[Mux.scala 19:72:@1173.4]
  assign _T_1135 = _T_1134 | _T_1025; // @[Mux.scala 19:72:@1174.4]
  assign _T_1136 = _T_1135 | _T_1027; // @[Mux.scala 19:72:@1175.4]
  assign _T_1137 = _T_1136 | _T_1029; // @[Mux.scala 19:72:@1176.4]
  assign _T_1138 = _T_1137 | _T_1031; // @[Mux.scala 19:72:@1177.4]
  assign _T_1139 = _T_1138 | _T_1033; // @[Mux.scala 19:72:@1178.4]
  assign _T_1140 = _T_1139 | _T_1035; // @[Mux.scala 19:72:@1179.4]
  assign _T_1141 = _T_1140 | _T_1037; // @[Mux.scala 19:72:@1180.4]
  assign _T_1142 = _T_1141 | _T_1039; // @[Mux.scala 19:72:@1181.4]
  assign _T_1143 = _T_1142 | _T_1041; // @[Mux.scala 19:72:@1182.4]
  assign _T_1144 = _T_1143 | _T_1043; // @[Mux.scala 19:72:@1183.4]
  assign _T_1145 = _T_1144 | _T_1045; // @[Mux.scala 19:72:@1184.4]
  assign _T_1146 = _T_1145 | _T_1047; // @[Mux.scala 19:72:@1185.4]
  assign _T_1147 = _T_1146 | _T_1049; // @[Mux.scala 19:72:@1186.4]
  assign _T_1148 = _T_1147 | _T_1051; // @[Mux.scala 19:72:@1187.4]
  assign _T_1149 = _T_1148 | _T_1053; // @[Mux.scala 19:72:@1188.4]
  assign _T_1150 = _T_1149 | _T_1055; // @[Mux.scala 19:72:@1189.4]
  assign _T_1151 = _T_1150 | _T_1057; // @[Mux.scala 19:72:@1190.4]
  assign _T_1152 = _T_1151 | _T_1059; // @[Mux.scala 19:72:@1191.4]
  assign _T_1153 = _T_1152 | _T_1061; // @[Mux.scala 19:72:@1192.4]
  assign _T_1154 = _T_1153 | _T_1063; // @[Mux.scala 19:72:@1193.4]
  assign _T_1155 = _T_1154 | _T_1065; // @[Mux.scala 19:72:@1194.4]
  assign _T_1156 = _T_1155 | _T_1067; // @[Mux.scala 19:72:@1195.4]
  assign _T_1157 = _T_1156 | _T_1069; // @[Mux.scala 19:72:@1196.4]
  assign _T_1158 = _T_1157 | _T_1071; // @[Mux.scala 19:72:@1197.4]
  assign _T_1159 = _T_1158 | _T_1073; // @[Mux.scala 19:72:@1198.4]
  assign _T_1160 = _T_1159 | _T_1075; // @[Mux.scala 19:72:@1199.4]
  assign _T_1161 = _T_1160 | _T_1077; // @[Mux.scala 19:72:@1200.4]
  assign _T_1162 = _T_1161 | _T_1079; // @[Mux.scala 19:72:@1201.4]
  assign _T_1163 = _T_1162 | _T_1081; // @[Mux.scala 19:72:@1202.4]
  assign _T_1164 = _T_1163 | _T_1083; // @[Mux.scala 19:72:@1203.4]
  assign _T_1165 = _T_1164 | _T_1085; // @[Mux.scala 19:72:@1204.4]
  assign _T_1166 = _T_1165 | _T_1087; // @[Mux.scala 19:72:@1205.4]
  assign _T_1167 = _T_1166 | _T_1089; // @[Mux.scala 19:72:@1206.4]
  assign _T_1168 = _T_1167 | _T_1091; // @[Mux.scala 19:72:@1207.4]
  assign _T_1169 = _T_1168 | _T_1093; // @[Mux.scala 19:72:@1208.4]
  assign _T_1170 = _T_1169 | _T_1095; // @[Mux.scala 19:72:@1209.4]
  assign _T_1171 = _T_1170 | _T_1097; // @[Mux.scala 19:72:@1210.4]
  assign _T_1172 = _T_1171 | _T_1099; // @[Mux.scala 19:72:@1211.4]
  assign _T_1173 = _T_1172 | _T_1101; // @[Mux.scala 19:72:@1212.4]
  assign _T_1174 = _T_1173 | _T_1103; // @[Mux.scala 19:72:@1213.4]
  assign _T_1175 = _T_1174 | _T_1105; // @[Mux.scala 19:72:@1214.4]
  assign _T_1176 = _T_1175 | _T_1107; // @[Mux.scala 19:72:@1215.4]
  assign _T_1177 = _T_1176 | _T_1109; // @[Mux.scala 19:72:@1216.4]
  assign _T_1178 = _T_1177 | _T_1111; // @[Mux.scala 19:72:@1217.4]
  assign _T_1179 = _T_1178 | _T_1113; // @[Mux.scala 19:72:@1218.4]
  assign _T_1180 = _T_1179 | _T_1115; // @[Mux.scala 19:72:@1219.4]
  assign _T_1181 = _T_1180 | _T_1117; // @[Mux.scala 19:72:@1220.4]
  assign predict_h_count = _T_1181 | _T_1119; // @[Mux.scala 19:72:@1221.4]
  assign _T_1186 = io_if_pc[11:2]; // @[BTB.scala 107:46:@1226.4]
  assign gshare_xor = gb_history ^ _T_1186; // @[BTB.scala 107:36:@1227.4]
  assign shift_wire = shift_reg & io_branch; // @[BTB.scala 111:30:@1233.4]
  assign _T_1191 = io_fb_type == 2'h2; // @[BTB.scala 113:22:@1235.6]
  assign _T_1192 = io_feedBack_history[8:0]; // @[BTB.scala 114:44:@1237.8]
  assign _T_1193 = {_T_1192,io_feedBack_redirect}; // @[Cat.scala 30:58:@1238.8]
  assign _GEN_0 = _T_1191 ? _T_1193 : io_feedBack_history; // @[BTB.scala 113:44:@1236.6]
  assign _T_1195 = predict_lookup != 64'h0; // @[BTB.scala 90:30:@1247.8]
  assign _T_1197 = predict_bj_type == 2'h2; // @[BTB.scala 97:41:@1248.8]
  assign _T_1198 = _T_1195 & _T_1197; // @[BTB.scala 97:30:@1249.8]
  assign _T_1200 = _T_1198 == 1'h0; // @[BTB.scala 119:18:@1250.8]
  assign _T_1201 = gb_history[8:0]; // @[BTB.scala 121:35:@1253.10]
  assign _T_1203 = {_T_1201,1'h0}; // @[Cat.scala 30:58:@1254.10]
  assign predict_gshare = bht__T_1188_data; // @[BTB.scala 88:21:@382.4 BTB.scala 109:20:@1231.4]
  assign _T_1210 = predict_gshare[1]; // @[BTB.scala 95:41:@1263.12]
  assign _T_1211 = predict_h_count[1]; // @[BTB.scala 95:53:@1264.12]
  assign predict_select = arb__T_1187_data; // @[BTB.scala 88:21:@382.4 BTB.scala 108:20:@1229.4]
  assign _T_1212 = predict_select ? _T_1210 : _T_1211; // @[BTB.scala 95:26:@1265.12]
  assign _T_1213 = {_T_1201,_T_1212}; // @[Cat.scala 30:58:@1266.12]
  assign _GEN_1 = _T_1198 ? _T_1213 : gb_history; // @[BTB.scala 122:32:@1261.10]
  assign _GEN_2 = shift_wire ? _T_1203 : _GEN_1; // @[BTB.scala 120:23:@1252.8]
  assign _GEN_3 = io_forward ? _T_1200 : shift_reg; // @[BTB.scala 118:26:@1246.6]
  assign _GEN_4 = io_forward ? _GEN_2 : gb_history; // @[BTB.scala 118:26:@1246.6]
  assign _GEN_5 = io_fb_miss ? _GEN_0 : _GEN_4; // @[BTB.scala 112:21:@1234.4]
  assign _T_1217 = predict_bj_type != 2'h2; // @[BTB.scala 98:44:@1271.4]
  assign _T_1221 = _T_1217 | _T_1212; // @[BTB.scala 98:65:@1275.4]
  assign _T_1222 = _T_1195 & _T_1221; // @[BTB.scala 98:32:@1276.4]
  assign _T_1227 = predict_bj_type == 2'h1; // @[BTB.scala 129:41:@1283.4]
  assign _T_1237 = _T_1222 ? predict_jump_tgt : predict_cont_tgt; // @[BTB.scala 130:8:@1291.4]
  assign _T_1247 = io_fb_pc[11:2]; // @[BTB.scala 167:57:@1313.4]
  assign _T_1248 = io_feedBack_history ^ _T_1247; // @[BTB.scala 167:47:@1314.4]
  assign _T_1249 = fb_reg_lfsr[0]; // @[BTB.scala 146:22:@1316.4]
  assign _T_1250 = fb_reg_lfsr[1]; // @[BTB.scala 146:32:@1317.4]
  assign _T_1251 = _T_1249 ^ _T_1250; // @[BTB.scala 146:26:@1318.4]
  assign _T_1252 = fb_reg_lfsr[5:1]; // @[BTB.scala 146:41:@1319.4]
  assign _T_1253 = {_T_1251,_T_1252}; // @[Cat.scala 30:58:@1320.4]
  assign _T_1255 = btb_pc_0 == fb_reg_pc; // @[BTB.scala 177:44:@1323.4]
  assign _T_1256 = btb_pc_1 == fb_reg_pc; // @[BTB.scala 177:44:@1324.4]
  assign _T_1257 = btb_pc_2 == fb_reg_pc; // @[BTB.scala 177:44:@1325.4]
  assign _T_1258 = btb_pc_3 == fb_reg_pc; // @[BTB.scala 177:44:@1326.4]
  assign _T_1259 = btb_pc_4 == fb_reg_pc; // @[BTB.scala 177:44:@1327.4]
  assign _T_1260 = btb_pc_5 == fb_reg_pc; // @[BTB.scala 177:44:@1328.4]
  assign _T_1261 = btb_pc_6 == fb_reg_pc; // @[BTB.scala 177:44:@1329.4]
  assign _T_1262 = btb_pc_7 == fb_reg_pc; // @[BTB.scala 177:44:@1330.4]
  assign _T_1263 = btb_pc_8 == fb_reg_pc; // @[BTB.scala 177:44:@1331.4]
  assign _T_1264 = btb_pc_9 == fb_reg_pc; // @[BTB.scala 177:44:@1332.4]
  assign _T_1265 = btb_pc_10 == fb_reg_pc; // @[BTB.scala 177:44:@1333.4]
  assign _T_1266 = btb_pc_11 == fb_reg_pc; // @[BTB.scala 177:44:@1334.4]
  assign _T_1267 = btb_pc_12 == fb_reg_pc; // @[BTB.scala 177:44:@1335.4]
  assign _T_1268 = btb_pc_13 == fb_reg_pc; // @[BTB.scala 177:44:@1336.4]
  assign _T_1269 = btb_pc_14 == fb_reg_pc; // @[BTB.scala 177:44:@1337.4]
  assign _T_1270 = btb_pc_15 == fb_reg_pc; // @[BTB.scala 177:44:@1338.4]
  assign _T_1271 = btb_pc_16 == fb_reg_pc; // @[BTB.scala 177:44:@1339.4]
  assign _T_1272 = btb_pc_17 == fb_reg_pc; // @[BTB.scala 177:44:@1340.4]
  assign _T_1273 = btb_pc_18 == fb_reg_pc; // @[BTB.scala 177:44:@1341.4]
  assign _T_1274 = btb_pc_19 == fb_reg_pc; // @[BTB.scala 177:44:@1342.4]
  assign _T_1275 = btb_pc_20 == fb_reg_pc; // @[BTB.scala 177:44:@1343.4]
  assign _T_1276 = btb_pc_21 == fb_reg_pc; // @[BTB.scala 177:44:@1344.4]
  assign _T_1277 = btb_pc_22 == fb_reg_pc; // @[BTB.scala 177:44:@1345.4]
  assign _T_1278 = btb_pc_23 == fb_reg_pc; // @[BTB.scala 177:44:@1346.4]
  assign _T_1279 = btb_pc_24 == fb_reg_pc; // @[BTB.scala 177:44:@1347.4]
  assign _T_1280 = btb_pc_25 == fb_reg_pc; // @[BTB.scala 177:44:@1348.4]
  assign _T_1281 = btb_pc_26 == fb_reg_pc; // @[BTB.scala 177:44:@1349.4]
  assign _T_1282 = btb_pc_27 == fb_reg_pc; // @[BTB.scala 177:44:@1350.4]
  assign _T_1283 = btb_pc_28 == fb_reg_pc; // @[BTB.scala 177:44:@1351.4]
  assign _T_1284 = btb_pc_29 == fb_reg_pc; // @[BTB.scala 177:44:@1352.4]
  assign _T_1285 = btb_pc_30 == fb_reg_pc; // @[BTB.scala 177:44:@1353.4]
  assign _T_1286 = btb_pc_31 == fb_reg_pc; // @[BTB.scala 177:44:@1354.4]
  assign _T_1287 = btb_pc_32 == fb_reg_pc; // @[BTB.scala 177:44:@1355.4]
  assign _T_1288 = btb_pc_33 == fb_reg_pc; // @[BTB.scala 177:44:@1356.4]
  assign _T_1289 = btb_pc_34 == fb_reg_pc; // @[BTB.scala 177:44:@1357.4]
  assign _T_1290 = btb_pc_35 == fb_reg_pc; // @[BTB.scala 177:44:@1358.4]
  assign _T_1291 = btb_pc_36 == fb_reg_pc; // @[BTB.scala 177:44:@1359.4]
  assign _T_1292 = btb_pc_37 == fb_reg_pc; // @[BTB.scala 177:44:@1360.4]
  assign _T_1293 = btb_pc_38 == fb_reg_pc; // @[BTB.scala 177:44:@1361.4]
  assign _T_1294 = btb_pc_39 == fb_reg_pc; // @[BTB.scala 177:44:@1362.4]
  assign _T_1295 = btb_pc_40 == fb_reg_pc; // @[BTB.scala 177:44:@1363.4]
  assign _T_1296 = btb_pc_41 == fb_reg_pc; // @[BTB.scala 177:44:@1364.4]
  assign _T_1297 = btb_pc_42 == fb_reg_pc; // @[BTB.scala 177:44:@1365.4]
  assign _T_1298 = btb_pc_43 == fb_reg_pc; // @[BTB.scala 177:44:@1366.4]
  assign _T_1299 = btb_pc_44 == fb_reg_pc; // @[BTB.scala 177:44:@1367.4]
  assign _T_1300 = btb_pc_45 == fb_reg_pc; // @[BTB.scala 177:44:@1368.4]
  assign _T_1301 = btb_pc_46 == fb_reg_pc; // @[BTB.scala 177:44:@1369.4]
  assign _T_1302 = btb_pc_47 == fb_reg_pc; // @[BTB.scala 177:44:@1370.4]
  assign _T_1303 = btb_pc_48 == fb_reg_pc; // @[BTB.scala 177:44:@1371.4]
  assign _T_1304 = btb_pc_49 == fb_reg_pc; // @[BTB.scala 177:44:@1372.4]
  assign _T_1305 = btb_pc_50 == fb_reg_pc; // @[BTB.scala 177:44:@1373.4]
  assign _T_1306 = btb_pc_51 == fb_reg_pc; // @[BTB.scala 177:44:@1374.4]
  assign _T_1307 = btb_pc_52 == fb_reg_pc; // @[BTB.scala 177:44:@1375.4]
  assign _T_1308 = btb_pc_53 == fb_reg_pc; // @[BTB.scala 177:44:@1376.4]
  assign _T_1309 = btb_pc_54 == fb_reg_pc; // @[BTB.scala 177:44:@1377.4]
  assign _T_1310 = btb_pc_55 == fb_reg_pc; // @[BTB.scala 177:44:@1378.4]
  assign _T_1311 = btb_pc_56 == fb_reg_pc; // @[BTB.scala 177:44:@1379.4]
  assign _T_1312 = btb_pc_57 == fb_reg_pc; // @[BTB.scala 177:44:@1380.4]
  assign _T_1313 = btb_pc_58 == fb_reg_pc; // @[BTB.scala 177:44:@1381.4]
  assign _T_1314 = btb_pc_59 == fb_reg_pc; // @[BTB.scala 177:44:@1382.4]
  assign _T_1315 = btb_pc_60 == fb_reg_pc; // @[BTB.scala 177:44:@1383.4]
  assign _T_1316 = btb_pc_61 == fb_reg_pc; // @[BTB.scala 177:44:@1384.4]
  assign _T_1317 = btb_pc_62 == fb_reg_pc; // @[BTB.scala 177:44:@1385.4]
  assign _T_1318 = btb_pc_63 == fb_reg_pc; // @[BTB.scala 177:44:@1386.4]
  assign _T_1395 = {_T_1262,_T_1261,_T_1260,_T_1259,_T_1258,_T_1257,_T_1256,_T_1255}; // @[BTB.scala 177:60:@1458.4]
  assign _T_1403 = {_T_1270,_T_1269,_T_1268,_T_1267,_T_1266,_T_1265,_T_1264,_T_1263,_T_1395}; // @[BTB.scala 177:60:@1466.4]
  assign _T_1410 = {_T_1278,_T_1277,_T_1276,_T_1275,_T_1274,_T_1273,_T_1272,_T_1271}; // @[BTB.scala 177:60:@1473.4]
  assign _T_1419 = {_T_1286,_T_1285,_T_1284,_T_1283,_T_1282,_T_1281,_T_1280,_T_1279,_T_1410,_T_1403}; // @[BTB.scala 177:60:@1482.4]
  assign _T_1426 = {_T_1294,_T_1293,_T_1292,_T_1291,_T_1290,_T_1289,_T_1288,_T_1287}; // @[BTB.scala 177:60:@1489.4]
  assign _T_1434 = {_T_1302,_T_1301,_T_1300,_T_1299,_T_1298,_T_1297,_T_1296,_T_1295,_T_1426}; // @[BTB.scala 177:60:@1497.4]
  assign _T_1441 = {_T_1310,_T_1309,_T_1308,_T_1307,_T_1306,_T_1305,_T_1304,_T_1303}; // @[BTB.scala 177:60:@1504.4]
  assign _T_1450 = {_T_1318,_T_1317,_T_1316,_T_1315,_T_1314,_T_1313,_T_1312,_T_1311,_T_1441,_T_1434}; // @[BTB.scala 177:60:@1513.4]
  assign _T_1451 = {_T_1450,_T_1419}; // @[BTB.scala 177:60:@1514.4]
  assign feedback_lookup = _T_1451 & _T_409; // @[BTB.scala 177:67:@1578.4]
  assign _T_1516 = feedback_lookup[0]; // @[Mux.scala 21:36:@1580.4]
  assign _T_1517 = feedback_lookup[1]; // @[Mux.scala 21:36:@1581.4]
  assign _T_1518 = feedback_lookup[2]; // @[Mux.scala 21:36:@1582.4]
  assign _T_1519 = feedback_lookup[3]; // @[Mux.scala 21:36:@1583.4]
  assign _T_1520 = feedback_lookup[4]; // @[Mux.scala 21:36:@1584.4]
  assign _T_1521 = feedback_lookup[5]; // @[Mux.scala 21:36:@1585.4]
  assign _T_1522 = feedback_lookup[6]; // @[Mux.scala 21:36:@1586.4]
  assign _T_1523 = feedback_lookup[7]; // @[Mux.scala 21:36:@1587.4]
  assign _T_1524 = feedback_lookup[8]; // @[Mux.scala 21:36:@1588.4]
  assign _T_1525 = feedback_lookup[9]; // @[Mux.scala 21:36:@1589.4]
  assign _T_1526 = feedback_lookup[10]; // @[Mux.scala 21:36:@1590.4]
  assign _T_1527 = feedback_lookup[11]; // @[Mux.scala 21:36:@1591.4]
  assign _T_1528 = feedback_lookup[12]; // @[Mux.scala 21:36:@1592.4]
  assign _T_1529 = feedback_lookup[13]; // @[Mux.scala 21:36:@1593.4]
  assign _T_1530 = feedback_lookup[14]; // @[Mux.scala 21:36:@1594.4]
  assign _T_1531 = feedback_lookup[15]; // @[Mux.scala 21:36:@1595.4]
  assign _T_1532 = feedback_lookup[16]; // @[Mux.scala 21:36:@1596.4]
  assign _T_1533 = feedback_lookup[17]; // @[Mux.scala 21:36:@1597.4]
  assign _T_1534 = feedback_lookup[18]; // @[Mux.scala 21:36:@1598.4]
  assign _T_1535 = feedback_lookup[19]; // @[Mux.scala 21:36:@1599.4]
  assign _T_1536 = feedback_lookup[20]; // @[Mux.scala 21:36:@1600.4]
  assign _T_1537 = feedback_lookup[21]; // @[Mux.scala 21:36:@1601.4]
  assign _T_1538 = feedback_lookup[22]; // @[Mux.scala 21:36:@1602.4]
  assign _T_1539 = feedback_lookup[23]; // @[Mux.scala 21:36:@1603.4]
  assign _T_1540 = feedback_lookup[24]; // @[Mux.scala 21:36:@1604.4]
  assign _T_1541 = feedback_lookup[25]; // @[Mux.scala 21:36:@1605.4]
  assign _T_1542 = feedback_lookup[26]; // @[Mux.scala 21:36:@1606.4]
  assign _T_1543 = feedback_lookup[27]; // @[Mux.scala 21:36:@1607.4]
  assign _T_1544 = feedback_lookup[28]; // @[Mux.scala 21:36:@1608.4]
  assign _T_1545 = feedback_lookup[29]; // @[Mux.scala 21:36:@1609.4]
  assign _T_1546 = feedback_lookup[30]; // @[Mux.scala 21:36:@1610.4]
  assign _T_1547 = feedback_lookup[31]; // @[Mux.scala 21:36:@1611.4]
  assign _T_1548 = feedback_lookup[32]; // @[Mux.scala 21:36:@1612.4]
  assign _T_1549 = feedback_lookup[33]; // @[Mux.scala 21:36:@1613.4]
  assign _T_1550 = feedback_lookup[34]; // @[Mux.scala 21:36:@1614.4]
  assign _T_1551 = feedback_lookup[35]; // @[Mux.scala 21:36:@1615.4]
  assign _T_1552 = feedback_lookup[36]; // @[Mux.scala 21:36:@1616.4]
  assign _T_1553 = feedback_lookup[37]; // @[Mux.scala 21:36:@1617.4]
  assign _T_1554 = feedback_lookup[38]; // @[Mux.scala 21:36:@1618.4]
  assign _T_1555 = feedback_lookup[39]; // @[Mux.scala 21:36:@1619.4]
  assign _T_1556 = feedback_lookup[40]; // @[Mux.scala 21:36:@1620.4]
  assign _T_1557 = feedback_lookup[41]; // @[Mux.scala 21:36:@1621.4]
  assign _T_1558 = feedback_lookup[42]; // @[Mux.scala 21:36:@1622.4]
  assign _T_1559 = feedback_lookup[43]; // @[Mux.scala 21:36:@1623.4]
  assign _T_1560 = feedback_lookup[44]; // @[Mux.scala 21:36:@1624.4]
  assign _T_1561 = feedback_lookup[45]; // @[Mux.scala 21:36:@1625.4]
  assign _T_1562 = feedback_lookup[46]; // @[Mux.scala 21:36:@1626.4]
  assign _T_1563 = feedback_lookup[47]; // @[Mux.scala 21:36:@1627.4]
  assign _T_1564 = feedback_lookup[48]; // @[Mux.scala 21:36:@1628.4]
  assign _T_1565 = feedback_lookup[49]; // @[Mux.scala 21:36:@1629.4]
  assign _T_1566 = feedback_lookup[50]; // @[Mux.scala 21:36:@1630.4]
  assign _T_1567 = feedback_lookup[51]; // @[Mux.scala 21:36:@1631.4]
  assign _T_1568 = feedback_lookup[52]; // @[Mux.scala 21:36:@1632.4]
  assign _T_1569 = feedback_lookup[53]; // @[Mux.scala 21:36:@1633.4]
  assign _T_1570 = feedback_lookup[54]; // @[Mux.scala 21:36:@1634.4]
  assign _T_1571 = feedback_lookup[55]; // @[Mux.scala 21:36:@1635.4]
  assign _T_1572 = feedback_lookup[56]; // @[Mux.scala 21:36:@1636.4]
  assign _T_1573 = feedback_lookup[57]; // @[Mux.scala 21:36:@1637.4]
  assign _T_1574 = feedback_lookup[58]; // @[Mux.scala 21:36:@1638.4]
  assign _T_1575 = feedback_lookup[59]; // @[Mux.scala 21:36:@1639.4]
  assign _T_1576 = feedback_lookup[60]; // @[Mux.scala 21:36:@1640.4]
  assign _T_1577 = feedback_lookup[61]; // @[Mux.scala 21:36:@1641.4]
  assign _T_1578 = feedback_lookup[62]; // @[Mux.scala 21:36:@1642.4]
  assign _T_1579 = feedback_lookup[63]; // @[Mux.scala 21:36:@1643.4]
  assign _T_1582 = _T_1516 ? btb_h_count_0 : 2'h0; // @[Mux.scala 19:72:@1644.4]
  assign _T_1584 = _T_1517 ? btb_h_count_1 : 2'h0; // @[Mux.scala 19:72:@1645.4]
  assign _T_1586 = _T_1518 ? btb_h_count_2 : 2'h0; // @[Mux.scala 19:72:@1646.4]
  assign _T_1588 = _T_1519 ? btb_h_count_3 : 2'h0; // @[Mux.scala 19:72:@1647.4]
  assign _T_1590 = _T_1520 ? btb_h_count_4 : 2'h0; // @[Mux.scala 19:72:@1648.4]
  assign _T_1592 = _T_1521 ? btb_h_count_5 : 2'h0; // @[Mux.scala 19:72:@1649.4]
  assign _T_1594 = _T_1522 ? btb_h_count_6 : 2'h0; // @[Mux.scala 19:72:@1650.4]
  assign _T_1596 = _T_1523 ? btb_h_count_7 : 2'h0; // @[Mux.scala 19:72:@1651.4]
  assign _T_1598 = _T_1524 ? btb_h_count_8 : 2'h0; // @[Mux.scala 19:72:@1652.4]
  assign _T_1600 = _T_1525 ? btb_h_count_9 : 2'h0; // @[Mux.scala 19:72:@1653.4]
  assign _T_1602 = _T_1526 ? btb_h_count_10 : 2'h0; // @[Mux.scala 19:72:@1654.4]
  assign _T_1604 = _T_1527 ? btb_h_count_11 : 2'h0; // @[Mux.scala 19:72:@1655.4]
  assign _T_1606 = _T_1528 ? btb_h_count_12 : 2'h0; // @[Mux.scala 19:72:@1656.4]
  assign _T_1608 = _T_1529 ? btb_h_count_13 : 2'h0; // @[Mux.scala 19:72:@1657.4]
  assign _T_1610 = _T_1530 ? btb_h_count_14 : 2'h0; // @[Mux.scala 19:72:@1658.4]
  assign _T_1612 = _T_1531 ? btb_h_count_15 : 2'h0; // @[Mux.scala 19:72:@1659.4]
  assign _T_1614 = _T_1532 ? btb_h_count_16 : 2'h0; // @[Mux.scala 19:72:@1660.4]
  assign _T_1616 = _T_1533 ? btb_h_count_17 : 2'h0; // @[Mux.scala 19:72:@1661.4]
  assign _T_1618 = _T_1534 ? btb_h_count_18 : 2'h0; // @[Mux.scala 19:72:@1662.4]
  assign _T_1620 = _T_1535 ? btb_h_count_19 : 2'h0; // @[Mux.scala 19:72:@1663.4]
  assign _T_1622 = _T_1536 ? btb_h_count_20 : 2'h0; // @[Mux.scala 19:72:@1664.4]
  assign _T_1624 = _T_1537 ? btb_h_count_21 : 2'h0; // @[Mux.scala 19:72:@1665.4]
  assign _T_1626 = _T_1538 ? btb_h_count_22 : 2'h0; // @[Mux.scala 19:72:@1666.4]
  assign _T_1628 = _T_1539 ? btb_h_count_23 : 2'h0; // @[Mux.scala 19:72:@1667.4]
  assign _T_1630 = _T_1540 ? btb_h_count_24 : 2'h0; // @[Mux.scala 19:72:@1668.4]
  assign _T_1632 = _T_1541 ? btb_h_count_25 : 2'h0; // @[Mux.scala 19:72:@1669.4]
  assign _T_1634 = _T_1542 ? btb_h_count_26 : 2'h0; // @[Mux.scala 19:72:@1670.4]
  assign _T_1636 = _T_1543 ? btb_h_count_27 : 2'h0; // @[Mux.scala 19:72:@1671.4]
  assign _T_1638 = _T_1544 ? btb_h_count_28 : 2'h0; // @[Mux.scala 19:72:@1672.4]
  assign _T_1640 = _T_1545 ? btb_h_count_29 : 2'h0; // @[Mux.scala 19:72:@1673.4]
  assign _T_1642 = _T_1546 ? btb_h_count_30 : 2'h0; // @[Mux.scala 19:72:@1674.4]
  assign _T_1644 = _T_1547 ? btb_h_count_31 : 2'h0; // @[Mux.scala 19:72:@1675.4]
  assign _T_1646 = _T_1548 ? btb_h_count_32 : 2'h0; // @[Mux.scala 19:72:@1676.4]
  assign _T_1648 = _T_1549 ? btb_h_count_33 : 2'h0; // @[Mux.scala 19:72:@1677.4]
  assign _T_1650 = _T_1550 ? btb_h_count_34 : 2'h0; // @[Mux.scala 19:72:@1678.4]
  assign _T_1652 = _T_1551 ? btb_h_count_35 : 2'h0; // @[Mux.scala 19:72:@1679.4]
  assign _T_1654 = _T_1552 ? btb_h_count_36 : 2'h0; // @[Mux.scala 19:72:@1680.4]
  assign _T_1656 = _T_1553 ? btb_h_count_37 : 2'h0; // @[Mux.scala 19:72:@1681.4]
  assign _T_1658 = _T_1554 ? btb_h_count_38 : 2'h0; // @[Mux.scala 19:72:@1682.4]
  assign _T_1660 = _T_1555 ? btb_h_count_39 : 2'h0; // @[Mux.scala 19:72:@1683.4]
  assign _T_1662 = _T_1556 ? btb_h_count_40 : 2'h0; // @[Mux.scala 19:72:@1684.4]
  assign _T_1664 = _T_1557 ? btb_h_count_41 : 2'h0; // @[Mux.scala 19:72:@1685.4]
  assign _T_1666 = _T_1558 ? btb_h_count_42 : 2'h0; // @[Mux.scala 19:72:@1686.4]
  assign _T_1668 = _T_1559 ? btb_h_count_43 : 2'h0; // @[Mux.scala 19:72:@1687.4]
  assign _T_1670 = _T_1560 ? btb_h_count_44 : 2'h0; // @[Mux.scala 19:72:@1688.4]
  assign _T_1672 = _T_1561 ? btb_h_count_45 : 2'h0; // @[Mux.scala 19:72:@1689.4]
  assign _T_1674 = _T_1562 ? btb_h_count_46 : 2'h0; // @[Mux.scala 19:72:@1690.4]
  assign _T_1676 = _T_1563 ? btb_h_count_47 : 2'h0; // @[Mux.scala 19:72:@1691.4]
  assign _T_1678 = _T_1564 ? btb_h_count_48 : 2'h0; // @[Mux.scala 19:72:@1692.4]
  assign _T_1680 = _T_1565 ? btb_h_count_49 : 2'h0; // @[Mux.scala 19:72:@1693.4]
  assign _T_1682 = _T_1566 ? btb_h_count_50 : 2'h0; // @[Mux.scala 19:72:@1694.4]
  assign _T_1684 = _T_1567 ? btb_h_count_51 : 2'h0; // @[Mux.scala 19:72:@1695.4]
  assign _T_1686 = _T_1568 ? btb_h_count_52 : 2'h0; // @[Mux.scala 19:72:@1696.4]
  assign _T_1688 = _T_1569 ? btb_h_count_53 : 2'h0; // @[Mux.scala 19:72:@1697.4]
  assign _T_1690 = _T_1570 ? btb_h_count_54 : 2'h0; // @[Mux.scala 19:72:@1698.4]
  assign _T_1692 = _T_1571 ? btb_h_count_55 : 2'h0; // @[Mux.scala 19:72:@1699.4]
  assign _T_1694 = _T_1572 ? btb_h_count_56 : 2'h0; // @[Mux.scala 19:72:@1700.4]
  assign _T_1696 = _T_1573 ? btb_h_count_57 : 2'h0; // @[Mux.scala 19:72:@1701.4]
  assign _T_1698 = _T_1574 ? btb_h_count_58 : 2'h0; // @[Mux.scala 19:72:@1702.4]
  assign _T_1700 = _T_1575 ? btb_h_count_59 : 2'h0; // @[Mux.scala 19:72:@1703.4]
  assign _T_1702 = _T_1576 ? btb_h_count_60 : 2'h0; // @[Mux.scala 19:72:@1704.4]
  assign _T_1704 = _T_1577 ? btb_h_count_61 : 2'h0; // @[Mux.scala 19:72:@1705.4]
  assign _T_1706 = _T_1578 ? btb_h_count_62 : 2'h0; // @[Mux.scala 19:72:@1706.4]
  assign _T_1708 = _T_1579 ? btb_h_count_63 : 2'h0; // @[Mux.scala 19:72:@1707.4]
  assign _T_1709 = _T_1582 | _T_1584; // @[Mux.scala 19:72:@1708.4]
  assign _T_1710 = _T_1709 | _T_1586; // @[Mux.scala 19:72:@1709.4]
  assign _T_1711 = _T_1710 | _T_1588; // @[Mux.scala 19:72:@1710.4]
  assign _T_1712 = _T_1711 | _T_1590; // @[Mux.scala 19:72:@1711.4]
  assign _T_1713 = _T_1712 | _T_1592; // @[Mux.scala 19:72:@1712.4]
  assign _T_1714 = _T_1713 | _T_1594; // @[Mux.scala 19:72:@1713.4]
  assign _T_1715 = _T_1714 | _T_1596; // @[Mux.scala 19:72:@1714.4]
  assign _T_1716 = _T_1715 | _T_1598; // @[Mux.scala 19:72:@1715.4]
  assign _T_1717 = _T_1716 | _T_1600; // @[Mux.scala 19:72:@1716.4]
  assign _T_1718 = _T_1717 | _T_1602; // @[Mux.scala 19:72:@1717.4]
  assign _T_1719 = _T_1718 | _T_1604; // @[Mux.scala 19:72:@1718.4]
  assign _T_1720 = _T_1719 | _T_1606; // @[Mux.scala 19:72:@1719.4]
  assign _T_1721 = _T_1720 | _T_1608; // @[Mux.scala 19:72:@1720.4]
  assign _T_1722 = _T_1721 | _T_1610; // @[Mux.scala 19:72:@1721.4]
  assign _T_1723 = _T_1722 | _T_1612; // @[Mux.scala 19:72:@1722.4]
  assign _T_1724 = _T_1723 | _T_1614; // @[Mux.scala 19:72:@1723.4]
  assign _T_1725 = _T_1724 | _T_1616; // @[Mux.scala 19:72:@1724.4]
  assign _T_1726 = _T_1725 | _T_1618; // @[Mux.scala 19:72:@1725.4]
  assign _T_1727 = _T_1726 | _T_1620; // @[Mux.scala 19:72:@1726.4]
  assign _T_1728 = _T_1727 | _T_1622; // @[Mux.scala 19:72:@1727.4]
  assign _T_1729 = _T_1728 | _T_1624; // @[Mux.scala 19:72:@1728.4]
  assign _T_1730 = _T_1729 | _T_1626; // @[Mux.scala 19:72:@1729.4]
  assign _T_1731 = _T_1730 | _T_1628; // @[Mux.scala 19:72:@1730.4]
  assign _T_1732 = _T_1731 | _T_1630; // @[Mux.scala 19:72:@1731.4]
  assign _T_1733 = _T_1732 | _T_1632; // @[Mux.scala 19:72:@1732.4]
  assign _T_1734 = _T_1733 | _T_1634; // @[Mux.scala 19:72:@1733.4]
  assign _T_1735 = _T_1734 | _T_1636; // @[Mux.scala 19:72:@1734.4]
  assign _T_1736 = _T_1735 | _T_1638; // @[Mux.scala 19:72:@1735.4]
  assign _T_1737 = _T_1736 | _T_1640; // @[Mux.scala 19:72:@1736.4]
  assign _T_1738 = _T_1737 | _T_1642; // @[Mux.scala 19:72:@1737.4]
  assign _T_1739 = _T_1738 | _T_1644; // @[Mux.scala 19:72:@1738.4]
  assign _T_1740 = _T_1739 | _T_1646; // @[Mux.scala 19:72:@1739.4]
  assign _T_1741 = _T_1740 | _T_1648; // @[Mux.scala 19:72:@1740.4]
  assign _T_1742 = _T_1741 | _T_1650; // @[Mux.scala 19:72:@1741.4]
  assign _T_1743 = _T_1742 | _T_1652; // @[Mux.scala 19:72:@1742.4]
  assign _T_1744 = _T_1743 | _T_1654; // @[Mux.scala 19:72:@1743.4]
  assign _T_1745 = _T_1744 | _T_1656; // @[Mux.scala 19:72:@1744.4]
  assign _T_1746 = _T_1745 | _T_1658; // @[Mux.scala 19:72:@1745.4]
  assign _T_1747 = _T_1746 | _T_1660; // @[Mux.scala 19:72:@1746.4]
  assign _T_1748 = _T_1747 | _T_1662; // @[Mux.scala 19:72:@1747.4]
  assign _T_1749 = _T_1748 | _T_1664; // @[Mux.scala 19:72:@1748.4]
  assign _T_1750 = _T_1749 | _T_1666; // @[Mux.scala 19:72:@1749.4]
  assign _T_1751 = _T_1750 | _T_1668; // @[Mux.scala 19:72:@1750.4]
  assign _T_1752 = _T_1751 | _T_1670; // @[Mux.scala 19:72:@1751.4]
  assign _T_1753 = _T_1752 | _T_1672; // @[Mux.scala 19:72:@1752.4]
  assign _T_1754 = _T_1753 | _T_1674; // @[Mux.scala 19:72:@1753.4]
  assign _T_1755 = _T_1754 | _T_1676; // @[Mux.scala 19:72:@1754.4]
  assign _T_1756 = _T_1755 | _T_1678; // @[Mux.scala 19:72:@1755.4]
  assign _T_1757 = _T_1756 | _T_1680; // @[Mux.scala 19:72:@1756.4]
  assign _T_1758 = _T_1757 | _T_1682; // @[Mux.scala 19:72:@1757.4]
  assign _T_1759 = _T_1758 | _T_1684; // @[Mux.scala 19:72:@1758.4]
  assign _T_1760 = _T_1759 | _T_1686; // @[Mux.scala 19:72:@1759.4]
  assign _T_1761 = _T_1760 | _T_1688; // @[Mux.scala 19:72:@1760.4]
  assign _T_1762 = _T_1761 | _T_1690; // @[Mux.scala 19:72:@1761.4]
  assign _T_1763 = _T_1762 | _T_1692; // @[Mux.scala 19:72:@1762.4]
  assign _T_1764 = _T_1763 | _T_1694; // @[Mux.scala 19:72:@1763.4]
  assign _T_1765 = _T_1764 | _T_1696; // @[Mux.scala 19:72:@1764.4]
  assign _T_1766 = _T_1765 | _T_1698; // @[Mux.scala 19:72:@1765.4]
  assign _T_1767 = _T_1766 | _T_1700; // @[Mux.scala 19:72:@1766.4]
  assign _T_1768 = _T_1767 | _T_1702; // @[Mux.scala 19:72:@1767.4]
  assign _T_1769 = _T_1768 | _T_1704; // @[Mux.scala 19:72:@1768.4]
  assign _T_1770 = _T_1769 | _T_1706; // @[Mux.scala 19:72:@1769.4]
  assign feedback_h_count = _T_1770 | _T_1708; // @[Mux.scala 19:72:@1770.4]
  assign _T_1776 = feedback_lookup != 64'h0; // @[BTB.scala 172:30:@1776.4]
  assign _T_1777 = feedback_lookup[63:32]; // @[OneHot.scala 26:18:@1777.4]
  assign _T_1778 = feedback_lookup[31:0]; // @[OneHot.scala 27:18:@1778.4]
  assign _T_1780 = _T_1777 != 32'h0; // @[OneHot.scala 28:14:@1779.4]
  assign _T_1781 = _T_1777 | _T_1778; // @[OneHot.scala 28:28:@1780.4]
  assign _T_1782 = _T_1781[31:16]; // @[OneHot.scala 26:18:@1781.4]
  assign _T_1783 = _T_1781[15:0]; // @[OneHot.scala 27:18:@1782.4]
  assign _T_1785 = _T_1782 != 16'h0; // @[OneHot.scala 28:14:@1783.4]
  assign _T_1786 = _T_1782 | _T_1783; // @[OneHot.scala 28:28:@1784.4]
  assign _T_1787 = _T_1786[15:8]; // @[OneHot.scala 26:18:@1785.4]
  assign _T_1788 = _T_1786[7:0]; // @[OneHot.scala 27:18:@1786.4]
  assign _T_1790 = _T_1787 != 8'h0; // @[OneHot.scala 28:14:@1787.4]
  assign _T_1791 = _T_1787 | _T_1788; // @[OneHot.scala 28:28:@1788.4]
  assign _T_1792 = _T_1791[7:4]; // @[OneHot.scala 26:18:@1789.4]
  assign _T_1793 = _T_1791[3:0]; // @[OneHot.scala 27:18:@1790.4]
  assign _T_1795 = _T_1792 != 4'h0; // @[OneHot.scala 28:14:@1791.4]
  assign _T_1796 = _T_1792 | _T_1793; // @[OneHot.scala 28:28:@1792.4]
  assign _T_1797 = _T_1796[3:2]; // @[OneHot.scala 26:18:@1793.4]
  assign _T_1798 = _T_1796[1:0]; // @[OneHot.scala 27:18:@1794.4]
  assign _T_1800 = _T_1797 != 2'h0; // @[OneHot.scala 28:14:@1795.4]
  assign _T_1801 = _T_1797 | _T_1798; // @[OneHot.scala 28:28:@1796.4]
  assign _T_1802 = _T_1801[1]; // @[CircuitMath.scala 30:8:@1797.4]
  assign _T_1807 = {_T_1780,_T_1785,_T_1790,_T_1795,_T_1800,_T_1802}; // @[Cat.scala 30:58:@1802.4]
  assign _T_1871 = ~ _T_409; // @[BTB.scala 181:26:@1866.4]
  assign _T_1873 = _T_1871 == 64'h0; // @[BTB.scala 181:26:@1867.4]
  assign _T_1938 = _T_1871[0]; // @[OneHot.scala 39:40:@1932.4]
  assign _T_1939 = _T_1871[1]; // @[OneHot.scala 39:40:@1933.4]
  assign _T_1940 = _T_1871[2]; // @[OneHot.scala 39:40:@1934.4]
  assign _T_1941 = _T_1871[3]; // @[OneHot.scala 39:40:@1935.4]
  assign _T_1942 = _T_1871[4]; // @[OneHot.scala 39:40:@1936.4]
  assign _T_1943 = _T_1871[5]; // @[OneHot.scala 39:40:@1937.4]
  assign _T_1944 = _T_1871[6]; // @[OneHot.scala 39:40:@1938.4]
  assign _T_1945 = _T_1871[7]; // @[OneHot.scala 39:40:@1939.4]
  assign _T_1946 = _T_1871[8]; // @[OneHot.scala 39:40:@1940.4]
  assign _T_1947 = _T_1871[9]; // @[OneHot.scala 39:40:@1941.4]
  assign _T_1948 = _T_1871[10]; // @[OneHot.scala 39:40:@1942.4]
  assign _T_1949 = _T_1871[11]; // @[OneHot.scala 39:40:@1943.4]
  assign _T_1950 = _T_1871[12]; // @[OneHot.scala 39:40:@1944.4]
  assign _T_1951 = _T_1871[13]; // @[OneHot.scala 39:40:@1945.4]
  assign _T_1952 = _T_1871[14]; // @[OneHot.scala 39:40:@1946.4]
  assign _T_1953 = _T_1871[15]; // @[OneHot.scala 39:40:@1947.4]
  assign _T_1954 = _T_1871[16]; // @[OneHot.scala 39:40:@1948.4]
  assign _T_1955 = _T_1871[17]; // @[OneHot.scala 39:40:@1949.4]
  assign _T_1956 = _T_1871[18]; // @[OneHot.scala 39:40:@1950.4]
  assign _T_1957 = _T_1871[19]; // @[OneHot.scala 39:40:@1951.4]
  assign _T_1958 = _T_1871[20]; // @[OneHot.scala 39:40:@1952.4]
  assign _T_1959 = _T_1871[21]; // @[OneHot.scala 39:40:@1953.4]
  assign _T_1960 = _T_1871[22]; // @[OneHot.scala 39:40:@1954.4]
  assign _T_1961 = _T_1871[23]; // @[OneHot.scala 39:40:@1955.4]
  assign _T_1962 = _T_1871[24]; // @[OneHot.scala 39:40:@1956.4]
  assign _T_1963 = _T_1871[25]; // @[OneHot.scala 39:40:@1957.4]
  assign _T_1964 = _T_1871[26]; // @[OneHot.scala 39:40:@1958.4]
  assign _T_1965 = _T_1871[27]; // @[OneHot.scala 39:40:@1959.4]
  assign _T_1966 = _T_1871[28]; // @[OneHot.scala 39:40:@1960.4]
  assign _T_1967 = _T_1871[29]; // @[OneHot.scala 39:40:@1961.4]
  assign _T_1968 = _T_1871[30]; // @[OneHot.scala 39:40:@1962.4]
  assign _T_1969 = _T_1871[31]; // @[OneHot.scala 39:40:@1963.4]
  assign _T_1970 = _T_1871[32]; // @[OneHot.scala 39:40:@1964.4]
  assign _T_1971 = _T_1871[33]; // @[OneHot.scala 39:40:@1965.4]
  assign _T_1972 = _T_1871[34]; // @[OneHot.scala 39:40:@1966.4]
  assign _T_1973 = _T_1871[35]; // @[OneHot.scala 39:40:@1967.4]
  assign _T_1974 = _T_1871[36]; // @[OneHot.scala 39:40:@1968.4]
  assign _T_1975 = _T_1871[37]; // @[OneHot.scala 39:40:@1969.4]
  assign _T_1976 = _T_1871[38]; // @[OneHot.scala 39:40:@1970.4]
  assign _T_1977 = _T_1871[39]; // @[OneHot.scala 39:40:@1971.4]
  assign _T_1978 = _T_1871[40]; // @[OneHot.scala 39:40:@1972.4]
  assign _T_1979 = _T_1871[41]; // @[OneHot.scala 39:40:@1973.4]
  assign _T_1980 = _T_1871[42]; // @[OneHot.scala 39:40:@1974.4]
  assign _T_1981 = _T_1871[43]; // @[OneHot.scala 39:40:@1975.4]
  assign _T_1982 = _T_1871[44]; // @[OneHot.scala 39:40:@1976.4]
  assign _T_1983 = _T_1871[45]; // @[OneHot.scala 39:40:@1977.4]
  assign _T_1984 = _T_1871[46]; // @[OneHot.scala 39:40:@1978.4]
  assign _T_1985 = _T_1871[47]; // @[OneHot.scala 39:40:@1979.4]
  assign _T_1986 = _T_1871[48]; // @[OneHot.scala 39:40:@1980.4]
  assign _T_1987 = _T_1871[49]; // @[OneHot.scala 39:40:@1981.4]
  assign _T_1988 = _T_1871[50]; // @[OneHot.scala 39:40:@1982.4]
  assign _T_1989 = _T_1871[51]; // @[OneHot.scala 39:40:@1983.4]
  assign _T_1990 = _T_1871[52]; // @[OneHot.scala 39:40:@1984.4]
  assign _T_1991 = _T_1871[53]; // @[OneHot.scala 39:40:@1985.4]
  assign _T_1992 = _T_1871[54]; // @[OneHot.scala 39:40:@1986.4]
  assign _T_1993 = _T_1871[55]; // @[OneHot.scala 39:40:@1987.4]
  assign _T_1994 = _T_1871[56]; // @[OneHot.scala 39:40:@1988.4]
  assign _T_1995 = _T_1871[57]; // @[OneHot.scala 39:40:@1989.4]
  assign _T_1996 = _T_1871[58]; // @[OneHot.scala 39:40:@1990.4]
  assign _T_1997 = _T_1871[59]; // @[OneHot.scala 39:40:@1991.4]
  assign _T_1998 = _T_1871[60]; // @[OneHot.scala 39:40:@1992.4]
  assign _T_1999 = _T_1871[61]; // @[OneHot.scala 39:40:@1993.4]
  assign _T_2000 = _T_1871[62]; // @[OneHot.scala 39:40:@1994.4]
  assign _T_2066 = _T_2000 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@1996.4]
  assign _T_2067 = _T_1999 ? 6'h3d : _T_2066; // @[Mux.scala 31:69:@1997.4]
  assign _T_2068 = _T_1998 ? 6'h3c : _T_2067; // @[Mux.scala 31:69:@1998.4]
  assign _T_2069 = _T_1997 ? 6'h3b : _T_2068; // @[Mux.scala 31:69:@1999.4]
  assign _T_2070 = _T_1996 ? 6'h3a : _T_2069; // @[Mux.scala 31:69:@2000.4]
  assign _T_2071 = _T_1995 ? 6'h39 : _T_2070; // @[Mux.scala 31:69:@2001.4]
  assign _T_2072 = _T_1994 ? 6'h38 : _T_2071; // @[Mux.scala 31:69:@2002.4]
  assign _T_2073 = _T_1993 ? 6'h37 : _T_2072; // @[Mux.scala 31:69:@2003.4]
  assign _T_2074 = _T_1992 ? 6'h36 : _T_2073; // @[Mux.scala 31:69:@2004.4]
  assign _T_2075 = _T_1991 ? 6'h35 : _T_2074; // @[Mux.scala 31:69:@2005.4]
  assign _T_2076 = _T_1990 ? 6'h34 : _T_2075; // @[Mux.scala 31:69:@2006.4]
  assign _T_2077 = _T_1989 ? 6'h33 : _T_2076; // @[Mux.scala 31:69:@2007.4]
  assign _T_2078 = _T_1988 ? 6'h32 : _T_2077; // @[Mux.scala 31:69:@2008.4]
  assign _T_2079 = _T_1987 ? 6'h31 : _T_2078; // @[Mux.scala 31:69:@2009.4]
  assign _T_2080 = _T_1986 ? 6'h30 : _T_2079; // @[Mux.scala 31:69:@2010.4]
  assign _T_2081 = _T_1985 ? 6'h2f : _T_2080; // @[Mux.scala 31:69:@2011.4]
  assign _T_2082 = _T_1984 ? 6'h2e : _T_2081; // @[Mux.scala 31:69:@2012.4]
  assign _T_2083 = _T_1983 ? 6'h2d : _T_2082; // @[Mux.scala 31:69:@2013.4]
  assign _T_2084 = _T_1982 ? 6'h2c : _T_2083; // @[Mux.scala 31:69:@2014.4]
  assign _T_2085 = _T_1981 ? 6'h2b : _T_2084; // @[Mux.scala 31:69:@2015.4]
  assign _T_2086 = _T_1980 ? 6'h2a : _T_2085; // @[Mux.scala 31:69:@2016.4]
  assign _T_2087 = _T_1979 ? 6'h29 : _T_2086; // @[Mux.scala 31:69:@2017.4]
  assign _T_2088 = _T_1978 ? 6'h28 : _T_2087; // @[Mux.scala 31:69:@2018.4]
  assign _T_2089 = _T_1977 ? 6'h27 : _T_2088; // @[Mux.scala 31:69:@2019.4]
  assign _T_2090 = _T_1976 ? 6'h26 : _T_2089; // @[Mux.scala 31:69:@2020.4]
  assign _T_2091 = _T_1975 ? 6'h25 : _T_2090; // @[Mux.scala 31:69:@2021.4]
  assign _T_2092 = _T_1974 ? 6'h24 : _T_2091; // @[Mux.scala 31:69:@2022.4]
  assign _T_2093 = _T_1973 ? 6'h23 : _T_2092; // @[Mux.scala 31:69:@2023.4]
  assign _T_2094 = _T_1972 ? 6'h22 : _T_2093; // @[Mux.scala 31:69:@2024.4]
  assign _T_2095 = _T_1971 ? 6'h21 : _T_2094; // @[Mux.scala 31:69:@2025.4]
  assign _T_2096 = _T_1970 ? 6'h20 : _T_2095; // @[Mux.scala 31:69:@2026.4]
  assign _T_2097 = _T_1969 ? 6'h1f : _T_2096; // @[Mux.scala 31:69:@2027.4]
  assign _T_2098 = _T_1968 ? 6'h1e : _T_2097; // @[Mux.scala 31:69:@2028.4]
  assign _T_2099 = _T_1967 ? 6'h1d : _T_2098; // @[Mux.scala 31:69:@2029.4]
  assign _T_2100 = _T_1966 ? 6'h1c : _T_2099; // @[Mux.scala 31:69:@2030.4]
  assign _T_2101 = _T_1965 ? 6'h1b : _T_2100; // @[Mux.scala 31:69:@2031.4]
  assign _T_2102 = _T_1964 ? 6'h1a : _T_2101; // @[Mux.scala 31:69:@2032.4]
  assign _T_2103 = _T_1963 ? 6'h19 : _T_2102; // @[Mux.scala 31:69:@2033.4]
  assign _T_2104 = _T_1962 ? 6'h18 : _T_2103; // @[Mux.scala 31:69:@2034.4]
  assign _T_2105 = _T_1961 ? 6'h17 : _T_2104; // @[Mux.scala 31:69:@2035.4]
  assign _T_2106 = _T_1960 ? 6'h16 : _T_2105; // @[Mux.scala 31:69:@2036.4]
  assign _T_2107 = _T_1959 ? 6'h15 : _T_2106; // @[Mux.scala 31:69:@2037.4]
  assign _T_2108 = _T_1958 ? 6'h14 : _T_2107; // @[Mux.scala 31:69:@2038.4]
  assign _T_2109 = _T_1957 ? 6'h13 : _T_2108; // @[Mux.scala 31:69:@2039.4]
  assign _T_2110 = _T_1956 ? 6'h12 : _T_2109; // @[Mux.scala 31:69:@2040.4]
  assign _T_2111 = _T_1955 ? 6'h11 : _T_2110; // @[Mux.scala 31:69:@2041.4]
  assign _T_2112 = _T_1954 ? 6'h10 : _T_2111; // @[Mux.scala 31:69:@2042.4]
  assign _T_2113 = _T_1953 ? 6'hf : _T_2112; // @[Mux.scala 31:69:@2043.4]
  assign _T_2114 = _T_1952 ? 6'he : _T_2113; // @[Mux.scala 31:69:@2044.4]
  assign _T_2115 = _T_1951 ? 6'hd : _T_2114; // @[Mux.scala 31:69:@2045.4]
  assign _T_2116 = _T_1950 ? 6'hc : _T_2115; // @[Mux.scala 31:69:@2046.4]
  assign _T_2117 = _T_1949 ? 6'hb : _T_2116; // @[Mux.scala 31:69:@2047.4]
  assign _T_2118 = _T_1948 ? 6'ha : _T_2117; // @[Mux.scala 31:69:@2048.4]
  assign _T_2119 = _T_1947 ? 6'h9 : _T_2118; // @[Mux.scala 31:69:@2049.4]
  assign _T_2120 = _T_1946 ? 6'h8 : _T_2119; // @[Mux.scala 31:69:@2050.4]
  assign _T_2121 = _T_1945 ? 6'h7 : _T_2120; // @[Mux.scala 31:69:@2051.4]
  assign _T_2122 = _T_1944 ? 6'h6 : _T_2121; // @[Mux.scala 31:69:@2052.4]
  assign _T_2123 = _T_1943 ? 6'h5 : _T_2122; // @[Mux.scala 31:69:@2053.4]
  assign _T_2124 = _T_1942 ? 6'h4 : _T_2123; // @[Mux.scala 31:69:@2054.4]
  assign _T_2125 = _T_1941 ? 6'h3 : _T_2124; // @[Mux.scala 31:69:@2055.4]
  assign _T_2126 = _T_1940 ? 6'h2 : _T_2125; // @[Mux.scala 31:69:@2056.4]
  assign _T_2127 = _T_1939 ? 6'h1 : _T_2126; // @[Mux.scala 31:69:@2057.4]
  assign _T_2128 = _T_1938 ? 6'h0 : _T_2127; // @[Mux.scala 31:69:@2058.4]
  assign _T_2129 = _T_1873 ? fb_reg_lfsr : _T_2128; // @[BTB.scala 181:8:@2059.4]
  assign feedback_idx = _T_1776 ? _T_1807 : _T_2129; // @[BTB.scala 180:22:@2060.4]
  assign _GEN_7 = 6'h0 == feedback_idx ? 1'h1 : btb_valid_0; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_8 = 6'h1 == feedback_idx ? 1'h1 : btb_valid_1; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_9 = 6'h2 == feedback_idx ? 1'h1 : btb_valid_2; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_10 = 6'h3 == feedback_idx ? 1'h1 : btb_valid_3; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_11 = 6'h4 == feedback_idx ? 1'h1 : btb_valid_4; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_12 = 6'h5 == feedback_idx ? 1'h1 : btb_valid_5; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_13 = 6'h6 == feedback_idx ? 1'h1 : btb_valid_6; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_14 = 6'h7 == feedback_idx ? 1'h1 : btb_valid_7; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_15 = 6'h8 == feedback_idx ? 1'h1 : btb_valid_8; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_16 = 6'h9 == feedback_idx ? 1'h1 : btb_valid_9; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_17 = 6'ha == feedback_idx ? 1'h1 : btb_valid_10; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_18 = 6'hb == feedback_idx ? 1'h1 : btb_valid_11; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_19 = 6'hc == feedback_idx ? 1'h1 : btb_valid_12; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_20 = 6'hd == feedback_idx ? 1'h1 : btb_valid_13; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_21 = 6'he == feedback_idx ? 1'h1 : btb_valid_14; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_22 = 6'hf == feedback_idx ? 1'h1 : btb_valid_15; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_23 = 6'h10 == feedback_idx ? 1'h1 : btb_valid_16; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_24 = 6'h11 == feedback_idx ? 1'h1 : btb_valid_17; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_25 = 6'h12 == feedback_idx ? 1'h1 : btb_valid_18; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_26 = 6'h13 == feedback_idx ? 1'h1 : btb_valid_19; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_27 = 6'h14 == feedback_idx ? 1'h1 : btb_valid_20; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_28 = 6'h15 == feedback_idx ? 1'h1 : btb_valid_21; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_29 = 6'h16 == feedback_idx ? 1'h1 : btb_valid_22; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_30 = 6'h17 == feedback_idx ? 1'h1 : btb_valid_23; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_31 = 6'h18 == feedback_idx ? 1'h1 : btb_valid_24; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_32 = 6'h19 == feedback_idx ? 1'h1 : btb_valid_25; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_33 = 6'h1a == feedback_idx ? 1'h1 : btb_valid_26; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_34 = 6'h1b == feedback_idx ? 1'h1 : btb_valid_27; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_35 = 6'h1c == feedback_idx ? 1'h1 : btb_valid_28; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_36 = 6'h1d == feedback_idx ? 1'h1 : btb_valid_29; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_37 = 6'h1e == feedback_idx ? 1'h1 : btb_valid_30; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_38 = 6'h1f == feedback_idx ? 1'h1 : btb_valid_31; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_39 = 6'h20 == feedback_idx ? 1'h1 : btb_valid_32; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_40 = 6'h21 == feedback_idx ? 1'h1 : btb_valid_33; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_41 = 6'h22 == feedback_idx ? 1'h1 : btb_valid_34; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_42 = 6'h23 == feedback_idx ? 1'h1 : btb_valid_35; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_43 = 6'h24 == feedback_idx ? 1'h1 : btb_valid_36; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_44 = 6'h25 == feedback_idx ? 1'h1 : btb_valid_37; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_45 = 6'h26 == feedback_idx ? 1'h1 : btb_valid_38; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_46 = 6'h27 == feedback_idx ? 1'h1 : btb_valid_39; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_47 = 6'h28 == feedback_idx ? 1'h1 : btb_valid_40; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_48 = 6'h29 == feedback_idx ? 1'h1 : btb_valid_41; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_49 = 6'h2a == feedback_idx ? 1'h1 : btb_valid_42; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_50 = 6'h2b == feedback_idx ? 1'h1 : btb_valid_43; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_51 = 6'h2c == feedback_idx ? 1'h1 : btb_valid_44; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_52 = 6'h2d == feedback_idx ? 1'h1 : btb_valid_45; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_53 = 6'h2e == feedback_idx ? 1'h1 : btb_valid_46; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_54 = 6'h2f == feedback_idx ? 1'h1 : btb_valid_47; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_55 = 6'h30 == feedback_idx ? 1'h1 : btb_valid_48; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_56 = 6'h31 == feedback_idx ? 1'h1 : btb_valid_49; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_57 = 6'h32 == feedback_idx ? 1'h1 : btb_valid_50; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_58 = 6'h33 == feedback_idx ? 1'h1 : btb_valid_51; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_59 = 6'h34 == feedback_idx ? 1'h1 : btb_valid_52; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_60 = 6'h35 == feedback_idx ? 1'h1 : btb_valid_53; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_61 = 6'h36 == feedback_idx ? 1'h1 : btb_valid_54; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_62 = 6'h37 == feedback_idx ? 1'h1 : btb_valid_55; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_63 = 6'h38 == feedback_idx ? 1'h1 : btb_valid_56; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_64 = 6'h39 == feedback_idx ? 1'h1 : btb_valid_57; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_65 = 6'h3a == feedback_idx ? 1'h1 : btb_valid_58; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_66 = 6'h3b == feedback_idx ? 1'h1 : btb_valid_59; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_67 = 6'h3c == feedback_idx ? 1'h1 : btb_valid_60; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_68 = 6'h3d == feedback_idx ? 1'h1 : btb_valid_61; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_69 = 6'h3e == feedback_idx ? 1'h1 : btb_valid_62; // @[BTB.scala 185:32:@2064.8]
  assign _GEN_70 = 6'h3f == feedback_idx ? 1'h1 : btb_valid_63; // @[BTB.scala 185:32:@2064.8]
  assign _T_2135 = fb_reg_btb_type == 2'h2; // @[BTB.scala 187:51:@2069.10]
  assign _GEN_71 = 6'h0 == feedback_idx ? _T_2135 : btb_valid_0; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_72 = 6'h1 == feedback_idx ? _T_2135 : btb_valid_1; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_73 = 6'h2 == feedback_idx ? _T_2135 : btb_valid_2; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_74 = 6'h3 == feedback_idx ? _T_2135 : btb_valid_3; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_75 = 6'h4 == feedback_idx ? _T_2135 : btb_valid_4; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_76 = 6'h5 == feedback_idx ? _T_2135 : btb_valid_5; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_77 = 6'h6 == feedback_idx ? _T_2135 : btb_valid_6; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_78 = 6'h7 == feedback_idx ? _T_2135 : btb_valid_7; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_79 = 6'h8 == feedback_idx ? _T_2135 : btb_valid_8; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_80 = 6'h9 == feedback_idx ? _T_2135 : btb_valid_9; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_81 = 6'ha == feedback_idx ? _T_2135 : btb_valid_10; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_82 = 6'hb == feedback_idx ? _T_2135 : btb_valid_11; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_83 = 6'hc == feedback_idx ? _T_2135 : btb_valid_12; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_84 = 6'hd == feedback_idx ? _T_2135 : btb_valid_13; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_85 = 6'he == feedback_idx ? _T_2135 : btb_valid_14; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_86 = 6'hf == feedback_idx ? _T_2135 : btb_valid_15; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_87 = 6'h10 == feedback_idx ? _T_2135 : btb_valid_16; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_88 = 6'h11 == feedback_idx ? _T_2135 : btb_valid_17; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_89 = 6'h12 == feedback_idx ? _T_2135 : btb_valid_18; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_90 = 6'h13 == feedback_idx ? _T_2135 : btb_valid_19; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_91 = 6'h14 == feedback_idx ? _T_2135 : btb_valid_20; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_92 = 6'h15 == feedback_idx ? _T_2135 : btb_valid_21; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_93 = 6'h16 == feedback_idx ? _T_2135 : btb_valid_22; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_94 = 6'h17 == feedback_idx ? _T_2135 : btb_valid_23; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_95 = 6'h18 == feedback_idx ? _T_2135 : btb_valid_24; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_96 = 6'h19 == feedback_idx ? _T_2135 : btb_valid_25; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_97 = 6'h1a == feedback_idx ? _T_2135 : btb_valid_26; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_98 = 6'h1b == feedback_idx ? _T_2135 : btb_valid_27; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_99 = 6'h1c == feedback_idx ? _T_2135 : btb_valid_28; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_100 = 6'h1d == feedback_idx ? _T_2135 : btb_valid_29; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_101 = 6'h1e == feedback_idx ? _T_2135 : btb_valid_30; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_102 = 6'h1f == feedback_idx ? _T_2135 : btb_valid_31; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_103 = 6'h20 == feedback_idx ? _T_2135 : btb_valid_32; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_104 = 6'h21 == feedback_idx ? _T_2135 : btb_valid_33; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_105 = 6'h22 == feedback_idx ? _T_2135 : btb_valid_34; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_106 = 6'h23 == feedback_idx ? _T_2135 : btb_valid_35; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_107 = 6'h24 == feedback_idx ? _T_2135 : btb_valid_36; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_108 = 6'h25 == feedback_idx ? _T_2135 : btb_valid_37; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_109 = 6'h26 == feedback_idx ? _T_2135 : btb_valid_38; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_110 = 6'h27 == feedback_idx ? _T_2135 : btb_valid_39; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_111 = 6'h28 == feedback_idx ? _T_2135 : btb_valid_40; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_112 = 6'h29 == feedback_idx ? _T_2135 : btb_valid_41; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_113 = 6'h2a == feedback_idx ? _T_2135 : btb_valid_42; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_114 = 6'h2b == feedback_idx ? _T_2135 : btb_valid_43; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_115 = 6'h2c == feedback_idx ? _T_2135 : btb_valid_44; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_116 = 6'h2d == feedback_idx ? _T_2135 : btb_valid_45; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_117 = 6'h2e == feedback_idx ? _T_2135 : btb_valid_46; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_118 = 6'h2f == feedback_idx ? _T_2135 : btb_valid_47; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_119 = 6'h30 == feedback_idx ? _T_2135 : btb_valid_48; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_120 = 6'h31 == feedback_idx ? _T_2135 : btb_valid_49; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_121 = 6'h32 == feedback_idx ? _T_2135 : btb_valid_50; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_122 = 6'h33 == feedback_idx ? _T_2135 : btb_valid_51; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_123 = 6'h34 == feedback_idx ? _T_2135 : btb_valid_52; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_124 = 6'h35 == feedback_idx ? _T_2135 : btb_valid_53; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_125 = 6'h36 == feedback_idx ? _T_2135 : btb_valid_54; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_126 = 6'h37 == feedback_idx ? _T_2135 : btb_valid_55; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_127 = 6'h38 == feedback_idx ? _T_2135 : btb_valid_56; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_128 = 6'h39 == feedback_idx ? _T_2135 : btb_valid_57; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_129 = 6'h3a == feedback_idx ? _T_2135 : btb_valid_58; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_130 = 6'h3b == feedback_idx ? _T_2135 : btb_valid_59; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_131 = 6'h3c == feedback_idx ? _T_2135 : btb_valid_60; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_132 = 6'h3d == feedback_idx ? _T_2135 : btb_valid_61; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_133 = 6'h3e == feedback_idx ? _T_2135 : btb_valid_62; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_134 = 6'h3f == feedback_idx ? _T_2135 : btb_valid_63; // @[BTB.scala 187:32:@2070.10]
  assign _GEN_135 = _T_1776 ? _GEN_71 : btb_valid_0; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_136 = _T_1776 ? _GEN_72 : btb_valid_1; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_137 = _T_1776 ? _GEN_73 : btb_valid_2; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_138 = _T_1776 ? _GEN_74 : btb_valid_3; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_139 = _T_1776 ? _GEN_75 : btb_valid_4; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_140 = _T_1776 ? _GEN_76 : btb_valid_5; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_141 = _T_1776 ? _GEN_77 : btb_valid_6; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_142 = _T_1776 ? _GEN_78 : btb_valid_7; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_143 = _T_1776 ? _GEN_79 : btb_valid_8; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_144 = _T_1776 ? _GEN_80 : btb_valid_9; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_145 = _T_1776 ? _GEN_81 : btb_valid_10; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_146 = _T_1776 ? _GEN_82 : btb_valid_11; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_147 = _T_1776 ? _GEN_83 : btb_valid_12; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_148 = _T_1776 ? _GEN_84 : btb_valid_13; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_149 = _T_1776 ? _GEN_85 : btb_valid_14; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_150 = _T_1776 ? _GEN_86 : btb_valid_15; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_151 = _T_1776 ? _GEN_87 : btb_valid_16; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_152 = _T_1776 ? _GEN_88 : btb_valid_17; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_153 = _T_1776 ? _GEN_89 : btb_valid_18; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_154 = _T_1776 ? _GEN_90 : btb_valid_19; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_155 = _T_1776 ? _GEN_91 : btb_valid_20; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_156 = _T_1776 ? _GEN_92 : btb_valid_21; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_157 = _T_1776 ? _GEN_93 : btb_valid_22; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_158 = _T_1776 ? _GEN_94 : btb_valid_23; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_159 = _T_1776 ? _GEN_95 : btb_valid_24; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_160 = _T_1776 ? _GEN_96 : btb_valid_25; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_161 = _T_1776 ? _GEN_97 : btb_valid_26; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_162 = _T_1776 ? _GEN_98 : btb_valid_27; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_163 = _T_1776 ? _GEN_99 : btb_valid_28; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_164 = _T_1776 ? _GEN_100 : btb_valid_29; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_165 = _T_1776 ? _GEN_101 : btb_valid_30; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_166 = _T_1776 ? _GEN_102 : btb_valid_31; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_167 = _T_1776 ? _GEN_103 : btb_valid_32; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_168 = _T_1776 ? _GEN_104 : btb_valid_33; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_169 = _T_1776 ? _GEN_105 : btb_valid_34; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_170 = _T_1776 ? _GEN_106 : btb_valid_35; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_171 = _T_1776 ? _GEN_107 : btb_valid_36; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_172 = _T_1776 ? _GEN_108 : btb_valid_37; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_173 = _T_1776 ? _GEN_109 : btb_valid_38; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_174 = _T_1776 ? _GEN_110 : btb_valid_39; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_175 = _T_1776 ? _GEN_111 : btb_valid_40; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_176 = _T_1776 ? _GEN_112 : btb_valid_41; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_177 = _T_1776 ? _GEN_113 : btb_valid_42; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_178 = _T_1776 ? _GEN_114 : btb_valid_43; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_179 = _T_1776 ? _GEN_115 : btb_valid_44; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_180 = _T_1776 ? _GEN_116 : btb_valid_45; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_181 = _T_1776 ? _GEN_117 : btb_valid_46; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_182 = _T_1776 ? _GEN_118 : btb_valid_47; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_183 = _T_1776 ? _GEN_119 : btb_valid_48; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_184 = _T_1776 ? _GEN_120 : btb_valid_49; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_185 = _T_1776 ? _GEN_121 : btb_valid_50; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_186 = _T_1776 ? _GEN_122 : btb_valid_51; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_187 = _T_1776 ? _GEN_123 : btb_valid_52; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_188 = _T_1776 ? _GEN_124 : btb_valid_53; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_189 = _T_1776 ? _GEN_125 : btb_valid_54; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_190 = _T_1776 ? _GEN_126 : btb_valid_55; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_191 = _T_1776 ? _GEN_127 : btb_valid_56; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_192 = _T_1776 ? _GEN_128 : btb_valid_57; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_193 = _T_1776 ? _GEN_129 : btb_valid_58; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_194 = _T_1776 ? _GEN_130 : btb_valid_59; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_195 = _T_1776 ? _GEN_131 : btb_valid_60; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_196 = _T_1776 ? _GEN_132 : btb_valid_61; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_197 = _T_1776 ? _GEN_133 : btb_valid_62; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_198 = _T_1776 ? _GEN_134 : btb_valid_63; // @[BTB.scala 186:32:@2068.8]
  assign _GEN_199 = fb_reg_redirect ? _GEN_7 : _GEN_135; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_200 = fb_reg_redirect ? _GEN_8 : _GEN_136; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_201 = fb_reg_redirect ? _GEN_9 : _GEN_137; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_202 = fb_reg_redirect ? _GEN_10 : _GEN_138; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_203 = fb_reg_redirect ? _GEN_11 : _GEN_139; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_204 = fb_reg_redirect ? _GEN_12 : _GEN_140; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_205 = fb_reg_redirect ? _GEN_13 : _GEN_141; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_206 = fb_reg_redirect ? _GEN_14 : _GEN_142; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_207 = fb_reg_redirect ? _GEN_15 : _GEN_143; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_208 = fb_reg_redirect ? _GEN_16 : _GEN_144; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_209 = fb_reg_redirect ? _GEN_17 : _GEN_145; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_210 = fb_reg_redirect ? _GEN_18 : _GEN_146; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_211 = fb_reg_redirect ? _GEN_19 : _GEN_147; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_212 = fb_reg_redirect ? _GEN_20 : _GEN_148; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_213 = fb_reg_redirect ? _GEN_21 : _GEN_149; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_214 = fb_reg_redirect ? _GEN_22 : _GEN_150; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_215 = fb_reg_redirect ? _GEN_23 : _GEN_151; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_216 = fb_reg_redirect ? _GEN_24 : _GEN_152; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_217 = fb_reg_redirect ? _GEN_25 : _GEN_153; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_218 = fb_reg_redirect ? _GEN_26 : _GEN_154; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_219 = fb_reg_redirect ? _GEN_27 : _GEN_155; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_220 = fb_reg_redirect ? _GEN_28 : _GEN_156; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_221 = fb_reg_redirect ? _GEN_29 : _GEN_157; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_222 = fb_reg_redirect ? _GEN_30 : _GEN_158; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_223 = fb_reg_redirect ? _GEN_31 : _GEN_159; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_224 = fb_reg_redirect ? _GEN_32 : _GEN_160; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_225 = fb_reg_redirect ? _GEN_33 : _GEN_161; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_226 = fb_reg_redirect ? _GEN_34 : _GEN_162; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_227 = fb_reg_redirect ? _GEN_35 : _GEN_163; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_228 = fb_reg_redirect ? _GEN_36 : _GEN_164; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_229 = fb_reg_redirect ? _GEN_37 : _GEN_165; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_230 = fb_reg_redirect ? _GEN_38 : _GEN_166; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_231 = fb_reg_redirect ? _GEN_39 : _GEN_167; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_232 = fb_reg_redirect ? _GEN_40 : _GEN_168; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_233 = fb_reg_redirect ? _GEN_41 : _GEN_169; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_234 = fb_reg_redirect ? _GEN_42 : _GEN_170; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_235 = fb_reg_redirect ? _GEN_43 : _GEN_171; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_236 = fb_reg_redirect ? _GEN_44 : _GEN_172; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_237 = fb_reg_redirect ? _GEN_45 : _GEN_173; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_238 = fb_reg_redirect ? _GEN_46 : _GEN_174; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_239 = fb_reg_redirect ? _GEN_47 : _GEN_175; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_240 = fb_reg_redirect ? _GEN_48 : _GEN_176; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_241 = fb_reg_redirect ? _GEN_49 : _GEN_177; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_242 = fb_reg_redirect ? _GEN_50 : _GEN_178; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_243 = fb_reg_redirect ? _GEN_51 : _GEN_179; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_244 = fb_reg_redirect ? _GEN_52 : _GEN_180; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_245 = fb_reg_redirect ? _GEN_53 : _GEN_181; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_246 = fb_reg_redirect ? _GEN_54 : _GEN_182; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_247 = fb_reg_redirect ? _GEN_55 : _GEN_183; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_248 = fb_reg_redirect ? _GEN_56 : _GEN_184; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_249 = fb_reg_redirect ? _GEN_57 : _GEN_185; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_250 = fb_reg_redirect ? _GEN_58 : _GEN_186; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_251 = fb_reg_redirect ? _GEN_59 : _GEN_187; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_252 = fb_reg_redirect ? _GEN_60 : _GEN_188; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_253 = fb_reg_redirect ? _GEN_61 : _GEN_189; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_254 = fb_reg_redirect ? _GEN_62 : _GEN_190; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_255 = fb_reg_redirect ? _GEN_63 : _GEN_191; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_256 = fb_reg_redirect ? _GEN_64 : _GEN_192; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_257 = fb_reg_redirect ? _GEN_65 : _GEN_193; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_258 = fb_reg_redirect ? _GEN_66 : _GEN_194; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_259 = fb_reg_redirect ? _GEN_67 : _GEN_195; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_260 = fb_reg_redirect ? _GEN_68 : _GEN_196; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_261 = fb_reg_redirect ? _GEN_69 : _GEN_197; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_262 = fb_reg_redirect ? _GEN_70 : _GEN_198; // @[BTB.scala 184:28:@2063.6]
  assign _GEN_263 = 6'h0 == feedback_idx ? fb_reg_pc : btb_pc_0; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_264 = 6'h1 == feedback_idx ? fb_reg_pc : btb_pc_1; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_265 = 6'h2 == feedback_idx ? fb_reg_pc : btb_pc_2; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_266 = 6'h3 == feedback_idx ? fb_reg_pc : btb_pc_3; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_267 = 6'h4 == feedback_idx ? fb_reg_pc : btb_pc_4; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_268 = 6'h5 == feedback_idx ? fb_reg_pc : btb_pc_5; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_269 = 6'h6 == feedback_idx ? fb_reg_pc : btb_pc_6; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_270 = 6'h7 == feedback_idx ? fb_reg_pc : btb_pc_7; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_271 = 6'h8 == feedback_idx ? fb_reg_pc : btb_pc_8; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_272 = 6'h9 == feedback_idx ? fb_reg_pc : btb_pc_9; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_273 = 6'ha == feedback_idx ? fb_reg_pc : btb_pc_10; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_274 = 6'hb == feedback_idx ? fb_reg_pc : btb_pc_11; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_275 = 6'hc == feedback_idx ? fb_reg_pc : btb_pc_12; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_276 = 6'hd == feedback_idx ? fb_reg_pc : btb_pc_13; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_277 = 6'he == feedback_idx ? fb_reg_pc : btb_pc_14; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_278 = 6'hf == feedback_idx ? fb_reg_pc : btb_pc_15; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_279 = 6'h10 == feedback_idx ? fb_reg_pc : btb_pc_16; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_280 = 6'h11 == feedback_idx ? fb_reg_pc : btb_pc_17; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_281 = 6'h12 == feedback_idx ? fb_reg_pc : btb_pc_18; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_282 = 6'h13 == feedback_idx ? fb_reg_pc : btb_pc_19; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_283 = 6'h14 == feedback_idx ? fb_reg_pc : btb_pc_20; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_284 = 6'h15 == feedback_idx ? fb_reg_pc : btb_pc_21; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_285 = 6'h16 == feedback_idx ? fb_reg_pc : btb_pc_22; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_286 = 6'h17 == feedback_idx ? fb_reg_pc : btb_pc_23; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_287 = 6'h18 == feedback_idx ? fb_reg_pc : btb_pc_24; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_288 = 6'h19 == feedback_idx ? fb_reg_pc : btb_pc_25; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_289 = 6'h1a == feedback_idx ? fb_reg_pc : btb_pc_26; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_290 = 6'h1b == feedback_idx ? fb_reg_pc : btb_pc_27; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_291 = 6'h1c == feedback_idx ? fb_reg_pc : btb_pc_28; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_292 = 6'h1d == feedback_idx ? fb_reg_pc : btb_pc_29; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_293 = 6'h1e == feedback_idx ? fb_reg_pc : btb_pc_30; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_294 = 6'h1f == feedback_idx ? fb_reg_pc : btb_pc_31; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_295 = 6'h20 == feedback_idx ? fb_reg_pc : btb_pc_32; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_296 = 6'h21 == feedback_idx ? fb_reg_pc : btb_pc_33; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_297 = 6'h22 == feedback_idx ? fb_reg_pc : btb_pc_34; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_298 = 6'h23 == feedback_idx ? fb_reg_pc : btb_pc_35; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_299 = 6'h24 == feedback_idx ? fb_reg_pc : btb_pc_36; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_300 = 6'h25 == feedback_idx ? fb_reg_pc : btb_pc_37; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_301 = 6'h26 == feedback_idx ? fb_reg_pc : btb_pc_38; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_302 = 6'h27 == feedback_idx ? fb_reg_pc : btb_pc_39; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_303 = 6'h28 == feedback_idx ? fb_reg_pc : btb_pc_40; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_304 = 6'h29 == feedback_idx ? fb_reg_pc : btb_pc_41; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_305 = 6'h2a == feedback_idx ? fb_reg_pc : btb_pc_42; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_306 = 6'h2b == feedback_idx ? fb_reg_pc : btb_pc_43; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_307 = 6'h2c == feedback_idx ? fb_reg_pc : btb_pc_44; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_308 = 6'h2d == feedback_idx ? fb_reg_pc : btb_pc_45; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_309 = 6'h2e == feedback_idx ? fb_reg_pc : btb_pc_46; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_310 = 6'h2f == feedback_idx ? fb_reg_pc : btb_pc_47; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_311 = 6'h30 == feedback_idx ? fb_reg_pc : btb_pc_48; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_312 = 6'h31 == feedback_idx ? fb_reg_pc : btb_pc_49; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_313 = 6'h32 == feedback_idx ? fb_reg_pc : btb_pc_50; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_314 = 6'h33 == feedback_idx ? fb_reg_pc : btb_pc_51; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_315 = 6'h34 == feedback_idx ? fb_reg_pc : btb_pc_52; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_316 = 6'h35 == feedback_idx ? fb_reg_pc : btb_pc_53; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_317 = 6'h36 == feedback_idx ? fb_reg_pc : btb_pc_54; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_318 = 6'h37 == feedback_idx ? fb_reg_pc : btb_pc_55; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_319 = 6'h38 == feedback_idx ? fb_reg_pc : btb_pc_56; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_320 = 6'h39 == feedback_idx ? fb_reg_pc : btb_pc_57; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_321 = 6'h3a == feedback_idx ? fb_reg_pc : btb_pc_58; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_322 = 6'h3b == feedback_idx ? fb_reg_pc : btb_pc_59; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_323 = 6'h3c == feedback_idx ? fb_reg_pc : btb_pc_60; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_324 = 6'h3d == feedback_idx ? fb_reg_pc : btb_pc_61; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_325 = 6'h3e == feedback_idx ? fb_reg_pc : btb_pc_62; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_326 = 6'h3f == feedback_idx ? fb_reg_pc : btb_pc_63; // @[BTB.scala 190:33:@2073.8]
  assign _GEN_327 = 6'h0 == feedback_idx ? fb_reg_tgt : btb_tgt_0; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_328 = 6'h1 == feedback_idx ? fb_reg_tgt : btb_tgt_1; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_329 = 6'h2 == feedback_idx ? fb_reg_tgt : btb_tgt_2; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_330 = 6'h3 == feedback_idx ? fb_reg_tgt : btb_tgt_3; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_331 = 6'h4 == feedback_idx ? fb_reg_tgt : btb_tgt_4; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_332 = 6'h5 == feedback_idx ? fb_reg_tgt : btb_tgt_5; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_333 = 6'h6 == feedback_idx ? fb_reg_tgt : btb_tgt_6; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_334 = 6'h7 == feedback_idx ? fb_reg_tgt : btb_tgt_7; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_335 = 6'h8 == feedback_idx ? fb_reg_tgt : btb_tgt_8; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_336 = 6'h9 == feedback_idx ? fb_reg_tgt : btb_tgt_9; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_337 = 6'ha == feedback_idx ? fb_reg_tgt : btb_tgt_10; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_338 = 6'hb == feedback_idx ? fb_reg_tgt : btb_tgt_11; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_339 = 6'hc == feedback_idx ? fb_reg_tgt : btb_tgt_12; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_340 = 6'hd == feedback_idx ? fb_reg_tgt : btb_tgt_13; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_341 = 6'he == feedback_idx ? fb_reg_tgt : btb_tgt_14; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_342 = 6'hf == feedback_idx ? fb_reg_tgt : btb_tgt_15; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_343 = 6'h10 == feedback_idx ? fb_reg_tgt : btb_tgt_16; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_344 = 6'h11 == feedback_idx ? fb_reg_tgt : btb_tgt_17; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_345 = 6'h12 == feedback_idx ? fb_reg_tgt : btb_tgt_18; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_346 = 6'h13 == feedback_idx ? fb_reg_tgt : btb_tgt_19; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_347 = 6'h14 == feedback_idx ? fb_reg_tgt : btb_tgt_20; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_348 = 6'h15 == feedback_idx ? fb_reg_tgt : btb_tgt_21; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_349 = 6'h16 == feedback_idx ? fb_reg_tgt : btb_tgt_22; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_350 = 6'h17 == feedback_idx ? fb_reg_tgt : btb_tgt_23; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_351 = 6'h18 == feedback_idx ? fb_reg_tgt : btb_tgt_24; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_352 = 6'h19 == feedback_idx ? fb_reg_tgt : btb_tgt_25; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_353 = 6'h1a == feedback_idx ? fb_reg_tgt : btb_tgt_26; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_354 = 6'h1b == feedback_idx ? fb_reg_tgt : btb_tgt_27; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_355 = 6'h1c == feedback_idx ? fb_reg_tgt : btb_tgt_28; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_356 = 6'h1d == feedback_idx ? fb_reg_tgt : btb_tgt_29; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_357 = 6'h1e == feedback_idx ? fb_reg_tgt : btb_tgt_30; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_358 = 6'h1f == feedback_idx ? fb_reg_tgt : btb_tgt_31; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_359 = 6'h20 == feedback_idx ? fb_reg_tgt : btb_tgt_32; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_360 = 6'h21 == feedback_idx ? fb_reg_tgt : btb_tgt_33; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_361 = 6'h22 == feedback_idx ? fb_reg_tgt : btb_tgt_34; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_362 = 6'h23 == feedback_idx ? fb_reg_tgt : btb_tgt_35; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_363 = 6'h24 == feedback_idx ? fb_reg_tgt : btb_tgt_36; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_364 = 6'h25 == feedback_idx ? fb_reg_tgt : btb_tgt_37; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_365 = 6'h26 == feedback_idx ? fb_reg_tgt : btb_tgt_38; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_366 = 6'h27 == feedback_idx ? fb_reg_tgt : btb_tgt_39; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_367 = 6'h28 == feedback_idx ? fb_reg_tgt : btb_tgt_40; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_368 = 6'h29 == feedback_idx ? fb_reg_tgt : btb_tgt_41; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_369 = 6'h2a == feedback_idx ? fb_reg_tgt : btb_tgt_42; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_370 = 6'h2b == feedback_idx ? fb_reg_tgt : btb_tgt_43; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_371 = 6'h2c == feedback_idx ? fb_reg_tgt : btb_tgt_44; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_372 = 6'h2d == feedback_idx ? fb_reg_tgt : btb_tgt_45; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_373 = 6'h2e == feedback_idx ? fb_reg_tgt : btb_tgt_46; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_374 = 6'h2f == feedback_idx ? fb_reg_tgt : btb_tgt_47; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_375 = 6'h30 == feedback_idx ? fb_reg_tgt : btb_tgt_48; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_376 = 6'h31 == feedback_idx ? fb_reg_tgt : btb_tgt_49; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_377 = 6'h32 == feedback_idx ? fb_reg_tgt : btb_tgt_50; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_378 = 6'h33 == feedback_idx ? fb_reg_tgt : btb_tgt_51; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_379 = 6'h34 == feedback_idx ? fb_reg_tgt : btb_tgt_52; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_380 = 6'h35 == feedback_idx ? fb_reg_tgt : btb_tgt_53; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_381 = 6'h36 == feedback_idx ? fb_reg_tgt : btb_tgt_54; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_382 = 6'h37 == feedback_idx ? fb_reg_tgt : btb_tgt_55; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_383 = 6'h38 == feedback_idx ? fb_reg_tgt : btb_tgt_56; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_384 = 6'h39 == feedback_idx ? fb_reg_tgt : btb_tgt_57; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_385 = 6'h3a == feedback_idx ? fb_reg_tgt : btb_tgt_58; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_386 = 6'h3b == feedback_idx ? fb_reg_tgt : btb_tgt_59; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_387 = 6'h3c == feedback_idx ? fb_reg_tgt : btb_tgt_60; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_388 = 6'h3d == feedback_idx ? fb_reg_tgt : btb_tgt_61; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_389 = 6'h3e == feedback_idx ? fb_reg_tgt : btb_tgt_62; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_390 = 6'h3f == feedback_idx ? fb_reg_tgt : btb_tgt_63; // @[BTB.scala 191:33:@2074.8]
  assign _GEN_391 = 6'h0 == feedback_idx ? fb_reg_btb_type : btb_bj_type_0; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_392 = 6'h1 == feedback_idx ? fb_reg_btb_type : btb_bj_type_1; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_393 = 6'h2 == feedback_idx ? fb_reg_btb_type : btb_bj_type_2; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_394 = 6'h3 == feedback_idx ? fb_reg_btb_type : btb_bj_type_3; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_395 = 6'h4 == feedback_idx ? fb_reg_btb_type : btb_bj_type_4; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_396 = 6'h5 == feedback_idx ? fb_reg_btb_type : btb_bj_type_5; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_397 = 6'h6 == feedback_idx ? fb_reg_btb_type : btb_bj_type_6; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_398 = 6'h7 == feedback_idx ? fb_reg_btb_type : btb_bj_type_7; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_399 = 6'h8 == feedback_idx ? fb_reg_btb_type : btb_bj_type_8; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_400 = 6'h9 == feedback_idx ? fb_reg_btb_type : btb_bj_type_9; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_401 = 6'ha == feedback_idx ? fb_reg_btb_type : btb_bj_type_10; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_402 = 6'hb == feedback_idx ? fb_reg_btb_type : btb_bj_type_11; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_403 = 6'hc == feedback_idx ? fb_reg_btb_type : btb_bj_type_12; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_404 = 6'hd == feedback_idx ? fb_reg_btb_type : btb_bj_type_13; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_405 = 6'he == feedback_idx ? fb_reg_btb_type : btb_bj_type_14; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_406 = 6'hf == feedback_idx ? fb_reg_btb_type : btb_bj_type_15; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_407 = 6'h10 == feedback_idx ? fb_reg_btb_type : btb_bj_type_16; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_408 = 6'h11 == feedback_idx ? fb_reg_btb_type : btb_bj_type_17; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_409 = 6'h12 == feedback_idx ? fb_reg_btb_type : btb_bj_type_18; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_410 = 6'h13 == feedback_idx ? fb_reg_btb_type : btb_bj_type_19; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_411 = 6'h14 == feedback_idx ? fb_reg_btb_type : btb_bj_type_20; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_412 = 6'h15 == feedback_idx ? fb_reg_btb_type : btb_bj_type_21; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_413 = 6'h16 == feedback_idx ? fb_reg_btb_type : btb_bj_type_22; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_414 = 6'h17 == feedback_idx ? fb_reg_btb_type : btb_bj_type_23; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_415 = 6'h18 == feedback_idx ? fb_reg_btb_type : btb_bj_type_24; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_416 = 6'h19 == feedback_idx ? fb_reg_btb_type : btb_bj_type_25; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_417 = 6'h1a == feedback_idx ? fb_reg_btb_type : btb_bj_type_26; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_418 = 6'h1b == feedback_idx ? fb_reg_btb_type : btb_bj_type_27; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_419 = 6'h1c == feedback_idx ? fb_reg_btb_type : btb_bj_type_28; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_420 = 6'h1d == feedback_idx ? fb_reg_btb_type : btb_bj_type_29; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_421 = 6'h1e == feedback_idx ? fb_reg_btb_type : btb_bj_type_30; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_422 = 6'h1f == feedback_idx ? fb_reg_btb_type : btb_bj_type_31; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_423 = 6'h20 == feedback_idx ? fb_reg_btb_type : btb_bj_type_32; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_424 = 6'h21 == feedback_idx ? fb_reg_btb_type : btb_bj_type_33; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_425 = 6'h22 == feedback_idx ? fb_reg_btb_type : btb_bj_type_34; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_426 = 6'h23 == feedback_idx ? fb_reg_btb_type : btb_bj_type_35; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_427 = 6'h24 == feedback_idx ? fb_reg_btb_type : btb_bj_type_36; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_428 = 6'h25 == feedback_idx ? fb_reg_btb_type : btb_bj_type_37; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_429 = 6'h26 == feedback_idx ? fb_reg_btb_type : btb_bj_type_38; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_430 = 6'h27 == feedback_idx ? fb_reg_btb_type : btb_bj_type_39; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_431 = 6'h28 == feedback_idx ? fb_reg_btb_type : btb_bj_type_40; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_432 = 6'h29 == feedback_idx ? fb_reg_btb_type : btb_bj_type_41; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_433 = 6'h2a == feedback_idx ? fb_reg_btb_type : btb_bj_type_42; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_434 = 6'h2b == feedback_idx ? fb_reg_btb_type : btb_bj_type_43; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_435 = 6'h2c == feedback_idx ? fb_reg_btb_type : btb_bj_type_44; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_436 = 6'h2d == feedback_idx ? fb_reg_btb_type : btb_bj_type_45; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_437 = 6'h2e == feedback_idx ? fb_reg_btb_type : btb_bj_type_46; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_438 = 6'h2f == feedback_idx ? fb_reg_btb_type : btb_bj_type_47; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_439 = 6'h30 == feedback_idx ? fb_reg_btb_type : btb_bj_type_48; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_440 = 6'h31 == feedback_idx ? fb_reg_btb_type : btb_bj_type_49; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_441 = 6'h32 == feedback_idx ? fb_reg_btb_type : btb_bj_type_50; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_442 = 6'h33 == feedback_idx ? fb_reg_btb_type : btb_bj_type_51; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_443 = 6'h34 == feedback_idx ? fb_reg_btb_type : btb_bj_type_52; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_444 = 6'h35 == feedback_idx ? fb_reg_btb_type : btb_bj_type_53; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_445 = 6'h36 == feedback_idx ? fb_reg_btb_type : btb_bj_type_54; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_446 = 6'h37 == feedback_idx ? fb_reg_btb_type : btb_bj_type_55; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_447 = 6'h38 == feedback_idx ? fb_reg_btb_type : btb_bj_type_56; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_448 = 6'h39 == feedback_idx ? fb_reg_btb_type : btb_bj_type_57; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_449 = 6'h3a == feedback_idx ? fb_reg_btb_type : btb_bj_type_58; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_450 = 6'h3b == feedback_idx ? fb_reg_btb_type : btb_bj_type_59; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_451 = 6'h3c == feedback_idx ? fb_reg_btb_type : btb_bj_type_60; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_452 = 6'h3d == feedback_idx ? fb_reg_btb_type : btb_bj_type_61; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_453 = 6'h3e == feedback_idx ? fb_reg_btb_type : btb_bj_type_62; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_454 = 6'h3f == feedback_idx ? fb_reg_btb_type : btb_bj_type_63; // @[BTB.scala 192:33:@2075.8]
  assign _GEN_455 = fb_reg_redirect ? _GEN_263 : btb_pc_0; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_456 = fb_reg_redirect ? _GEN_264 : btb_pc_1; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_457 = fb_reg_redirect ? _GEN_265 : btb_pc_2; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_458 = fb_reg_redirect ? _GEN_266 : btb_pc_3; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_459 = fb_reg_redirect ? _GEN_267 : btb_pc_4; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_460 = fb_reg_redirect ? _GEN_268 : btb_pc_5; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_461 = fb_reg_redirect ? _GEN_269 : btb_pc_6; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_462 = fb_reg_redirect ? _GEN_270 : btb_pc_7; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_463 = fb_reg_redirect ? _GEN_271 : btb_pc_8; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_464 = fb_reg_redirect ? _GEN_272 : btb_pc_9; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_465 = fb_reg_redirect ? _GEN_273 : btb_pc_10; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_466 = fb_reg_redirect ? _GEN_274 : btb_pc_11; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_467 = fb_reg_redirect ? _GEN_275 : btb_pc_12; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_468 = fb_reg_redirect ? _GEN_276 : btb_pc_13; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_469 = fb_reg_redirect ? _GEN_277 : btb_pc_14; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_470 = fb_reg_redirect ? _GEN_278 : btb_pc_15; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_471 = fb_reg_redirect ? _GEN_279 : btb_pc_16; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_472 = fb_reg_redirect ? _GEN_280 : btb_pc_17; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_473 = fb_reg_redirect ? _GEN_281 : btb_pc_18; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_474 = fb_reg_redirect ? _GEN_282 : btb_pc_19; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_475 = fb_reg_redirect ? _GEN_283 : btb_pc_20; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_476 = fb_reg_redirect ? _GEN_284 : btb_pc_21; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_477 = fb_reg_redirect ? _GEN_285 : btb_pc_22; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_478 = fb_reg_redirect ? _GEN_286 : btb_pc_23; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_479 = fb_reg_redirect ? _GEN_287 : btb_pc_24; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_480 = fb_reg_redirect ? _GEN_288 : btb_pc_25; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_481 = fb_reg_redirect ? _GEN_289 : btb_pc_26; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_482 = fb_reg_redirect ? _GEN_290 : btb_pc_27; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_483 = fb_reg_redirect ? _GEN_291 : btb_pc_28; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_484 = fb_reg_redirect ? _GEN_292 : btb_pc_29; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_485 = fb_reg_redirect ? _GEN_293 : btb_pc_30; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_486 = fb_reg_redirect ? _GEN_294 : btb_pc_31; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_487 = fb_reg_redirect ? _GEN_295 : btb_pc_32; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_488 = fb_reg_redirect ? _GEN_296 : btb_pc_33; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_489 = fb_reg_redirect ? _GEN_297 : btb_pc_34; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_490 = fb_reg_redirect ? _GEN_298 : btb_pc_35; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_491 = fb_reg_redirect ? _GEN_299 : btb_pc_36; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_492 = fb_reg_redirect ? _GEN_300 : btb_pc_37; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_493 = fb_reg_redirect ? _GEN_301 : btb_pc_38; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_494 = fb_reg_redirect ? _GEN_302 : btb_pc_39; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_495 = fb_reg_redirect ? _GEN_303 : btb_pc_40; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_496 = fb_reg_redirect ? _GEN_304 : btb_pc_41; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_497 = fb_reg_redirect ? _GEN_305 : btb_pc_42; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_498 = fb_reg_redirect ? _GEN_306 : btb_pc_43; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_499 = fb_reg_redirect ? _GEN_307 : btb_pc_44; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_500 = fb_reg_redirect ? _GEN_308 : btb_pc_45; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_501 = fb_reg_redirect ? _GEN_309 : btb_pc_46; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_502 = fb_reg_redirect ? _GEN_310 : btb_pc_47; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_503 = fb_reg_redirect ? _GEN_311 : btb_pc_48; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_504 = fb_reg_redirect ? _GEN_312 : btb_pc_49; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_505 = fb_reg_redirect ? _GEN_313 : btb_pc_50; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_506 = fb_reg_redirect ? _GEN_314 : btb_pc_51; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_507 = fb_reg_redirect ? _GEN_315 : btb_pc_52; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_508 = fb_reg_redirect ? _GEN_316 : btb_pc_53; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_509 = fb_reg_redirect ? _GEN_317 : btb_pc_54; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_510 = fb_reg_redirect ? _GEN_318 : btb_pc_55; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_511 = fb_reg_redirect ? _GEN_319 : btb_pc_56; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_512 = fb_reg_redirect ? _GEN_320 : btb_pc_57; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_513 = fb_reg_redirect ? _GEN_321 : btb_pc_58; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_514 = fb_reg_redirect ? _GEN_322 : btb_pc_59; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_515 = fb_reg_redirect ? _GEN_323 : btb_pc_60; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_516 = fb_reg_redirect ? _GEN_324 : btb_pc_61; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_517 = fb_reg_redirect ? _GEN_325 : btb_pc_62; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_518 = fb_reg_redirect ? _GEN_326 : btb_pc_63; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_519 = fb_reg_redirect ? _GEN_327 : btb_tgt_0; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_520 = fb_reg_redirect ? _GEN_328 : btb_tgt_1; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_521 = fb_reg_redirect ? _GEN_329 : btb_tgt_2; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_522 = fb_reg_redirect ? _GEN_330 : btb_tgt_3; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_523 = fb_reg_redirect ? _GEN_331 : btb_tgt_4; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_524 = fb_reg_redirect ? _GEN_332 : btb_tgt_5; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_525 = fb_reg_redirect ? _GEN_333 : btb_tgt_6; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_526 = fb_reg_redirect ? _GEN_334 : btb_tgt_7; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_527 = fb_reg_redirect ? _GEN_335 : btb_tgt_8; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_528 = fb_reg_redirect ? _GEN_336 : btb_tgt_9; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_529 = fb_reg_redirect ? _GEN_337 : btb_tgt_10; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_530 = fb_reg_redirect ? _GEN_338 : btb_tgt_11; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_531 = fb_reg_redirect ? _GEN_339 : btb_tgt_12; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_532 = fb_reg_redirect ? _GEN_340 : btb_tgt_13; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_533 = fb_reg_redirect ? _GEN_341 : btb_tgt_14; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_534 = fb_reg_redirect ? _GEN_342 : btb_tgt_15; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_535 = fb_reg_redirect ? _GEN_343 : btb_tgt_16; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_536 = fb_reg_redirect ? _GEN_344 : btb_tgt_17; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_537 = fb_reg_redirect ? _GEN_345 : btb_tgt_18; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_538 = fb_reg_redirect ? _GEN_346 : btb_tgt_19; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_539 = fb_reg_redirect ? _GEN_347 : btb_tgt_20; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_540 = fb_reg_redirect ? _GEN_348 : btb_tgt_21; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_541 = fb_reg_redirect ? _GEN_349 : btb_tgt_22; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_542 = fb_reg_redirect ? _GEN_350 : btb_tgt_23; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_543 = fb_reg_redirect ? _GEN_351 : btb_tgt_24; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_544 = fb_reg_redirect ? _GEN_352 : btb_tgt_25; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_545 = fb_reg_redirect ? _GEN_353 : btb_tgt_26; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_546 = fb_reg_redirect ? _GEN_354 : btb_tgt_27; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_547 = fb_reg_redirect ? _GEN_355 : btb_tgt_28; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_548 = fb_reg_redirect ? _GEN_356 : btb_tgt_29; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_549 = fb_reg_redirect ? _GEN_357 : btb_tgt_30; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_550 = fb_reg_redirect ? _GEN_358 : btb_tgt_31; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_551 = fb_reg_redirect ? _GEN_359 : btb_tgt_32; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_552 = fb_reg_redirect ? _GEN_360 : btb_tgt_33; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_553 = fb_reg_redirect ? _GEN_361 : btb_tgt_34; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_554 = fb_reg_redirect ? _GEN_362 : btb_tgt_35; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_555 = fb_reg_redirect ? _GEN_363 : btb_tgt_36; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_556 = fb_reg_redirect ? _GEN_364 : btb_tgt_37; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_557 = fb_reg_redirect ? _GEN_365 : btb_tgt_38; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_558 = fb_reg_redirect ? _GEN_366 : btb_tgt_39; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_559 = fb_reg_redirect ? _GEN_367 : btb_tgt_40; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_560 = fb_reg_redirect ? _GEN_368 : btb_tgt_41; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_561 = fb_reg_redirect ? _GEN_369 : btb_tgt_42; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_562 = fb_reg_redirect ? _GEN_370 : btb_tgt_43; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_563 = fb_reg_redirect ? _GEN_371 : btb_tgt_44; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_564 = fb_reg_redirect ? _GEN_372 : btb_tgt_45; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_565 = fb_reg_redirect ? _GEN_373 : btb_tgt_46; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_566 = fb_reg_redirect ? _GEN_374 : btb_tgt_47; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_567 = fb_reg_redirect ? _GEN_375 : btb_tgt_48; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_568 = fb_reg_redirect ? _GEN_376 : btb_tgt_49; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_569 = fb_reg_redirect ? _GEN_377 : btb_tgt_50; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_570 = fb_reg_redirect ? _GEN_378 : btb_tgt_51; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_571 = fb_reg_redirect ? _GEN_379 : btb_tgt_52; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_572 = fb_reg_redirect ? _GEN_380 : btb_tgt_53; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_573 = fb_reg_redirect ? _GEN_381 : btb_tgt_54; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_574 = fb_reg_redirect ? _GEN_382 : btb_tgt_55; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_575 = fb_reg_redirect ? _GEN_383 : btb_tgt_56; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_576 = fb_reg_redirect ? _GEN_384 : btb_tgt_57; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_577 = fb_reg_redirect ? _GEN_385 : btb_tgt_58; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_578 = fb_reg_redirect ? _GEN_386 : btb_tgt_59; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_579 = fb_reg_redirect ? _GEN_387 : btb_tgt_60; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_580 = fb_reg_redirect ? _GEN_388 : btb_tgt_61; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_581 = fb_reg_redirect ? _GEN_389 : btb_tgt_62; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_582 = fb_reg_redirect ? _GEN_390 : btb_tgt_63; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_583 = fb_reg_redirect ? _GEN_391 : btb_bj_type_0; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_584 = fb_reg_redirect ? _GEN_392 : btb_bj_type_1; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_585 = fb_reg_redirect ? _GEN_393 : btb_bj_type_2; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_586 = fb_reg_redirect ? _GEN_394 : btb_bj_type_3; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_587 = fb_reg_redirect ? _GEN_395 : btb_bj_type_4; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_588 = fb_reg_redirect ? _GEN_396 : btb_bj_type_5; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_589 = fb_reg_redirect ? _GEN_397 : btb_bj_type_6; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_590 = fb_reg_redirect ? _GEN_398 : btb_bj_type_7; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_591 = fb_reg_redirect ? _GEN_399 : btb_bj_type_8; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_592 = fb_reg_redirect ? _GEN_400 : btb_bj_type_9; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_593 = fb_reg_redirect ? _GEN_401 : btb_bj_type_10; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_594 = fb_reg_redirect ? _GEN_402 : btb_bj_type_11; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_595 = fb_reg_redirect ? _GEN_403 : btb_bj_type_12; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_596 = fb_reg_redirect ? _GEN_404 : btb_bj_type_13; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_597 = fb_reg_redirect ? _GEN_405 : btb_bj_type_14; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_598 = fb_reg_redirect ? _GEN_406 : btb_bj_type_15; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_599 = fb_reg_redirect ? _GEN_407 : btb_bj_type_16; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_600 = fb_reg_redirect ? _GEN_408 : btb_bj_type_17; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_601 = fb_reg_redirect ? _GEN_409 : btb_bj_type_18; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_602 = fb_reg_redirect ? _GEN_410 : btb_bj_type_19; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_603 = fb_reg_redirect ? _GEN_411 : btb_bj_type_20; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_604 = fb_reg_redirect ? _GEN_412 : btb_bj_type_21; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_605 = fb_reg_redirect ? _GEN_413 : btb_bj_type_22; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_606 = fb_reg_redirect ? _GEN_414 : btb_bj_type_23; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_607 = fb_reg_redirect ? _GEN_415 : btb_bj_type_24; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_608 = fb_reg_redirect ? _GEN_416 : btb_bj_type_25; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_609 = fb_reg_redirect ? _GEN_417 : btb_bj_type_26; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_610 = fb_reg_redirect ? _GEN_418 : btb_bj_type_27; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_611 = fb_reg_redirect ? _GEN_419 : btb_bj_type_28; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_612 = fb_reg_redirect ? _GEN_420 : btb_bj_type_29; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_613 = fb_reg_redirect ? _GEN_421 : btb_bj_type_30; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_614 = fb_reg_redirect ? _GEN_422 : btb_bj_type_31; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_615 = fb_reg_redirect ? _GEN_423 : btb_bj_type_32; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_616 = fb_reg_redirect ? _GEN_424 : btb_bj_type_33; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_617 = fb_reg_redirect ? _GEN_425 : btb_bj_type_34; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_618 = fb_reg_redirect ? _GEN_426 : btb_bj_type_35; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_619 = fb_reg_redirect ? _GEN_427 : btb_bj_type_36; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_620 = fb_reg_redirect ? _GEN_428 : btb_bj_type_37; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_621 = fb_reg_redirect ? _GEN_429 : btb_bj_type_38; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_622 = fb_reg_redirect ? _GEN_430 : btb_bj_type_39; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_623 = fb_reg_redirect ? _GEN_431 : btb_bj_type_40; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_624 = fb_reg_redirect ? _GEN_432 : btb_bj_type_41; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_625 = fb_reg_redirect ? _GEN_433 : btb_bj_type_42; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_626 = fb_reg_redirect ? _GEN_434 : btb_bj_type_43; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_627 = fb_reg_redirect ? _GEN_435 : btb_bj_type_44; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_628 = fb_reg_redirect ? _GEN_436 : btb_bj_type_45; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_629 = fb_reg_redirect ? _GEN_437 : btb_bj_type_46; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_630 = fb_reg_redirect ? _GEN_438 : btb_bj_type_47; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_631 = fb_reg_redirect ? _GEN_439 : btb_bj_type_48; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_632 = fb_reg_redirect ? _GEN_440 : btb_bj_type_49; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_633 = fb_reg_redirect ? _GEN_441 : btb_bj_type_50; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_634 = fb_reg_redirect ? _GEN_442 : btb_bj_type_51; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_635 = fb_reg_redirect ? _GEN_443 : btb_bj_type_52; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_636 = fb_reg_redirect ? _GEN_444 : btb_bj_type_53; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_637 = fb_reg_redirect ? _GEN_445 : btb_bj_type_54; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_638 = fb_reg_redirect ? _GEN_446 : btb_bj_type_55; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_639 = fb_reg_redirect ? _GEN_447 : btb_bj_type_56; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_640 = fb_reg_redirect ? _GEN_448 : btb_bj_type_57; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_641 = fb_reg_redirect ? _GEN_449 : btb_bj_type_58; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_642 = fb_reg_redirect ? _GEN_450 : btb_bj_type_59; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_643 = fb_reg_redirect ? _GEN_451 : btb_bj_type_60; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_644 = fb_reg_redirect ? _GEN_452 : btb_bj_type_61; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_645 = fb_reg_redirect ? _GEN_453 : btb_bj_type_62; // @[BTB.scala 189:28:@2072.6]
  assign _GEN_646 = fb_reg_redirect ? _GEN_454 : btb_bj_type_63; // @[BTB.scala 189:28:@2072.6]
  assign _T_2141 = feedback_h_count != 2'h0; // @[BTB.scala 62:38:@2082.12]
  assign _T_2142 = feedback_h_count[1]; // @[BTB.scala 62:45:@2083.12]
  assign _T_2143 = feedback_h_count[0]; // @[BTB.scala 62:54:@2084.12]
  assign _T_2145 = _T_2143 == 1'h0; // @[BTB.scala 62:52:@2085.12]
  assign _T_2146 = _T_2142 | _T_2145; // @[BTB.scala 62:49:@2086.12]
  assign _T_2147 = {_T_2141,_T_2146}; // @[Cat.scala 30:58:@2087.12]
  assign _GEN_647 = 6'h0 == feedback_idx ? _T_2147 : btb_h_count_0; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_648 = 6'h1 == feedback_idx ? _T_2147 : btb_h_count_1; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_649 = 6'h2 == feedback_idx ? _T_2147 : btb_h_count_2; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_650 = 6'h3 == feedback_idx ? _T_2147 : btb_h_count_3; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_651 = 6'h4 == feedback_idx ? _T_2147 : btb_h_count_4; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_652 = 6'h5 == feedback_idx ? _T_2147 : btb_h_count_5; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_653 = 6'h6 == feedback_idx ? _T_2147 : btb_h_count_6; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_654 = 6'h7 == feedback_idx ? _T_2147 : btb_h_count_7; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_655 = 6'h8 == feedback_idx ? _T_2147 : btb_h_count_8; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_656 = 6'h9 == feedback_idx ? _T_2147 : btb_h_count_9; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_657 = 6'ha == feedback_idx ? _T_2147 : btb_h_count_10; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_658 = 6'hb == feedback_idx ? _T_2147 : btb_h_count_11; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_659 = 6'hc == feedback_idx ? _T_2147 : btb_h_count_12; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_660 = 6'hd == feedback_idx ? _T_2147 : btb_h_count_13; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_661 = 6'he == feedback_idx ? _T_2147 : btb_h_count_14; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_662 = 6'hf == feedback_idx ? _T_2147 : btb_h_count_15; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_663 = 6'h10 == feedback_idx ? _T_2147 : btb_h_count_16; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_664 = 6'h11 == feedback_idx ? _T_2147 : btb_h_count_17; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_665 = 6'h12 == feedback_idx ? _T_2147 : btb_h_count_18; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_666 = 6'h13 == feedback_idx ? _T_2147 : btb_h_count_19; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_667 = 6'h14 == feedback_idx ? _T_2147 : btb_h_count_20; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_668 = 6'h15 == feedback_idx ? _T_2147 : btb_h_count_21; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_669 = 6'h16 == feedback_idx ? _T_2147 : btb_h_count_22; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_670 = 6'h17 == feedback_idx ? _T_2147 : btb_h_count_23; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_671 = 6'h18 == feedback_idx ? _T_2147 : btb_h_count_24; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_672 = 6'h19 == feedback_idx ? _T_2147 : btb_h_count_25; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_673 = 6'h1a == feedback_idx ? _T_2147 : btb_h_count_26; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_674 = 6'h1b == feedback_idx ? _T_2147 : btb_h_count_27; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_675 = 6'h1c == feedback_idx ? _T_2147 : btb_h_count_28; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_676 = 6'h1d == feedback_idx ? _T_2147 : btb_h_count_29; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_677 = 6'h1e == feedback_idx ? _T_2147 : btb_h_count_30; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_678 = 6'h1f == feedback_idx ? _T_2147 : btb_h_count_31; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_679 = 6'h20 == feedback_idx ? _T_2147 : btb_h_count_32; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_680 = 6'h21 == feedback_idx ? _T_2147 : btb_h_count_33; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_681 = 6'h22 == feedback_idx ? _T_2147 : btb_h_count_34; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_682 = 6'h23 == feedback_idx ? _T_2147 : btb_h_count_35; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_683 = 6'h24 == feedback_idx ? _T_2147 : btb_h_count_36; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_684 = 6'h25 == feedback_idx ? _T_2147 : btb_h_count_37; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_685 = 6'h26 == feedback_idx ? _T_2147 : btb_h_count_38; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_686 = 6'h27 == feedback_idx ? _T_2147 : btb_h_count_39; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_687 = 6'h28 == feedback_idx ? _T_2147 : btb_h_count_40; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_688 = 6'h29 == feedback_idx ? _T_2147 : btb_h_count_41; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_689 = 6'h2a == feedback_idx ? _T_2147 : btb_h_count_42; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_690 = 6'h2b == feedback_idx ? _T_2147 : btb_h_count_43; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_691 = 6'h2c == feedback_idx ? _T_2147 : btb_h_count_44; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_692 = 6'h2d == feedback_idx ? _T_2147 : btb_h_count_45; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_693 = 6'h2e == feedback_idx ? _T_2147 : btb_h_count_46; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_694 = 6'h2f == feedback_idx ? _T_2147 : btb_h_count_47; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_695 = 6'h30 == feedback_idx ? _T_2147 : btb_h_count_48; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_696 = 6'h31 == feedback_idx ? _T_2147 : btb_h_count_49; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_697 = 6'h32 == feedback_idx ? _T_2147 : btb_h_count_50; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_698 = 6'h33 == feedback_idx ? _T_2147 : btb_h_count_51; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_699 = 6'h34 == feedback_idx ? _T_2147 : btb_h_count_52; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_700 = 6'h35 == feedback_idx ? _T_2147 : btb_h_count_53; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_701 = 6'h36 == feedback_idx ? _T_2147 : btb_h_count_54; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_702 = 6'h37 == feedback_idx ? _T_2147 : btb_h_count_55; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_703 = 6'h38 == feedback_idx ? _T_2147 : btb_h_count_56; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_704 = 6'h39 == feedback_idx ? _T_2147 : btb_h_count_57; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_705 = 6'h3a == feedback_idx ? _T_2147 : btb_h_count_58; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_706 = 6'h3b == feedback_idx ? _T_2147 : btb_h_count_59; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_707 = 6'h3c == feedback_idx ? _T_2147 : btb_h_count_60; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_708 = 6'h3d == feedback_idx ? _T_2147 : btb_h_count_61; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_709 = 6'h3e == feedback_idx ? _T_2147 : btb_h_count_62; // @[BTB.scala 198:37:@2088.12]
  assign _GEN_710 = 6'h3f == feedback_idx ? _T_2147 : btb_h_count_63; // @[BTB.scala 198:37:@2088.12]
  assign feedback_gshare = bht__T_1774_data; // @[BTB.scala 170:22:@1322.4 BTB.scala 179:20:@1775.4]
  assign _T_2150 = feedback_gshare != 2'h0; // @[BTB.scala 62:38:@2090.12]
  assign _T_2151 = feedback_gshare[1]; // @[BTB.scala 62:45:@2091.12]
  assign _T_2152 = feedback_gshare[0]; // @[BTB.scala 62:54:@2092.12]
  assign _T_2154 = _T_2152 == 1'h0; // @[BTB.scala 62:52:@2093.12]
  assign _T_2155 = _T_2151 | _T_2154; // @[BTB.scala 62:49:@2094.12]
  assign _T_2157 = ~ feedback_h_count; // @[BTB.scala 64:38:@2099.12]
  assign _T_2159 = _T_2157 == 2'h0; // @[BTB.scala 64:38:@2100.12]
  assign _T_2164 = _T_2142 & _T_2145; // @[BTB.scala 64:49:@2104.12]
  assign _T_2165 = {_T_2159,_T_2164}; // @[Cat.scala 30:58:@2105.12]
  assign _GEN_711 = 6'h0 == feedback_idx ? _T_2165 : btb_h_count_0; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_712 = 6'h1 == feedback_idx ? _T_2165 : btb_h_count_1; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_713 = 6'h2 == feedback_idx ? _T_2165 : btb_h_count_2; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_714 = 6'h3 == feedback_idx ? _T_2165 : btb_h_count_3; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_715 = 6'h4 == feedback_idx ? _T_2165 : btb_h_count_4; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_716 = 6'h5 == feedback_idx ? _T_2165 : btb_h_count_5; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_717 = 6'h6 == feedback_idx ? _T_2165 : btb_h_count_6; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_718 = 6'h7 == feedback_idx ? _T_2165 : btb_h_count_7; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_719 = 6'h8 == feedback_idx ? _T_2165 : btb_h_count_8; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_720 = 6'h9 == feedback_idx ? _T_2165 : btb_h_count_9; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_721 = 6'ha == feedback_idx ? _T_2165 : btb_h_count_10; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_722 = 6'hb == feedback_idx ? _T_2165 : btb_h_count_11; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_723 = 6'hc == feedback_idx ? _T_2165 : btb_h_count_12; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_724 = 6'hd == feedback_idx ? _T_2165 : btb_h_count_13; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_725 = 6'he == feedback_idx ? _T_2165 : btb_h_count_14; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_726 = 6'hf == feedback_idx ? _T_2165 : btb_h_count_15; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_727 = 6'h10 == feedback_idx ? _T_2165 : btb_h_count_16; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_728 = 6'h11 == feedback_idx ? _T_2165 : btb_h_count_17; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_729 = 6'h12 == feedback_idx ? _T_2165 : btb_h_count_18; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_730 = 6'h13 == feedback_idx ? _T_2165 : btb_h_count_19; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_731 = 6'h14 == feedback_idx ? _T_2165 : btb_h_count_20; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_732 = 6'h15 == feedback_idx ? _T_2165 : btb_h_count_21; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_733 = 6'h16 == feedback_idx ? _T_2165 : btb_h_count_22; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_734 = 6'h17 == feedback_idx ? _T_2165 : btb_h_count_23; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_735 = 6'h18 == feedback_idx ? _T_2165 : btb_h_count_24; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_736 = 6'h19 == feedback_idx ? _T_2165 : btb_h_count_25; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_737 = 6'h1a == feedback_idx ? _T_2165 : btb_h_count_26; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_738 = 6'h1b == feedback_idx ? _T_2165 : btb_h_count_27; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_739 = 6'h1c == feedback_idx ? _T_2165 : btb_h_count_28; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_740 = 6'h1d == feedback_idx ? _T_2165 : btb_h_count_29; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_741 = 6'h1e == feedback_idx ? _T_2165 : btb_h_count_30; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_742 = 6'h1f == feedback_idx ? _T_2165 : btb_h_count_31; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_743 = 6'h20 == feedback_idx ? _T_2165 : btb_h_count_32; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_744 = 6'h21 == feedback_idx ? _T_2165 : btb_h_count_33; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_745 = 6'h22 == feedback_idx ? _T_2165 : btb_h_count_34; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_746 = 6'h23 == feedback_idx ? _T_2165 : btb_h_count_35; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_747 = 6'h24 == feedback_idx ? _T_2165 : btb_h_count_36; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_748 = 6'h25 == feedback_idx ? _T_2165 : btb_h_count_37; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_749 = 6'h26 == feedback_idx ? _T_2165 : btb_h_count_38; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_750 = 6'h27 == feedback_idx ? _T_2165 : btb_h_count_39; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_751 = 6'h28 == feedback_idx ? _T_2165 : btb_h_count_40; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_752 = 6'h29 == feedback_idx ? _T_2165 : btb_h_count_41; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_753 = 6'h2a == feedback_idx ? _T_2165 : btb_h_count_42; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_754 = 6'h2b == feedback_idx ? _T_2165 : btb_h_count_43; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_755 = 6'h2c == feedback_idx ? _T_2165 : btb_h_count_44; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_756 = 6'h2d == feedback_idx ? _T_2165 : btb_h_count_45; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_757 = 6'h2e == feedback_idx ? _T_2165 : btb_h_count_46; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_758 = 6'h2f == feedback_idx ? _T_2165 : btb_h_count_47; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_759 = 6'h30 == feedback_idx ? _T_2165 : btb_h_count_48; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_760 = 6'h31 == feedback_idx ? _T_2165 : btb_h_count_49; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_761 = 6'h32 == feedback_idx ? _T_2165 : btb_h_count_50; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_762 = 6'h33 == feedback_idx ? _T_2165 : btb_h_count_51; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_763 = 6'h34 == feedback_idx ? _T_2165 : btb_h_count_52; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_764 = 6'h35 == feedback_idx ? _T_2165 : btb_h_count_53; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_765 = 6'h36 == feedback_idx ? _T_2165 : btb_h_count_54; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_766 = 6'h37 == feedback_idx ? _T_2165 : btb_h_count_55; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_767 = 6'h38 == feedback_idx ? _T_2165 : btb_h_count_56; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_768 = 6'h39 == feedback_idx ? _T_2165 : btb_h_count_57; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_769 = 6'h3a == feedback_idx ? _T_2165 : btb_h_count_58; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_770 = 6'h3b == feedback_idx ? _T_2165 : btb_h_count_59; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_771 = 6'h3c == feedback_idx ? _T_2165 : btb_h_count_60; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_772 = 6'h3d == feedback_idx ? _T_2165 : btb_h_count_61; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_773 = 6'h3e == feedback_idx ? _T_2165 : btb_h_count_62; // @[BTB.scala 201:37:@2106.12]
  assign _GEN_774 = 6'h3f == feedback_idx ? _T_2165 : btb_h_count_63; // @[BTB.scala 201:37:@2106.12]
  assign _T_2167 = ~ feedback_gshare; // @[BTB.scala 64:38:@2108.12]
  assign _T_2169 = _T_2167 == 2'h0; // @[BTB.scala 64:38:@2109.12]
  assign _T_2174 = _T_2151 & _T_2154; // @[BTB.scala 64:49:@2113.12]
  assign _GEN_775 = fb_reg_redirect ? _GEN_647 : _GEN_711; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_776 = fb_reg_redirect ? _GEN_648 : _GEN_712; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_777 = fb_reg_redirect ? _GEN_649 : _GEN_713; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_778 = fb_reg_redirect ? _GEN_650 : _GEN_714; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_779 = fb_reg_redirect ? _GEN_651 : _GEN_715; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_780 = fb_reg_redirect ? _GEN_652 : _GEN_716; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_781 = fb_reg_redirect ? _GEN_653 : _GEN_717; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_782 = fb_reg_redirect ? _GEN_654 : _GEN_718; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_783 = fb_reg_redirect ? _GEN_655 : _GEN_719; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_784 = fb_reg_redirect ? _GEN_656 : _GEN_720; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_785 = fb_reg_redirect ? _GEN_657 : _GEN_721; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_786 = fb_reg_redirect ? _GEN_658 : _GEN_722; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_787 = fb_reg_redirect ? _GEN_659 : _GEN_723; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_788 = fb_reg_redirect ? _GEN_660 : _GEN_724; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_789 = fb_reg_redirect ? _GEN_661 : _GEN_725; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_790 = fb_reg_redirect ? _GEN_662 : _GEN_726; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_791 = fb_reg_redirect ? _GEN_663 : _GEN_727; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_792 = fb_reg_redirect ? _GEN_664 : _GEN_728; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_793 = fb_reg_redirect ? _GEN_665 : _GEN_729; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_794 = fb_reg_redirect ? _GEN_666 : _GEN_730; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_795 = fb_reg_redirect ? _GEN_667 : _GEN_731; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_796 = fb_reg_redirect ? _GEN_668 : _GEN_732; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_797 = fb_reg_redirect ? _GEN_669 : _GEN_733; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_798 = fb_reg_redirect ? _GEN_670 : _GEN_734; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_799 = fb_reg_redirect ? _GEN_671 : _GEN_735; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_800 = fb_reg_redirect ? _GEN_672 : _GEN_736; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_801 = fb_reg_redirect ? _GEN_673 : _GEN_737; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_802 = fb_reg_redirect ? _GEN_674 : _GEN_738; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_803 = fb_reg_redirect ? _GEN_675 : _GEN_739; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_804 = fb_reg_redirect ? _GEN_676 : _GEN_740; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_805 = fb_reg_redirect ? _GEN_677 : _GEN_741; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_806 = fb_reg_redirect ? _GEN_678 : _GEN_742; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_807 = fb_reg_redirect ? _GEN_679 : _GEN_743; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_808 = fb_reg_redirect ? _GEN_680 : _GEN_744; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_809 = fb_reg_redirect ? _GEN_681 : _GEN_745; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_810 = fb_reg_redirect ? _GEN_682 : _GEN_746; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_811 = fb_reg_redirect ? _GEN_683 : _GEN_747; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_812 = fb_reg_redirect ? _GEN_684 : _GEN_748; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_813 = fb_reg_redirect ? _GEN_685 : _GEN_749; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_814 = fb_reg_redirect ? _GEN_686 : _GEN_750; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_815 = fb_reg_redirect ? _GEN_687 : _GEN_751; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_816 = fb_reg_redirect ? _GEN_688 : _GEN_752; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_817 = fb_reg_redirect ? _GEN_689 : _GEN_753; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_818 = fb_reg_redirect ? _GEN_690 : _GEN_754; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_819 = fb_reg_redirect ? _GEN_691 : _GEN_755; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_820 = fb_reg_redirect ? _GEN_692 : _GEN_756; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_821 = fb_reg_redirect ? _GEN_693 : _GEN_757; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_822 = fb_reg_redirect ? _GEN_694 : _GEN_758; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_823 = fb_reg_redirect ? _GEN_695 : _GEN_759; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_824 = fb_reg_redirect ? _GEN_696 : _GEN_760; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_825 = fb_reg_redirect ? _GEN_697 : _GEN_761; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_826 = fb_reg_redirect ? _GEN_698 : _GEN_762; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_827 = fb_reg_redirect ? _GEN_699 : _GEN_763; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_828 = fb_reg_redirect ? _GEN_700 : _GEN_764; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_829 = fb_reg_redirect ? _GEN_701 : _GEN_765; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_830 = fb_reg_redirect ? _GEN_702 : _GEN_766; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_831 = fb_reg_redirect ? _GEN_703 : _GEN_767; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_832 = fb_reg_redirect ? _GEN_704 : _GEN_768; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_833 = fb_reg_redirect ? _GEN_705 : _GEN_769; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_834 = fb_reg_redirect ? _GEN_706 : _GEN_770; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_835 = fb_reg_redirect ? _GEN_707 : _GEN_771; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_836 = fb_reg_redirect ? _GEN_708 : _GEN_772; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_837 = fb_reg_redirect ? _GEN_709 : _GEN_773; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_838 = fb_reg_redirect ? _GEN_710 : _GEN_774; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_846 = fb_reg_redirect ? 1'h0 : 1'h1; // @[BTB.scala 197:32:@2081.10]
  assign _GEN_849 = 6'h0 == feedback_idx ? 2'h2 : btb_h_count_0; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_850 = 6'h1 == feedback_idx ? 2'h2 : btb_h_count_1; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_851 = 6'h2 == feedback_idx ? 2'h2 : btb_h_count_2; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_852 = 6'h3 == feedback_idx ? 2'h2 : btb_h_count_3; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_853 = 6'h4 == feedback_idx ? 2'h2 : btb_h_count_4; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_854 = 6'h5 == feedback_idx ? 2'h2 : btb_h_count_5; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_855 = 6'h6 == feedback_idx ? 2'h2 : btb_h_count_6; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_856 = 6'h7 == feedback_idx ? 2'h2 : btb_h_count_7; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_857 = 6'h8 == feedback_idx ? 2'h2 : btb_h_count_8; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_858 = 6'h9 == feedback_idx ? 2'h2 : btb_h_count_9; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_859 = 6'ha == feedback_idx ? 2'h2 : btb_h_count_10; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_860 = 6'hb == feedback_idx ? 2'h2 : btb_h_count_11; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_861 = 6'hc == feedback_idx ? 2'h2 : btb_h_count_12; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_862 = 6'hd == feedback_idx ? 2'h2 : btb_h_count_13; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_863 = 6'he == feedback_idx ? 2'h2 : btb_h_count_14; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_864 = 6'hf == feedback_idx ? 2'h2 : btb_h_count_15; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_865 = 6'h10 == feedback_idx ? 2'h2 : btb_h_count_16; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_866 = 6'h11 == feedback_idx ? 2'h2 : btb_h_count_17; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_867 = 6'h12 == feedback_idx ? 2'h2 : btb_h_count_18; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_868 = 6'h13 == feedback_idx ? 2'h2 : btb_h_count_19; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_869 = 6'h14 == feedback_idx ? 2'h2 : btb_h_count_20; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_870 = 6'h15 == feedback_idx ? 2'h2 : btb_h_count_21; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_871 = 6'h16 == feedback_idx ? 2'h2 : btb_h_count_22; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_872 = 6'h17 == feedback_idx ? 2'h2 : btb_h_count_23; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_873 = 6'h18 == feedback_idx ? 2'h2 : btb_h_count_24; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_874 = 6'h19 == feedback_idx ? 2'h2 : btb_h_count_25; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_875 = 6'h1a == feedback_idx ? 2'h2 : btb_h_count_26; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_876 = 6'h1b == feedback_idx ? 2'h2 : btb_h_count_27; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_877 = 6'h1c == feedback_idx ? 2'h2 : btb_h_count_28; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_878 = 6'h1d == feedback_idx ? 2'h2 : btb_h_count_29; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_879 = 6'h1e == feedback_idx ? 2'h2 : btb_h_count_30; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_880 = 6'h1f == feedback_idx ? 2'h2 : btb_h_count_31; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_881 = 6'h20 == feedback_idx ? 2'h2 : btb_h_count_32; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_882 = 6'h21 == feedback_idx ? 2'h2 : btb_h_count_33; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_883 = 6'h22 == feedback_idx ? 2'h2 : btb_h_count_34; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_884 = 6'h23 == feedback_idx ? 2'h2 : btb_h_count_35; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_885 = 6'h24 == feedback_idx ? 2'h2 : btb_h_count_36; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_886 = 6'h25 == feedback_idx ? 2'h2 : btb_h_count_37; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_887 = 6'h26 == feedback_idx ? 2'h2 : btb_h_count_38; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_888 = 6'h27 == feedback_idx ? 2'h2 : btb_h_count_39; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_889 = 6'h28 == feedback_idx ? 2'h2 : btb_h_count_40; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_890 = 6'h29 == feedback_idx ? 2'h2 : btb_h_count_41; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_891 = 6'h2a == feedback_idx ? 2'h2 : btb_h_count_42; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_892 = 6'h2b == feedback_idx ? 2'h2 : btb_h_count_43; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_893 = 6'h2c == feedback_idx ? 2'h2 : btb_h_count_44; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_894 = 6'h2d == feedback_idx ? 2'h2 : btb_h_count_45; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_895 = 6'h2e == feedback_idx ? 2'h2 : btb_h_count_46; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_896 = 6'h2f == feedback_idx ? 2'h2 : btb_h_count_47; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_897 = 6'h30 == feedback_idx ? 2'h2 : btb_h_count_48; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_898 = 6'h31 == feedback_idx ? 2'h2 : btb_h_count_49; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_899 = 6'h32 == feedback_idx ? 2'h2 : btb_h_count_50; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_900 = 6'h33 == feedback_idx ? 2'h2 : btb_h_count_51; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_901 = 6'h34 == feedback_idx ? 2'h2 : btb_h_count_52; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_902 = 6'h35 == feedback_idx ? 2'h2 : btb_h_count_53; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_903 = 6'h36 == feedback_idx ? 2'h2 : btb_h_count_54; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_904 = 6'h37 == feedback_idx ? 2'h2 : btb_h_count_55; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_905 = 6'h38 == feedback_idx ? 2'h2 : btb_h_count_56; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_906 = 6'h39 == feedback_idx ? 2'h2 : btb_h_count_57; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_907 = 6'h3a == feedback_idx ? 2'h2 : btb_h_count_58; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_908 = 6'h3b == feedback_idx ? 2'h2 : btb_h_count_59; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_909 = 6'h3c == feedback_idx ? 2'h2 : btb_h_count_60; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_910 = 6'h3d == feedback_idx ? 2'h2 : btb_h_count_61; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_911 = 6'h3e == feedback_idx ? 2'h2 : btb_h_count_62; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_912 = 6'h3f == feedback_idx ? 2'h2 : btb_h_count_63; // @[BTB.scala 205:35:@2120.12]
  assign _GEN_913 = fb_reg_redirect ? _GEN_849 : btb_h_count_0; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_914 = fb_reg_redirect ? _GEN_850 : btb_h_count_1; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_915 = fb_reg_redirect ? _GEN_851 : btb_h_count_2; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_916 = fb_reg_redirect ? _GEN_852 : btb_h_count_3; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_917 = fb_reg_redirect ? _GEN_853 : btb_h_count_4; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_918 = fb_reg_redirect ? _GEN_854 : btb_h_count_5; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_919 = fb_reg_redirect ? _GEN_855 : btb_h_count_6; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_920 = fb_reg_redirect ? _GEN_856 : btb_h_count_7; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_921 = fb_reg_redirect ? _GEN_857 : btb_h_count_8; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_922 = fb_reg_redirect ? _GEN_858 : btb_h_count_9; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_923 = fb_reg_redirect ? _GEN_859 : btb_h_count_10; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_924 = fb_reg_redirect ? _GEN_860 : btb_h_count_11; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_925 = fb_reg_redirect ? _GEN_861 : btb_h_count_12; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_926 = fb_reg_redirect ? _GEN_862 : btb_h_count_13; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_927 = fb_reg_redirect ? _GEN_863 : btb_h_count_14; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_928 = fb_reg_redirect ? _GEN_864 : btb_h_count_15; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_929 = fb_reg_redirect ? _GEN_865 : btb_h_count_16; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_930 = fb_reg_redirect ? _GEN_866 : btb_h_count_17; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_931 = fb_reg_redirect ? _GEN_867 : btb_h_count_18; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_932 = fb_reg_redirect ? _GEN_868 : btb_h_count_19; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_933 = fb_reg_redirect ? _GEN_869 : btb_h_count_20; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_934 = fb_reg_redirect ? _GEN_870 : btb_h_count_21; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_935 = fb_reg_redirect ? _GEN_871 : btb_h_count_22; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_936 = fb_reg_redirect ? _GEN_872 : btb_h_count_23; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_937 = fb_reg_redirect ? _GEN_873 : btb_h_count_24; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_938 = fb_reg_redirect ? _GEN_874 : btb_h_count_25; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_939 = fb_reg_redirect ? _GEN_875 : btb_h_count_26; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_940 = fb_reg_redirect ? _GEN_876 : btb_h_count_27; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_941 = fb_reg_redirect ? _GEN_877 : btb_h_count_28; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_942 = fb_reg_redirect ? _GEN_878 : btb_h_count_29; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_943 = fb_reg_redirect ? _GEN_879 : btb_h_count_30; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_944 = fb_reg_redirect ? _GEN_880 : btb_h_count_31; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_945 = fb_reg_redirect ? _GEN_881 : btb_h_count_32; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_946 = fb_reg_redirect ? _GEN_882 : btb_h_count_33; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_947 = fb_reg_redirect ? _GEN_883 : btb_h_count_34; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_948 = fb_reg_redirect ? _GEN_884 : btb_h_count_35; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_949 = fb_reg_redirect ? _GEN_885 : btb_h_count_36; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_950 = fb_reg_redirect ? _GEN_886 : btb_h_count_37; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_951 = fb_reg_redirect ? _GEN_887 : btb_h_count_38; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_952 = fb_reg_redirect ? _GEN_888 : btb_h_count_39; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_953 = fb_reg_redirect ? _GEN_889 : btb_h_count_40; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_954 = fb_reg_redirect ? _GEN_890 : btb_h_count_41; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_955 = fb_reg_redirect ? _GEN_891 : btb_h_count_42; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_956 = fb_reg_redirect ? _GEN_892 : btb_h_count_43; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_957 = fb_reg_redirect ? _GEN_893 : btb_h_count_44; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_958 = fb_reg_redirect ? _GEN_894 : btb_h_count_45; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_959 = fb_reg_redirect ? _GEN_895 : btb_h_count_46; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_960 = fb_reg_redirect ? _GEN_896 : btb_h_count_47; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_961 = fb_reg_redirect ? _GEN_897 : btb_h_count_48; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_962 = fb_reg_redirect ? _GEN_898 : btb_h_count_49; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_963 = fb_reg_redirect ? _GEN_899 : btb_h_count_50; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_964 = fb_reg_redirect ? _GEN_900 : btb_h_count_51; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_965 = fb_reg_redirect ? _GEN_901 : btb_h_count_52; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_966 = fb_reg_redirect ? _GEN_902 : btb_h_count_53; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_967 = fb_reg_redirect ? _GEN_903 : btb_h_count_54; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_968 = fb_reg_redirect ? _GEN_904 : btb_h_count_55; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_969 = fb_reg_redirect ? _GEN_905 : btb_h_count_56; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_970 = fb_reg_redirect ? _GEN_906 : btb_h_count_57; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_971 = fb_reg_redirect ? _GEN_907 : btb_h_count_58; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_972 = fb_reg_redirect ? _GEN_908 : btb_h_count_59; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_973 = fb_reg_redirect ? _GEN_909 : btb_h_count_60; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_974 = fb_reg_redirect ? _GEN_910 : btb_h_count_61; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_975 = fb_reg_redirect ? _GEN_911 : btb_h_count_62; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_976 = fb_reg_redirect ? _GEN_912 : btb_h_count_63; // @[BTB.scala 204:35:@2119.10]
  assign _GEN_978 = _T_1776 ? _GEN_775 : _GEN_913; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_979 = _T_1776 ? _GEN_776 : _GEN_914; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_980 = _T_1776 ? _GEN_777 : _GEN_915; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_981 = _T_1776 ? _GEN_778 : _GEN_916; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_982 = _T_1776 ? _GEN_779 : _GEN_917; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_983 = _T_1776 ? _GEN_780 : _GEN_918; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_984 = _T_1776 ? _GEN_781 : _GEN_919; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_985 = _T_1776 ? _GEN_782 : _GEN_920; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_986 = _T_1776 ? _GEN_783 : _GEN_921; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_987 = _T_1776 ? _GEN_784 : _GEN_922; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_988 = _T_1776 ? _GEN_785 : _GEN_923; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_989 = _T_1776 ? _GEN_786 : _GEN_924; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_990 = _T_1776 ? _GEN_787 : _GEN_925; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_991 = _T_1776 ? _GEN_788 : _GEN_926; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_992 = _T_1776 ? _GEN_789 : _GEN_927; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_993 = _T_1776 ? _GEN_790 : _GEN_928; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_994 = _T_1776 ? _GEN_791 : _GEN_929; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_995 = _T_1776 ? _GEN_792 : _GEN_930; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_996 = _T_1776 ? _GEN_793 : _GEN_931; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_997 = _T_1776 ? _GEN_794 : _GEN_932; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_998 = _T_1776 ? _GEN_795 : _GEN_933; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_999 = _T_1776 ? _GEN_796 : _GEN_934; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1000 = _T_1776 ? _GEN_797 : _GEN_935; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1001 = _T_1776 ? _GEN_798 : _GEN_936; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1002 = _T_1776 ? _GEN_799 : _GEN_937; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1003 = _T_1776 ? _GEN_800 : _GEN_938; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1004 = _T_1776 ? _GEN_801 : _GEN_939; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1005 = _T_1776 ? _GEN_802 : _GEN_940; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1006 = _T_1776 ? _GEN_803 : _GEN_941; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1007 = _T_1776 ? _GEN_804 : _GEN_942; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1008 = _T_1776 ? _GEN_805 : _GEN_943; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1009 = _T_1776 ? _GEN_806 : _GEN_944; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1010 = _T_1776 ? _GEN_807 : _GEN_945; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1011 = _T_1776 ? _GEN_808 : _GEN_946; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1012 = _T_1776 ? _GEN_809 : _GEN_947; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1013 = _T_1776 ? _GEN_810 : _GEN_948; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1014 = _T_1776 ? _GEN_811 : _GEN_949; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1015 = _T_1776 ? _GEN_812 : _GEN_950; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1016 = _T_1776 ? _GEN_813 : _GEN_951; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1017 = _T_1776 ? _GEN_814 : _GEN_952; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1018 = _T_1776 ? _GEN_815 : _GEN_953; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1019 = _T_1776 ? _GEN_816 : _GEN_954; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1020 = _T_1776 ? _GEN_817 : _GEN_955; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1021 = _T_1776 ? _GEN_818 : _GEN_956; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1022 = _T_1776 ? _GEN_819 : _GEN_957; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1023 = _T_1776 ? _GEN_820 : _GEN_958; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1024 = _T_1776 ? _GEN_821 : _GEN_959; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1025 = _T_1776 ? _GEN_822 : _GEN_960; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1026 = _T_1776 ? _GEN_823 : _GEN_961; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1027 = _T_1776 ? _GEN_824 : _GEN_962; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1028 = _T_1776 ? _GEN_825 : _GEN_963; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1029 = _T_1776 ? _GEN_826 : _GEN_964; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1030 = _T_1776 ? _GEN_827 : _GEN_965; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1031 = _T_1776 ? _GEN_828 : _GEN_966; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1032 = _T_1776 ? _GEN_829 : _GEN_967; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1033 = _T_1776 ? _GEN_830 : _GEN_968; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1034 = _T_1776 ? _GEN_831 : _GEN_969; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1035 = _T_1776 ? _GEN_832 : _GEN_970; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1036 = _T_1776 ? _GEN_833 : _GEN_971; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1037 = _T_1776 ? _GEN_834 : _GEN_972; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1038 = _T_1776 ? _GEN_835 : _GEN_973; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1039 = _T_1776 ? _GEN_836 : _GEN_974; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1040 = _T_1776 ? _GEN_837 : _GEN_975; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1041 = _T_1776 ? _GEN_838 : _GEN_976; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1044 = _T_1776 ? fb_reg_redirect : 1'h0; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1049 = _T_1776 ? _GEN_846 : 1'h0; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1054 = _T_1776 ? 1'h0 : fb_reg_redirect; // @[BTB.scala 196:29:@2080.8]
  assign _GEN_1057 = _T_2135 ? _GEN_978 : btb_h_count_0; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1058 = _T_2135 ? _GEN_979 : btb_h_count_1; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1059 = _T_2135 ? _GEN_980 : btb_h_count_2; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1060 = _T_2135 ? _GEN_981 : btb_h_count_3; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1061 = _T_2135 ? _GEN_982 : btb_h_count_4; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1062 = _T_2135 ? _GEN_983 : btb_h_count_5; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1063 = _T_2135 ? _GEN_984 : btb_h_count_6; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1064 = _T_2135 ? _GEN_985 : btb_h_count_7; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1065 = _T_2135 ? _GEN_986 : btb_h_count_8; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1066 = _T_2135 ? _GEN_987 : btb_h_count_9; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1067 = _T_2135 ? _GEN_988 : btb_h_count_10; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1068 = _T_2135 ? _GEN_989 : btb_h_count_11; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1069 = _T_2135 ? _GEN_990 : btb_h_count_12; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1070 = _T_2135 ? _GEN_991 : btb_h_count_13; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1071 = _T_2135 ? _GEN_992 : btb_h_count_14; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1072 = _T_2135 ? _GEN_993 : btb_h_count_15; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1073 = _T_2135 ? _GEN_994 : btb_h_count_16; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1074 = _T_2135 ? _GEN_995 : btb_h_count_17; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1075 = _T_2135 ? _GEN_996 : btb_h_count_18; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1076 = _T_2135 ? _GEN_997 : btb_h_count_19; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1077 = _T_2135 ? _GEN_998 : btb_h_count_20; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1078 = _T_2135 ? _GEN_999 : btb_h_count_21; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1079 = _T_2135 ? _GEN_1000 : btb_h_count_22; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1080 = _T_2135 ? _GEN_1001 : btb_h_count_23; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1081 = _T_2135 ? _GEN_1002 : btb_h_count_24; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1082 = _T_2135 ? _GEN_1003 : btb_h_count_25; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1083 = _T_2135 ? _GEN_1004 : btb_h_count_26; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1084 = _T_2135 ? _GEN_1005 : btb_h_count_27; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1085 = _T_2135 ? _GEN_1006 : btb_h_count_28; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1086 = _T_2135 ? _GEN_1007 : btb_h_count_29; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1087 = _T_2135 ? _GEN_1008 : btb_h_count_30; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1088 = _T_2135 ? _GEN_1009 : btb_h_count_31; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1089 = _T_2135 ? _GEN_1010 : btb_h_count_32; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1090 = _T_2135 ? _GEN_1011 : btb_h_count_33; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1091 = _T_2135 ? _GEN_1012 : btb_h_count_34; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1092 = _T_2135 ? _GEN_1013 : btb_h_count_35; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1093 = _T_2135 ? _GEN_1014 : btb_h_count_36; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1094 = _T_2135 ? _GEN_1015 : btb_h_count_37; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1095 = _T_2135 ? _GEN_1016 : btb_h_count_38; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1096 = _T_2135 ? _GEN_1017 : btb_h_count_39; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1097 = _T_2135 ? _GEN_1018 : btb_h_count_40; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1098 = _T_2135 ? _GEN_1019 : btb_h_count_41; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1099 = _T_2135 ? _GEN_1020 : btb_h_count_42; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1100 = _T_2135 ? _GEN_1021 : btb_h_count_43; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1101 = _T_2135 ? _GEN_1022 : btb_h_count_44; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1102 = _T_2135 ? _GEN_1023 : btb_h_count_45; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1103 = _T_2135 ? _GEN_1024 : btb_h_count_46; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1104 = _T_2135 ? _GEN_1025 : btb_h_count_47; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1105 = _T_2135 ? _GEN_1026 : btb_h_count_48; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1106 = _T_2135 ? _GEN_1027 : btb_h_count_49; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1107 = _T_2135 ? _GEN_1028 : btb_h_count_50; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1108 = _T_2135 ? _GEN_1029 : btb_h_count_51; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1109 = _T_2135 ? _GEN_1030 : btb_h_count_52; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1110 = _T_2135 ? _GEN_1031 : btb_h_count_53; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1111 = _T_2135 ? _GEN_1032 : btb_h_count_54; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1112 = _T_2135 ? _GEN_1033 : btb_h_count_55; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1113 = _T_2135 ? _GEN_1034 : btb_h_count_56; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1114 = _T_2135 ? _GEN_1035 : btb_h_count_57; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1115 = _T_2135 ? _GEN_1036 : btb_h_count_58; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1116 = _T_2135 ? _GEN_1037 : btb_h_count_59; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1117 = _T_2135 ? _GEN_1038 : btb_h_count_60; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1118 = _T_2135 ? _GEN_1039 : btb_h_count_61; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1119 = _T_2135 ? _GEN_1040 : btb_h_count_62; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1120 = _T_2135 ? _GEN_1041 : btb_h_count_63; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1123 = _T_2135 ? _GEN_1044 : 1'h0; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1128 = _T_2135 ? _GEN_1049 : 1'h0; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1133 = _T_2135 ? _GEN_1054 : 1'h0; // @[BTB.scala 195:49:@2078.6]
  assign _GEN_1136 = fb_reg_valid ? _GEN_199 : btb_valid_0; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1137 = fb_reg_valid ? _GEN_200 : btb_valid_1; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1138 = fb_reg_valid ? _GEN_201 : btb_valid_2; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1139 = fb_reg_valid ? _GEN_202 : btb_valid_3; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1140 = fb_reg_valid ? _GEN_203 : btb_valid_4; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1141 = fb_reg_valid ? _GEN_204 : btb_valid_5; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1142 = fb_reg_valid ? _GEN_205 : btb_valid_6; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1143 = fb_reg_valid ? _GEN_206 : btb_valid_7; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1144 = fb_reg_valid ? _GEN_207 : btb_valid_8; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1145 = fb_reg_valid ? _GEN_208 : btb_valid_9; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1146 = fb_reg_valid ? _GEN_209 : btb_valid_10; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1147 = fb_reg_valid ? _GEN_210 : btb_valid_11; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1148 = fb_reg_valid ? _GEN_211 : btb_valid_12; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1149 = fb_reg_valid ? _GEN_212 : btb_valid_13; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1150 = fb_reg_valid ? _GEN_213 : btb_valid_14; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1151 = fb_reg_valid ? _GEN_214 : btb_valid_15; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1152 = fb_reg_valid ? _GEN_215 : btb_valid_16; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1153 = fb_reg_valid ? _GEN_216 : btb_valid_17; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1154 = fb_reg_valid ? _GEN_217 : btb_valid_18; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1155 = fb_reg_valid ? _GEN_218 : btb_valid_19; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1156 = fb_reg_valid ? _GEN_219 : btb_valid_20; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1157 = fb_reg_valid ? _GEN_220 : btb_valid_21; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1158 = fb_reg_valid ? _GEN_221 : btb_valid_22; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1159 = fb_reg_valid ? _GEN_222 : btb_valid_23; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1160 = fb_reg_valid ? _GEN_223 : btb_valid_24; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1161 = fb_reg_valid ? _GEN_224 : btb_valid_25; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1162 = fb_reg_valid ? _GEN_225 : btb_valid_26; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1163 = fb_reg_valid ? _GEN_226 : btb_valid_27; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1164 = fb_reg_valid ? _GEN_227 : btb_valid_28; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1165 = fb_reg_valid ? _GEN_228 : btb_valid_29; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1166 = fb_reg_valid ? _GEN_229 : btb_valid_30; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1167 = fb_reg_valid ? _GEN_230 : btb_valid_31; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1168 = fb_reg_valid ? _GEN_231 : btb_valid_32; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1169 = fb_reg_valid ? _GEN_232 : btb_valid_33; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1170 = fb_reg_valid ? _GEN_233 : btb_valid_34; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1171 = fb_reg_valid ? _GEN_234 : btb_valid_35; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1172 = fb_reg_valid ? _GEN_235 : btb_valid_36; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1173 = fb_reg_valid ? _GEN_236 : btb_valid_37; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1174 = fb_reg_valid ? _GEN_237 : btb_valid_38; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1175 = fb_reg_valid ? _GEN_238 : btb_valid_39; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1176 = fb_reg_valid ? _GEN_239 : btb_valid_40; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1177 = fb_reg_valid ? _GEN_240 : btb_valid_41; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1178 = fb_reg_valid ? _GEN_241 : btb_valid_42; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1179 = fb_reg_valid ? _GEN_242 : btb_valid_43; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1180 = fb_reg_valid ? _GEN_243 : btb_valid_44; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1181 = fb_reg_valid ? _GEN_244 : btb_valid_45; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1182 = fb_reg_valid ? _GEN_245 : btb_valid_46; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1183 = fb_reg_valid ? _GEN_246 : btb_valid_47; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1184 = fb_reg_valid ? _GEN_247 : btb_valid_48; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1185 = fb_reg_valid ? _GEN_248 : btb_valid_49; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1186 = fb_reg_valid ? _GEN_249 : btb_valid_50; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1187 = fb_reg_valid ? _GEN_250 : btb_valid_51; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1188 = fb_reg_valid ? _GEN_251 : btb_valid_52; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1189 = fb_reg_valid ? _GEN_252 : btb_valid_53; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1190 = fb_reg_valid ? _GEN_253 : btb_valid_54; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1191 = fb_reg_valid ? _GEN_254 : btb_valid_55; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1192 = fb_reg_valid ? _GEN_255 : btb_valid_56; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1193 = fb_reg_valid ? _GEN_256 : btb_valid_57; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1194 = fb_reg_valid ? _GEN_257 : btb_valid_58; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1195 = fb_reg_valid ? _GEN_258 : btb_valid_59; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1196 = fb_reg_valid ? _GEN_259 : btb_valid_60; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1197 = fb_reg_valid ? _GEN_260 : btb_valid_61; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1198 = fb_reg_valid ? _GEN_261 : btb_valid_62; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1199 = fb_reg_valid ? _GEN_262 : btb_valid_63; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1200 = fb_reg_valid ? _GEN_455 : btb_pc_0; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1201 = fb_reg_valid ? _GEN_456 : btb_pc_1; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1202 = fb_reg_valid ? _GEN_457 : btb_pc_2; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1203 = fb_reg_valid ? _GEN_458 : btb_pc_3; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1204 = fb_reg_valid ? _GEN_459 : btb_pc_4; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1205 = fb_reg_valid ? _GEN_460 : btb_pc_5; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1206 = fb_reg_valid ? _GEN_461 : btb_pc_6; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1207 = fb_reg_valid ? _GEN_462 : btb_pc_7; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1208 = fb_reg_valid ? _GEN_463 : btb_pc_8; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1209 = fb_reg_valid ? _GEN_464 : btb_pc_9; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1210 = fb_reg_valid ? _GEN_465 : btb_pc_10; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1211 = fb_reg_valid ? _GEN_466 : btb_pc_11; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1212 = fb_reg_valid ? _GEN_467 : btb_pc_12; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1213 = fb_reg_valid ? _GEN_468 : btb_pc_13; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1214 = fb_reg_valid ? _GEN_469 : btb_pc_14; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1215 = fb_reg_valid ? _GEN_470 : btb_pc_15; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1216 = fb_reg_valid ? _GEN_471 : btb_pc_16; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1217 = fb_reg_valid ? _GEN_472 : btb_pc_17; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1218 = fb_reg_valid ? _GEN_473 : btb_pc_18; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1219 = fb_reg_valid ? _GEN_474 : btb_pc_19; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1220 = fb_reg_valid ? _GEN_475 : btb_pc_20; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1221 = fb_reg_valid ? _GEN_476 : btb_pc_21; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1222 = fb_reg_valid ? _GEN_477 : btb_pc_22; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1223 = fb_reg_valid ? _GEN_478 : btb_pc_23; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1224 = fb_reg_valid ? _GEN_479 : btb_pc_24; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1225 = fb_reg_valid ? _GEN_480 : btb_pc_25; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1226 = fb_reg_valid ? _GEN_481 : btb_pc_26; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1227 = fb_reg_valid ? _GEN_482 : btb_pc_27; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1228 = fb_reg_valid ? _GEN_483 : btb_pc_28; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1229 = fb_reg_valid ? _GEN_484 : btb_pc_29; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1230 = fb_reg_valid ? _GEN_485 : btb_pc_30; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1231 = fb_reg_valid ? _GEN_486 : btb_pc_31; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1232 = fb_reg_valid ? _GEN_487 : btb_pc_32; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1233 = fb_reg_valid ? _GEN_488 : btb_pc_33; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1234 = fb_reg_valid ? _GEN_489 : btb_pc_34; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1235 = fb_reg_valid ? _GEN_490 : btb_pc_35; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1236 = fb_reg_valid ? _GEN_491 : btb_pc_36; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1237 = fb_reg_valid ? _GEN_492 : btb_pc_37; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1238 = fb_reg_valid ? _GEN_493 : btb_pc_38; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1239 = fb_reg_valid ? _GEN_494 : btb_pc_39; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1240 = fb_reg_valid ? _GEN_495 : btb_pc_40; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1241 = fb_reg_valid ? _GEN_496 : btb_pc_41; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1242 = fb_reg_valid ? _GEN_497 : btb_pc_42; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1243 = fb_reg_valid ? _GEN_498 : btb_pc_43; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1244 = fb_reg_valid ? _GEN_499 : btb_pc_44; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1245 = fb_reg_valid ? _GEN_500 : btb_pc_45; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1246 = fb_reg_valid ? _GEN_501 : btb_pc_46; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1247 = fb_reg_valid ? _GEN_502 : btb_pc_47; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1248 = fb_reg_valid ? _GEN_503 : btb_pc_48; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1249 = fb_reg_valid ? _GEN_504 : btb_pc_49; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1250 = fb_reg_valid ? _GEN_505 : btb_pc_50; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1251 = fb_reg_valid ? _GEN_506 : btb_pc_51; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1252 = fb_reg_valid ? _GEN_507 : btb_pc_52; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1253 = fb_reg_valid ? _GEN_508 : btb_pc_53; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1254 = fb_reg_valid ? _GEN_509 : btb_pc_54; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1255 = fb_reg_valid ? _GEN_510 : btb_pc_55; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1256 = fb_reg_valid ? _GEN_511 : btb_pc_56; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1257 = fb_reg_valid ? _GEN_512 : btb_pc_57; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1258 = fb_reg_valid ? _GEN_513 : btb_pc_58; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1259 = fb_reg_valid ? _GEN_514 : btb_pc_59; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1260 = fb_reg_valid ? _GEN_515 : btb_pc_60; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1261 = fb_reg_valid ? _GEN_516 : btb_pc_61; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1262 = fb_reg_valid ? _GEN_517 : btb_pc_62; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1263 = fb_reg_valid ? _GEN_518 : btb_pc_63; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1264 = fb_reg_valid ? _GEN_519 : btb_tgt_0; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1265 = fb_reg_valid ? _GEN_520 : btb_tgt_1; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1266 = fb_reg_valid ? _GEN_521 : btb_tgt_2; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1267 = fb_reg_valid ? _GEN_522 : btb_tgt_3; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1268 = fb_reg_valid ? _GEN_523 : btb_tgt_4; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1269 = fb_reg_valid ? _GEN_524 : btb_tgt_5; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1270 = fb_reg_valid ? _GEN_525 : btb_tgt_6; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1271 = fb_reg_valid ? _GEN_526 : btb_tgt_7; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1272 = fb_reg_valid ? _GEN_527 : btb_tgt_8; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1273 = fb_reg_valid ? _GEN_528 : btb_tgt_9; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1274 = fb_reg_valid ? _GEN_529 : btb_tgt_10; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1275 = fb_reg_valid ? _GEN_530 : btb_tgt_11; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1276 = fb_reg_valid ? _GEN_531 : btb_tgt_12; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1277 = fb_reg_valid ? _GEN_532 : btb_tgt_13; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1278 = fb_reg_valid ? _GEN_533 : btb_tgt_14; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1279 = fb_reg_valid ? _GEN_534 : btb_tgt_15; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1280 = fb_reg_valid ? _GEN_535 : btb_tgt_16; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1281 = fb_reg_valid ? _GEN_536 : btb_tgt_17; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1282 = fb_reg_valid ? _GEN_537 : btb_tgt_18; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1283 = fb_reg_valid ? _GEN_538 : btb_tgt_19; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1284 = fb_reg_valid ? _GEN_539 : btb_tgt_20; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1285 = fb_reg_valid ? _GEN_540 : btb_tgt_21; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1286 = fb_reg_valid ? _GEN_541 : btb_tgt_22; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1287 = fb_reg_valid ? _GEN_542 : btb_tgt_23; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1288 = fb_reg_valid ? _GEN_543 : btb_tgt_24; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1289 = fb_reg_valid ? _GEN_544 : btb_tgt_25; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1290 = fb_reg_valid ? _GEN_545 : btb_tgt_26; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1291 = fb_reg_valid ? _GEN_546 : btb_tgt_27; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1292 = fb_reg_valid ? _GEN_547 : btb_tgt_28; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1293 = fb_reg_valid ? _GEN_548 : btb_tgt_29; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1294 = fb_reg_valid ? _GEN_549 : btb_tgt_30; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1295 = fb_reg_valid ? _GEN_550 : btb_tgt_31; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1296 = fb_reg_valid ? _GEN_551 : btb_tgt_32; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1297 = fb_reg_valid ? _GEN_552 : btb_tgt_33; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1298 = fb_reg_valid ? _GEN_553 : btb_tgt_34; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1299 = fb_reg_valid ? _GEN_554 : btb_tgt_35; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1300 = fb_reg_valid ? _GEN_555 : btb_tgt_36; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1301 = fb_reg_valid ? _GEN_556 : btb_tgt_37; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1302 = fb_reg_valid ? _GEN_557 : btb_tgt_38; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1303 = fb_reg_valid ? _GEN_558 : btb_tgt_39; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1304 = fb_reg_valid ? _GEN_559 : btb_tgt_40; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1305 = fb_reg_valid ? _GEN_560 : btb_tgt_41; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1306 = fb_reg_valid ? _GEN_561 : btb_tgt_42; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1307 = fb_reg_valid ? _GEN_562 : btb_tgt_43; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1308 = fb_reg_valid ? _GEN_563 : btb_tgt_44; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1309 = fb_reg_valid ? _GEN_564 : btb_tgt_45; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1310 = fb_reg_valid ? _GEN_565 : btb_tgt_46; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1311 = fb_reg_valid ? _GEN_566 : btb_tgt_47; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1312 = fb_reg_valid ? _GEN_567 : btb_tgt_48; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1313 = fb_reg_valid ? _GEN_568 : btb_tgt_49; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1314 = fb_reg_valid ? _GEN_569 : btb_tgt_50; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1315 = fb_reg_valid ? _GEN_570 : btb_tgt_51; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1316 = fb_reg_valid ? _GEN_571 : btb_tgt_52; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1317 = fb_reg_valid ? _GEN_572 : btb_tgt_53; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1318 = fb_reg_valid ? _GEN_573 : btb_tgt_54; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1319 = fb_reg_valid ? _GEN_574 : btb_tgt_55; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1320 = fb_reg_valid ? _GEN_575 : btb_tgt_56; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1321 = fb_reg_valid ? _GEN_576 : btb_tgt_57; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1322 = fb_reg_valid ? _GEN_577 : btb_tgt_58; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1323 = fb_reg_valid ? _GEN_578 : btb_tgt_59; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1324 = fb_reg_valid ? _GEN_579 : btb_tgt_60; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1325 = fb_reg_valid ? _GEN_580 : btb_tgt_61; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1326 = fb_reg_valid ? _GEN_581 : btb_tgt_62; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1327 = fb_reg_valid ? _GEN_582 : btb_tgt_63; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1328 = fb_reg_valid ? _GEN_583 : btb_bj_type_0; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1329 = fb_reg_valid ? _GEN_584 : btb_bj_type_1; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1330 = fb_reg_valid ? _GEN_585 : btb_bj_type_2; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1331 = fb_reg_valid ? _GEN_586 : btb_bj_type_3; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1332 = fb_reg_valid ? _GEN_587 : btb_bj_type_4; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1333 = fb_reg_valid ? _GEN_588 : btb_bj_type_5; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1334 = fb_reg_valid ? _GEN_589 : btb_bj_type_6; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1335 = fb_reg_valid ? _GEN_590 : btb_bj_type_7; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1336 = fb_reg_valid ? _GEN_591 : btb_bj_type_8; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1337 = fb_reg_valid ? _GEN_592 : btb_bj_type_9; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1338 = fb_reg_valid ? _GEN_593 : btb_bj_type_10; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1339 = fb_reg_valid ? _GEN_594 : btb_bj_type_11; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1340 = fb_reg_valid ? _GEN_595 : btb_bj_type_12; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1341 = fb_reg_valid ? _GEN_596 : btb_bj_type_13; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1342 = fb_reg_valid ? _GEN_597 : btb_bj_type_14; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1343 = fb_reg_valid ? _GEN_598 : btb_bj_type_15; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1344 = fb_reg_valid ? _GEN_599 : btb_bj_type_16; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1345 = fb_reg_valid ? _GEN_600 : btb_bj_type_17; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1346 = fb_reg_valid ? _GEN_601 : btb_bj_type_18; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1347 = fb_reg_valid ? _GEN_602 : btb_bj_type_19; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1348 = fb_reg_valid ? _GEN_603 : btb_bj_type_20; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1349 = fb_reg_valid ? _GEN_604 : btb_bj_type_21; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1350 = fb_reg_valid ? _GEN_605 : btb_bj_type_22; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1351 = fb_reg_valid ? _GEN_606 : btb_bj_type_23; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1352 = fb_reg_valid ? _GEN_607 : btb_bj_type_24; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1353 = fb_reg_valid ? _GEN_608 : btb_bj_type_25; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1354 = fb_reg_valid ? _GEN_609 : btb_bj_type_26; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1355 = fb_reg_valid ? _GEN_610 : btb_bj_type_27; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1356 = fb_reg_valid ? _GEN_611 : btb_bj_type_28; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1357 = fb_reg_valid ? _GEN_612 : btb_bj_type_29; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1358 = fb_reg_valid ? _GEN_613 : btb_bj_type_30; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1359 = fb_reg_valid ? _GEN_614 : btb_bj_type_31; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1360 = fb_reg_valid ? _GEN_615 : btb_bj_type_32; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1361 = fb_reg_valid ? _GEN_616 : btb_bj_type_33; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1362 = fb_reg_valid ? _GEN_617 : btb_bj_type_34; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1363 = fb_reg_valid ? _GEN_618 : btb_bj_type_35; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1364 = fb_reg_valid ? _GEN_619 : btb_bj_type_36; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1365 = fb_reg_valid ? _GEN_620 : btb_bj_type_37; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1366 = fb_reg_valid ? _GEN_621 : btb_bj_type_38; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1367 = fb_reg_valid ? _GEN_622 : btb_bj_type_39; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1368 = fb_reg_valid ? _GEN_623 : btb_bj_type_40; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1369 = fb_reg_valid ? _GEN_624 : btb_bj_type_41; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1370 = fb_reg_valid ? _GEN_625 : btb_bj_type_42; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1371 = fb_reg_valid ? _GEN_626 : btb_bj_type_43; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1372 = fb_reg_valid ? _GEN_627 : btb_bj_type_44; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1373 = fb_reg_valid ? _GEN_628 : btb_bj_type_45; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1374 = fb_reg_valid ? _GEN_629 : btb_bj_type_46; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1375 = fb_reg_valid ? _GEN_630 : btb_bj_type_47; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1376 = fb_reg_valid ? _GEN_631 : btb_bj_type_48; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1377 = fb_reg_valid ? _GEN_632 : btb_bj_type_49; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1378 = fb_reg_valid ? _GEN_633 : btb_bj_type_50; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1379 = fb_reg_valid ? _GEN_634 : btb_bj_type_51; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1380 = fb_reg_valid ? _GEN_635 : btb_bj_type_52; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1381 = fb_reg_valid ? _GEN_636 : btb_bj_type_53; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1382 = fb_reg_valid ? _GEN_637 : btb_bj_type_54; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1383 = fb_reg_valid ? _GEN_638 : btb_bj_type_55; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1384 = fb_reg_valid ? _GEN_639 : btb_bj_type_56; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1385 = fb_reg_valid ? _GEN_640 : btb_bj_type_57; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1386 = fb_reg_valid ? _GEN_641 : btb_bj_type_58; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1387 = fb_reg_valid ? _GEN_642 : btb_bj_type_59; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1388 = fb_reg_valid ? _GEN_643 : btb_bj_type_60; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1389 = fb_reg_valid ? _GEN_644 : btb_bj_type_61; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1390 = fb_reg_valid ? _GEN_645 : btb_bj_type_62; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1391 = fb_reg_valid ? _GEN_646 : btb_bj_type_63; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1392 = fb_reg_valid ? _GEN_1057 : btb_h_count_0; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1393 = fb_reg_valid ? _GEN_1058 : btb_h_count_1; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1394 = fb_reg_valid ? _GEN_1059 : btb_h_count_2; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1395 = fb_reg_valid ? _GEN_1060 : btb_h_count_3; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1396 = fb_reg_valid ? _GEN_1061 : btb_h_count_4; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1397 = fb_reg_valid ? _GEN_1062 : btb_h_count_5; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1398 = fb_reg_valid ? _GEN_1063 : btb_h_count_6; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1399 = fb_reg_valid ? _GEN_1064 : btb_h_count_7; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1400 = fb_reg_valid ? _GEN_1065 : btb_h_count_8; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1401 = fb_reg_valid ? _GEN_1066 : btb_h_count_9; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1402 = fb_reg_valid ? _GEN_1067 : btb_h_count_10; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1403 = fb_reg_valid ? _GEN_1068 : btb_h_count_11; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1404 = fb_reg_valid ? _GEN_1069 : btb_h_count_12; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1405 = fb_reg_valid ? _GEN_1070 : btb_h_count_13; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1406 = fb_reg_valid ? _GEN_1071 : btb_h_count_14; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1407 = fb_reg_valid ? _GEN_1072 : btb_h_count_15; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1408 = fb_reg_valid ? _GEN_1073 : btb_h_count_16; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1409 = fb_reg_valid ? _GEN_1074 : btb_h_count_17; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1410 = fb_reg_valid ? _GEN_1075 : btb_h_count_18; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1411 = fb_reg_valid ? _GEN_1076 : btb_h_count_19; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1412 = fb_reg_valid ? _GEN_1077 : btb_h_count_20; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1413 = fb_reg_valid ? _GEN_1078 : btb_h_count_21; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1414 = fb_reg_valid ? _GEN_1079 : btb_h_count_22; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1415 = fb_reg_valid ? _GEN_1080 : btb_h_count_23; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1416 = fb_reg_valid ? _GEN_1081 : btb_h_count_24; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1417 = fb_reg_valid ? _GEN_1082 : btb_h_count_25; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1418 = fb_reg_valid ? _GEN_1083 : btb_h_count_26; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1419 = fb_reg_valid ? _GEN_1084 : btb_h_count_27; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1420 = fb_reg_valid ? _GEN_1085 : btb_h_count_28; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1421 = fb_reg_valid ? _GEN_1086 : btb_h_count_29; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1422 = fb_reg_valid ? _GEN_1087 : btb_h_count_30; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1423 = fb_reg_valid ? _GEN_1088 : btb_h_count_31; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1424 = fb_reg_valid ? _GEN_1089 : btb_h_count_32; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1425 = fb_reg_valid ? _GEN_1090 : btb_h_count_33; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1426 = fb_reg_valid ? _GEN_1091 : btb_h_count_34; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1427 = fb_reg_valid ? _GEN_1092 : btb_h_count_35; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1428 = fb_reg_valid ? _GEN_1093 : btb_h_count_36; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1429 = fb_reg_valid ? _GEN_1094 : btb_h_count_37; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1430 = fb_reg_valid ? _GEN_1095 : btb_h_count_38; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1431 = fb_reg_valid ? _GEN_1096 : btb_h_count_39; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1432 = fb_reg_valid ? _GEN_1097 : btb_h_count_40; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1433 = fb_reg_valid ? _GEN_1098 : btb_h_count_41; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1434 = fb_reg_valid ? _GEN_1099 : btb_h_count_42; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1435 = fb_reg_valid ? _GEN_1100 : btb_h_count_43; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1436 = fb_reg_valid ? _GEN_1101 : btb_h_count_44; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1437 = fb_reg_valid ? _GEN_1102 : btb_h_count_45; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1438 = fb_reg_valid ? _GEN_1103 : btb_h_count_46; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1439 = fb_reg_valid ? _GEN_1104 : btb_h_count_47; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1440 = fb_reg_valid ? _GEN_1105 : btb_h_count_48; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1441 = fb_reg_valid ? _GEN_1106 : btb_h_count_49; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1442 = fb_reg_valid ? _GEN_1107 : btb_h_count_50; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1443 = fb_reg_valid ? _GEN_1108 : btb_h_count_51; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1444 = fb_reg_valid ? _GEN_1109 : btb_h_count_52; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1445 = fb_reg_valid ? _GEN_1110 : btb_h_count_53; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1446 = fb_reg_valid ? _GEN_1111 : btb_h_count_54; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1447 = fb_reg_valid ? _GEN_1112 : btb_h_count_55; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1448 = fb_reg_valid ? _GEN_1113 : btb_h_count_56; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1449 = fb_reg_valid ? _GEN_1114 : btb_h_count_57; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1450 = fb_reg_valid ? _GEN_1115 : btb_h_count_58; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1451 = fb_reg_valid ? _GEN_1116 : btb_h_count_59; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1452 = fb_reg_valid ? _GEN_1117 : btb_h_count_60; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1453 = fb_reg_valid ? _GEN_1118 : btb_h_count_61; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1454 = fb_reg_valid ? _GEN_1119 : btb_h_count_62; // @[BTB.scala 183:23:@2062.4]
  assign _GEN_1455 = fb_reg_valid ? _GEN_1120 : btb_h_count_63; // @[BTB.scala 183:23:@2062.4]
  assign _T_2181 = fb_reg_miss & _T_1776; // @[BTB.scala 212:21:@2128.4]
  assign _T_2183 = arb_gshare_sel_data == 1'h0; // @[BTB.scala 213:26:@2130.6]
  assign _T_2184 = fb_reg_diff & _T_2183; // @[BTB.scala 213:23:@2131.6]
  assign _GEN_1477 = _T_2184 ? 1'h0 : 1'h1; // @[BTB.scala 213:39:@2132.6]
  assign _T_2191 = predict_lookup[63:32]; // @[OneHot.scala 26:18:@2143.6]
  assign _T_2192 = predict_lookup[31:0]; // @[OneHot.scala 27:18:@2144.6]
  assign _T_2194 = _T_2191 != 32'h0; // @[OneHot.scala 28:14:@2145.6]
  assign _T_2195 = _T_2191 | _T_2192; // @[OneHot.scala 28:28:@2146.6]
  assign _T_2196 = _T_2195[31:16]; // @[OneHot.scala 26:18:@2147.6]
  assign _T_2197 = _T_2195[15:0]; // @[OneHot.scala 27:18:@2148.6]
  assign _T_2199 = _T_2196 != 16'h0; // @[OneHot.scala 28:14:@2149.6]
  assign _T_2200 = _T_2196 | _T_2197; // @[OneHot.scala 28:28:@2150.6]
  assign _T_2201 = _T_2200[15:8]; // @[OneHot.scala 26:18:@2151.6]
  assign _T_2202 = _T_2200[7:0]; // @[OneHot.scala 27:18:@2152.6]
  assign _T_2204 = _T_2201 != 8'h0; // @[OneHot.scala 28:14:@2153.6]
  assign _T_2205 = _T_2201 | _T_2202; // @[OneHot.scala 28:28:@2154.6]
  assign _T_2206 = _T_2205[7:4]; // @[OneHot.scala 26:18:@2155.6]
  assign _T_2207 = _T_2205[3:0]; // @[OneHot.scala 27:18:@2156.6]
  assign _T_2209 = _T_2206 != 4'h0; // @[OneHot.scala 28:14:@2157.6]
  assign _T_2210 = _T_2206 | _T_2207; // @[OneHot.scala 28:28:@2158.6]
  assign _T_2211 = _T_2210[3:2]; // @[OneHot.scala 26:18:@2159.6]
  assign _T_2212 = _T_2210[1:0]; // @[OneHot.scala 27:18:@2160.6]
  assign _T_2214 = _T_2211 != 2'h0; // @[OneHot.scala 28:14:@2161.6]
  assign _T_2215 = _T_2211 | _T_2212; // @[OneHot.scala 28:28:@2162.6]
  assign _T_2216 = _T_2215[1]; // @[CircuitMath.scala 30:8:@2163.6]
  assign _T_2221 = {_T_2194,_T_2199,_T_2204,_T_2209,_T_2214,_T_2216}; // @[Cat.scala 30:58:@2168.6]
  assign _T_2224 = reset == 1'h0; // @[BTB.scala 221:11:@2170.6]
  assign _T_2225 = gb_history[0]; // @[BTB.scala 231:47:@2174.6]
  assign _T_2229 = gb_history[1]; // @[BTB.scala 231:47:@2180.6]
  assign _T_2233 = gb_history[2]; // @[BTB.scala 231:47:@2186.6]
  assign _T_2237 = gb_history[3]; // @[BTB.scala 231:47:@2192.6]
  assign _T_2241 = gb_history[4]; // @[BTB.scala 231:47:@2198.6]
  assign _T_2245 = gb_history[5]; // @[BTB.scala 231:47:@2204.6]
  assign _T_2249 = gb_history[6]; // @[BTB.scala 231:47:@2210.6]
  assign _T_2253 = gb_history[7]; // @[BTB.scala 231:47:@2216.6]
  assign _T_2257 = gb_history[8]; // @[BTB.scala 231:47:@2222.6]
  assign _T_2261 = gb_history[9]; // @[BTB.scala 232:26:@2228.6]
  assign io_predict_redirect = _T_1195 & _T_1221; // @[BTB.scala 126:23:@1277.4]
  assign io_predict_history = gb_history; // @[BTB.scala 128:23:@1282.4]
  assign io_predict_diff = _T_1210 ^ _T_1211; // @[BTB.scala 127:23:@1281.4]
  assign io_predict_tgt = _T_1227 ? RAS_io_peek : _T_1237; // @[BTB.scala 129:18:@1293.4]
  assign RAS_clock = clock; // @[:@55.4]
  assign RAS_reset = reset; // @[:@56.4]
  assign RAS_io_push_valid = io_ras_push_valid; // @[BTB.scala 71:12:@59.4]
  assign RAS_io_push_bits = io_ras_push_bits; // @[BTB.scala 71:12:@58.4]
  assign RAS_io_pop = io_ras_pop; // @[BTB.scala 70:12:@57.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    bht[initvar] = _RAND_0[1:0];
  `endif // RANDOMIZE_MEM_INIT
  _RAND_1 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 1024; initvar = initvar+1)
    arb[initvar] = _RAND_1[0:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  gb_history = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  btb_valid_0 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  btb_valid_1 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  btb_valid_2 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  btb_valid_3 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  btb_valid_4 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  btb_valid_5 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  btb_valid_6 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  btb_valid_7 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  btb_valid_8 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  btb_valid_9 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  btb_valid_10 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  btb_valid_11 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  btb_valid_12 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  btb_valid_13 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  btb_valid_14 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  btb_valid_15 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  btb_valid_16 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  btb_valid_17 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  btb_valid_18 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  btb_valid_19 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  btb_valid_20 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  btb_valid_21 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  btb_valid_22 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  btb_valid_23 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  btb_valid_24 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  btb_valid_25 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  btb_valid_26 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  btb_valid_27 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  btb_valid_28 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  btb_valid_29 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  btb_valid_30 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  btb_valid_31 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  btb_valid_32 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  btb_valid_33 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  btb_valid_34 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  btb_valid_35 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  btb_valid_36 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  btb_valid_37 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  btb_valid_38 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  btb_valid_39 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  btb_valid_40 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  btb_valid_41 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  btb_valid_42 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  btb_valid_43 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  btb_valid_44 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  btb_valid_45 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  btb_valid_46 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  btb_valid_47 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  btb_valid_48 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  btb_valid_49 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  btb_valid_50 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  btb_valid_51 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  btb_valid_52 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  btb_valid_53 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  btb_valid_54 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  btb_valid_55 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  btb_valid_56 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  btb_valid_57 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  btb_valid_58 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  btb_valid_59 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  btb_valid_60 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  btb_valid_61 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  btb_valid_62 = _RAND_65[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  btb_valid_63 = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  btb_pc_0 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  btb_pc_1 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  btb_pc_2 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  btb_pc_3 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  btb_pc_4 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  btb_pc_5 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  btb_pc_6 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  btb_pc_7 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  btb_pc_8 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  btb_pc_9 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  btb_pc_10 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  btb_pc_11 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  btb_pc_12 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  btb_pc_13 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  btb_pc_14 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  btb_pc_15 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  btb_pc_16 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  btb_pc_17 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  btb_pc_18 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  btb_pc_19 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  btb_pc_20 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  btb_pc_21 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  btb_pc_22 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  btb_pc_23 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  btb_pc_24 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  btb_pc_25 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  btb_pc_26 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  btb_pc_27 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  btb_pc_28 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  btb_pc_29 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  btb_pc_30 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  btb_pc_31 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  btb_pc_32 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  btb_pc_33 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  btb_pc_34 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  btb_pc_35 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  btb_pc_36 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  btb_pc_37 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  btb_pc_38 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  btb_pc_39 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  btb_pc_40 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  btb_pc_41 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  btb_pc_42 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  btb_pc_43 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  btb_pc_44 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  btb_pc_45 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  btb_pc_46 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  btb_pc_47 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  btb_pc_48 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  btb_pc_49 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  btb_pc_50 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  btb_pc_51 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  btb_pc_52 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  btb_pc_53 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  btb_pc_54 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  btb_pc_55 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  btb_pc_56 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  btb_pc_57 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  btb_pc_58 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  btb_pc_59 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  btb_pc_60 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  btb_pc_61 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  btb_pc_62 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  btb_pc_63 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  btb_tgt_0 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  btb_tgt_1 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  btb_tgt_2 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  btb_tgt_3 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  btb_tgt_4 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  btb_tgt_5 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  btb_tgt_6 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  btb_tgt_7 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  btb_tgt_8 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  btb_tgt_9 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  btb_tgt_10 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  btb_tgt_11 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  btb_tgt_12 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  btb_tgt_13 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  btb_tgt_14 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  btb_tgt_15 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  btb_tgt_16 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  btb_tgt_17 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  btb_tgt_18 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  btb_tgt_19 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  btb_tgt_20 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  btb_tgt_21 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  btb_tgt_22 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  btb_tgt_23 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  btb_tgt_24 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  btb_tgt_25 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  btb_tgt_26 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  btb_tgt_27 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  btb_tgt_28 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  btb_tgt_29 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  btb_tgt_30 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  btb_tgt_31 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  btb_tgt_32 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  btb_tgt_33 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  btb_tgt_34 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  btb_tgt_35 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  btb_tgt_36 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  btb_tgt_37 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  btb_tgt_38 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  btb_tgt_39 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  btb_tgt_40 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  btb_tgt_41 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  btb_tgt_42 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  btb_tgt_43 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  btb_tgt_44 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  btb_tgt_45 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  btb_tgt_46 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  btb_tgt_47 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  btb_tgt_48 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  btb_tgt_49 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  btb_tgt_50 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  btb_tgt_51 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  btb_tgt_52 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  btb_tgt_53 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  btb_tgt_54 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  btb_tgt_55 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  btb_tgt_56 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  btb_tgt_57 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  btb_tgt_58 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  btb_tgt_59 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  btb_tgt_60 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  btb_tgt_61 = _RAND_192[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  btb_tgt_62 = _RAND_193[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  btb_tgt_63 = _RAND_194[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  btb_bj_type_0 = _RAND_195[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  btb_bj_type_1 = _RAND_196[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  btb_bj_type_2 = _RAND_197[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  btb_bj_type_3 = _RAND_198[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  btb_bj_type_4 = _RAND_199[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  btb_bj_type_5 = _RAND_200[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  btb_bj_type_6 = _RAND_201[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  btb_bj_type_7 = _RAND_202[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  btb_bj_type_8 = _RAND_203[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  btb_bj_type_9 = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  btb_bj_type_10 = _RAND_205[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  btb_bj_type_11 = _RAND_206[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  btb_bj_type_12 = _RAND_207[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  btb_bj_type_13 = _RAND_208[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  btb_bj_type_14 = _RAND_209[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  btb_bj_type_15 = _RAND_210[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  btb_bj_type_16 = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  btb_bj_type_17 = _RAND_212[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  btb_bj_type_18 = _RAND_213[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  btb_bj_type_19 = _RAND_214[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  btb_bj_type_20 = _RAND_215[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  btb_bj_type_21 = _RAND_216[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  btb_bj_type_22 = _RAND_217[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  btb_bj_type_23 = _RAND_218[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  btb_bj_type_24 = _RAND_219[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  btb_bj_type_25 = _RAND_220[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  btb_bj_type_26 = _RAND_221[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  btb_bj_type_27 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  btb_bj_type_28 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  btb_bj_type_29 = _RAND_224[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  btb_bj_type_30 = _RAND_225[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  btb_bj_type_31 = _RAND_226[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  btb_bj_type_32 = _RAND_227[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  btb_bj_type_33 = _RAND_228[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  btb_bj_type_34 = _RAND_229[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  btb_bj_type_35 = _RAND_230[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  btb_bj_type_36 = _RAND_231[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  btb_bj_type_37 = _RAND_232[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  btb_bj_type_38 = _RAND_233[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  btb_bj_type_39 = _RAND_234[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  btb_bj_type_40 = _RAND_235[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  btb_bj_type_41 = _RAND_236[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  btb_bj_type_42 = _RAND_237[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  btb_bj_type_43 = _RAND_238[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  btb_bj_type_44 = _RAND_239[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  btb_bj_type_45 = _RAND_240[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  btb_bj_type_46 = _RAND_241[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  btb_bj_type_47 = _RAND_242[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  btb_bj_type_48 = _RAND_243[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  btb_bj_type_49 = _RAND_244[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  btb_bj_type_50 = _RAND_245[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  btb_bj_type_51 = _RAND_246[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  btb_bj_type_52 = _RAND_247[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  btb_bj_type_53 = _RAND_248[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  btb_bj_type_54 = _RAND_249[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  btb_bj_type_55 = _RAND_250[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  btb_bj_type_56 = _RAND_251[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  btb_bj_type_57 = _RAND_252[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  btb_bj_type_58 = _RAND_253[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  btb_bj_type_59 = _RAND_254[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  btb_bj_type_60 = _RAND_255[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  btb_bj_type_61 = _RAND_256[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  btb_bj_type_62 = _RAND_257[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  btb_bj_type_63 = _RAND_258[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  btb_h_count_0 = _RAND_259[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  btb_h_count_1 = _RAND_260[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  btb_h_count_2 = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_262 = {1{`RANDOM}};
  btb_h_count_3 = _RAND_262[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_263 = {1{`RANDOM}};
  btb_h_count_4 = _RAND_263[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_264 = {1{`RANDOM}};
  btb_h_count_5 = _RAND_264[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_265 = {1{`RANDOM}};
  btb_h_count_6 = _RAND_265[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_266 = {1{`RANDOM}};
  btb_h_count_7 = _RAND_266[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_267 = {1{`RANDOM}};
  btb_h_count_8 = _RAND_267[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_268 = {1{`RANDOM}};
  btb_h_count_9 = _RAND_268[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_269 = {1{`RANDOM}};
  btb_h_count_10 = _RAND_269[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_270 = {1{`RANDOM}};
  btb_h_count_11 = _RAND_270[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_271 = {1{`RANDOM}};
  btb_h_count_12 = _RAND_271[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_272 = {1{`RANDOM}};
  btb_h_count_13 = _RAND_272[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_273 = {1{`RANDOM}};
  btb_h_count_14 = _RAND_273[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_274 = {1{`RANDOM}};
  btb_h_count_15 = _RAND_274[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_275 = {1{`RANDOM}};
  btb_h_count_16 = _RAND_275[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_276 = {1{`RANDOM}};
  btb_h_count_17 = _RAND_276[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_277 = {1{`RANDOM}};
  btb_h_count_18 = _RAND_277[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_278 = {1{`RANDOM}};
  btb_h_count_19 = _RAND_278[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_279 = {1{`RANDOM}};
  btb_h_count_20 = _RAND_279[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_280 = {1{`RANDOM}};
  btb_h_count_21 = _RAND_280[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_281 = {1{`RANDOM}};
  btb_h_count_22 = _RAND_281[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_282 = {1{`RANDOM}};
  btb_h_count_23 = _RAND_282[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_283 = {1{`RANDOM}};
  btb_h_count_24 = _RAND_283[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_284 = {1{`RANDOM}};
  btb_h_count_25 = _RAND_284[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_285 = {1{`RANDOM}};
  btb_h_count_26 = _RAND_285[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_286 = {1{`RANDOM}};
  btb_h_count_27 = _RAND_286[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_287 = {1{`RANDOM}};
  btb_h_count_28 = _RAND_287[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_288 = {1{`RANDOM}};
  btb_h_count_29 = _RAND_288[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_289 = {1{`RANDOM}};
  btb_h_count_30 = _RAND_289[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_290 = {1{`RANDOM}};
  btb_h_count_31 = _RAND_290[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_291 = {1{`RANDOM}};
  btb_h_count_32 = _RAND_291[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_292 = {1{`RANDOM}};
  btb_h_count_33 = _RAND_292[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_293 = {1{`RANDOM}};
  btb_h_count_34 = _RAND_293[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_294 = {1{`RANDOM}};
  btb_h_count_35 = _RAND_294[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_295 = {1{`RANDOM}};
  btb_h_count_36 = _RAND_295[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_296 = {1{`RANDOM}};
  btb_h_count_37 = _RAND_296[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_297 = {1{`RANDOM}};
  btb_h_count_38 = _RAND_297[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_298 = {1{`RANDOM}};
  btb_h_count_39 = _RAND_298[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_299 = {1{`RANDOM}};
  btb_h_count_40 = _RAND_299[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_300 = {1{`RANDOM}};
  btb_h_count_41 = _RAND_300[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_301 = {1{`RANDOM}};
  btb_h_count_42 = _RAND_301[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_302 = {1{`RANDOM}};
  btb_h_count_43 = _RAND_302[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_303 = {1{`RANDOM}};
  btb_h_count_44 = _RAND_303[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_304 = {1{`RANDOM}};
  btb_h_count_45 = _RAND_304[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_305 = {1{`RANDOM}};
  btb_h_count_46 = _RAND_305[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_306 = {1{`RANDOM}};
  btb_h_count_47 = _RAND_306[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_307 = {1{`RANDOM}};
  btb_h_count_48 = _RAND_307[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_308 = {1{`RANDOM}};
  btb_h_count_49 = _RAND_308[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_309 = {1{`RANDOM}};
  btb_h_count_50 = _RAND_309[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_310 = {1{`RANDOM}};
  btb_h_count_51 = _RAND_310[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_311 = {1{`RANDOM}};
  btb_h_count_52 = _RAND_311[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_312 = {1{`RANDOM}};
  btb_h_count_53 = _RAND_312[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_313 = {1{`RANDOM}};
  btb_h_count_54 = _RAND_313[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_314 = {1{`RANDOM}};
  btb_h_count_55 = _RAND_314[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_315 = {1{`RANDOM}};
  btb_h_count_56 = _RAND_315[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_316 = {1{`RANDOM}};
  btb_h_count_57 = _RAND_316[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_317 = {1{`RANDOM}};
  btb_h_count_58 = _RAND_317[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_318 = {1{`RANDOM}};
  btb_h_count_59 = _RAND_318[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_319 = {1{`RANDOM}};
  btb_h_count_60 = _RAND_319[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_320 = {1{`RANDOM}};
  btb_h_count_61 = _RAND_320[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_321 = {1{`RANDOM}};
  btb_h_count_62 = _RAND_321[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_322 = {1{`RANDOM}};
  btb_h_count_63 = _RAND_322[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_323 = {1{`RANDOM}};
  shift_reg = _RAND_323[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_324 = {1{`RANDOM}};
  fb_reg_valid = _RAND_324[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_325 = {1{`RANDOM}};
  fb_reg_miss = _RAND_325[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_326 = {1{`RANDOM}};
  fb_reg_redirect = _RAND_326[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_327 = {1{`RANDOM}};
  fb_reg_btb_type = _RAND_327[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_328 = {1{`RANDOM}};
  fb_reg_pc = _RAND_328[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_329 = {1{`RANDOM}};
  fb_reg_tgt = _RAND_329[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_330 = {1{`RANDOM}};
  fb_reg_diff = _RAND_330[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_331 = {1{`RANDOM}};
  fb_reg_gshare = _RAND_331[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_332 = {1{`RANDOM}};
  fb_reg_lfsr = _RAND_332[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(bht__T_2148_en & bht__T_2148_mask) begin
      bht[bht__T_2148_addr] <= bht__T_2148_data; // @[BTB.scala 67:16:@52.4]
    end
    if(bht__T_2166_en & bht__T_2166_mask) begin
      bht[bht__T_2166_addr] <= bht__T_2166_data; // @[BTB.scala 67:16:@52.4]
    end
    if(bht__T_2177_en & bht__T_2177_mask) begin
      bht[bht__T_2177_addr] <= bht__T_2177_data; // @[BTB.scala 67:16:@52.4]
    end
    if(arb__T_2185_en & arb__T_2185_mask) begin
      arb[arb__T_2185_addr] <= arb__T_2185_data; // @[BTB.scala 68:16:@53.4]
    end
    if(arb__T_2187_en & arb__T_2187_mask) begin
      arb[arb__T_2187_addr] <= arb__T_2187_data; // @[BTB.scala 68:16:@53.4]
    end
    if (reset) begin
      gb_history <= 10'h0;
    end else begin
      if (io_fb_miss) begin
        if (_T_1191) begin
          gb_history <= _T_1193;
        end else begin
          gb_history <= io_feedBack_history;
        end
      end else begin
        if (io_forward) begin
          if (shift_wire) begin
            gb_history <= _T_1203;
          end else begin
            if (_T_1198) begin
              gb_history <= _T_1213;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_0 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_valid_0 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h0 == feedback_idx) begin
              btb_valid_0 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_1 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_valid_1 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1 == feedback_idx) begin
              btb_valid_1 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_2 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_valid_2 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2 == feedback_idx) begin
              btb_valid_2 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_3 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_valid_3 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3 == feedback_idx) begin
              btb_valid_3 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_4 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_valid_4 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h4 == feedback_idx) begin
              btb_valid_4 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_5 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_valid_5 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h5 == feedback_idx) begin
              btb_valid_5 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_6 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_valid_6 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h6 == feedback_idx) begin
              btb_valid_6 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_7 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_valid_7 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h7 == feedback_idx) begin
              btb_valid_7 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_8 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_valid_8 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h8 == feedback_idx) begin
              btb_valid_8 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_9 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_valid_9 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h9 == feedback_idx) begin
              btb_valid_9 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_10 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_valid_10 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'ha == feedback_idx) begin
              btb_valid_10 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_11 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_valid_11 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'hb == feedback_idx) begin
              btb_valid_11 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_12 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_valid_12 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'hc == feedback_idx) begin
              btb_valid_12 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_13 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_valid_13 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'hd == feedback_idx) begin
              btb_valid_13 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_14 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_valid_14 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'he == feedback_idx) begin
              btb_valid_14 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_15 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_valid_15 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'hf == feedback_idx) begin
              btb_valid_15 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_16 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_valid_16 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h10 == feedback_idx) begin
              btb_valid_16 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_17 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_valid_17 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h11 == feedback_idx) begin
              btb_valid_17 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_18 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_valid_18 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h12 == feedback_idx) begin
              btb_valid_18 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_19 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_valid_19 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h13 == feedback_idx) begin
              btb_valid_19 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_20 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_valid_20 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h14 == feedback_idx) begin
              btb_valid_20 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_21 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_valid_21 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h15 == feedback_idx) begin
              btb_valid_21 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_22 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_valid_22 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h16 == feedback_idx) begin
              btb_valid_22 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_23 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_valid_23 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h17 == feedback_idx) begin
              btb_valid_23 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_24 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_valid_24 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h18 == feedback_idx) begin
              btb_valid_24 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_25 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_valid_25 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h19 == feedback_idx) begin
              btb_valid_25 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_26 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_valid_26 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1a == feedback_idx) begin
              btb_valid_26 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_27 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_valid_27 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1b == feedback_idx) begin
              btb_valid_27 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_28 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_valid_28 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1c == feedback_idx) begin
              btb_valid_28 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_29 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_valid_29 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1d == feedback_idx) begin
              btb_valid_29 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_30 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_valid_30 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1e == feedback_idx) begin
              btb_valid_30 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_31 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_valid_31 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h1f == feedback_idx) begin
              btb_valid_31 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_32 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_valid_32 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h20 == feedback_idx) begin
              btb_valid_32 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_33 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_valid_33 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h21 == feedback_idx) begin
              btb_valid_33 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_34 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_valid_34 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h22 == feedback_idx) begin
              btb_valid_34 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_35 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_valid_35 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h23 == feedback_idx) begin
              btb_valid_35 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_36 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_valid_36 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h24 == feedback_idx) begin
              btb_valid_36 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_37 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_valid_37 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h25 == feedback_idx) begin
              btb_valid_37 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_38 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_valid_38 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h26 == feedback_idx) begin
              btb_valid_38 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_39 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_valid_39 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h27 == feedback_idx) begin
              btb_valid_39 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_40 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_valid_40 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h28 == feedback_idx) begin
              btb_valid_40 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_41 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_valid_41 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h29 == feedback_idx) begin
              btb_valid_41 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_42 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_valid_42 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2a == feedback_idx) begin
              btb_valid_42 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_43 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_valid_43 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2b == feedback_idx) begin
              btb_valid_43 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_44 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_valid_44 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2c == feedback_idx) begin
              btb_valid_44 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_45 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_valid_45 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2d == feedback_idx) begin
              btb_valid_45 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_46 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_valid_46 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2e == feedback_idx) begin
              btb_valid_46 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_47 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_valid_47 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h2f == feedback_idx) begin
              btb_valid_47 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_48 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_valid_48 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h30 == feedback_idx) begin
              btb_valid_48 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_49 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_valid_49 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h31 == feedback_idx) begin
              btb_valid_49 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_50 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_valid_50 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h32 == feedback_idx) begin
              btb_valid_50 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_51 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_valid_51 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h33 == feedback_idx) begin
              btb_valid_51 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_52 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_valid_52 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h34 == feedback_idx) begin
              btb_valid_52 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_53 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_valid_53 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h35 == feedback_idx) begin
              btb_valid_53 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_54 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_valid_54 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h36 == feedback_idx) begin
              btb_valid_54 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_55 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_valid_55 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h37 == feedback_idx) begin
              btb_valid_55 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_56 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_valid_56 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h38 == feedback_idx) begin
              btb_valid_56 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_57 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_valid_57 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h39 == feedback_idx) begin
              btb_valid_57 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_58 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_valid_58 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3a == feedback_idx) begin
              btb_valid_58 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_59 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_valid_59 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3b == feedback_idx) begin
              btb_valid_59 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_60 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_valid_60 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3c == feedback_idx) begin
              btb_valid_60 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_61 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_valid_61 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3d == feedback_idx) begin
              btb_valid_61 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_62 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_valid_62 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3e == feedback_idx) begin
              btb_valid_62 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_valid_63 <= 1'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_valid_63 <= 1'h1;
          end
        end else begin
          if (_T_1776) begin
            if (6'h3f == feedback_idx) begin
              btb_valid_63 <= _T_2135;
            end
          end
        end
      end
    end
    if (reset) begin
      btb_pc_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_pc_0 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_pc_1 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_pc_2 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_pc_3 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_pc_4 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_pc_5 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_pc_6 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_pc_7 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_pc_8 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_pc_9 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_pc_10 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_pc_11 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_pc_12 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_pc_13 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_pc_14 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_pc_15 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_pc_16 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_pc_17 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_pc_18 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_pc_19 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_pc_20 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_pc_21 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_pc_22 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_pc_23 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_pc_24 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_pc_25 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_pc_26 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_pc_27 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_pc_28 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_pc_29 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_pc_30 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_pc_31 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_pc_32 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_pc_33 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_pc_34 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_pc_35 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_pc_36 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_pc_37 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_pc_38 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_pc_39 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_pc_40 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_pc_41 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_pc_42 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_pc_43 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_pc_44 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_pc_45 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_pc_46 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_pc_47 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_pc_48 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_pc_49 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_pc_50 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_pc_51 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_pc_52 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_pc_53 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_pc_54 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_pc_55 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_pc_56 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_pc_57 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_pc_58 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_pc_59 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_pc_60 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_pc_61 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_pc_62 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_pc_63 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_tgt_0 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_tgt_1 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_tgt_2 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_tgt_3 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_tgt_4 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_tgt_5 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_tgt_6 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_tgt_7 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_tgt_8 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_tgt_9 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_tgt_10 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_tgt_11 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_tgt_12 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_tgt_13 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_tgt_14 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_tgt_15 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_tgt_16 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_tgt_17 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_tgt_18 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_tgt_19 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_tgt_20 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_tgt_21 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_tgt_22 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_tgt_23 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_tgt_24 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_tgt_25 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_tgt_26 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_tgt_27 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_tgt_28 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_tgt_29 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_tgt_30 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_tgt_31 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_tgt_32 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_tgt_33 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_tgt_34 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_tgt_35 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_tgt_36 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_tgt_37 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_tgt_38 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_tgt_39 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_tgt_40 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_tgt_41 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_tgt_42 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_tgt_43 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_tgt_44 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_tgt_45 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_tgt_46 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_tgt_47 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_tgt_48 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_tgt_49 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_tgt_50 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_tgt_51 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_tgt_52 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_tgt_53 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_tgt_54 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_tgt_55 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_tgt_56 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_tgt_57 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_tgt_58 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_tgt_59 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_tgt_60 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_tgt_61 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_tgt_62 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_tgt_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_tgt_63 <= fb_reg_tgt;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == feedback_idx) begin
            btb_bj_type_0 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == feedback_idx) begin
            btb_bj_type_1 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == feedback_idx) begin
            btb_bj_type_2 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == feedback_idx) begin
            btb_bj_type_3 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == feedback_idx) begin
            btb_bj_type_4 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == feedback_idx) begin
            btb_bj_type_5 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == feedback_idx) begin
            btb_bj_type_6 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == feedback_idx) begin
            btb_bj_type_7 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == feedback_idx) begin
            btb_bj_type_8 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == feedback_idx) begin
            btb_bj_type_9 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == feedback_idx) begin
            btb_bj_type_10 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == feedback_idx) begin
            btb_bj_type_11 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == feedback_idx) begin
            btb_bj_type_12 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == feedback_idx) begin
            btb_bj_type_13 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == feedback_idx) begin
            btb_bj_type_14 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == feedback_idx) begin
            btb_bj_type_15 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == feedback_idx) begin
            btb_bj_type_16 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == feedback_idx) begin
            btb_bj_type_17 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == feedback_idx) begin
            btb_bj_type_18 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == feedback_idx) begin
            btb_bj_type_19 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == feedback_idx) begin
            btb_bj_type_20 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == feedback_idx) begin
            btb_bj_type_21 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == feedback_idx) begin
            btb_bj_type_22 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == feedback_idx) begin
            btb_bj_type_23 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == feedback_idx) begin
            btb_bj_type_24 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == feedback_idx) begin
            btb_bj_type_25 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == feedback_idx) begin
            btb_bj_type_26 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == feedback_idx) begin
            btb_bj_type_27 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == feedback_idx) begin
            btb_bj_type_28 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == feedback_idx) begin
            btb_bj_type_29 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == feedback_idx) begin
            btb_bj_type_30 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == feedback_idx) begin
            btb_bj_type_31 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == feedback_idx) begin
            btb_bj_type_32 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == feedback_idx) begin
            btb_bj_type_33 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == feedback_idx) begin
            btb_bj_type_34 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == feedback_idx) begin
            btb_bj_type_35 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == feedback_idx) begin
            btb_bj_type_36 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == feedback_idx) begin
            btb_bj_type_37 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == feedback_idx) begin
            btb_bj_type_38 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == feedback_idx) begin
            btb_bj_type_39 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == feedback_idx) begin
            btb_bj_type_40 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == feedback_idx) begin
            btb_bj_type_41 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == feedback_idx) begin
            btb_bj_type_42 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == feedback_idx) begin
            btb_bj_type_43 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == feedback_idx) begin
            btb_bj_type_44 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == feedback_idx) begin
            btb_bj_type_45 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == feedback_idx) begin
            btb_bj_type_46 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == feedback_idx) begin
            btb_bj_type_47 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == feedback_idx) begin
            btb_bj_type_48 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == feedback_idx) begin
            btb_bj_type_49 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == feedback_idx) begin
            btb_bj_type_50 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == feedback_idx) begin
            btb_bj_type_51 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == feedback_idx) begin
            btb_bj_type_52 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == feedback_idx) begin
            btb_bj_type_53 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == feedback_idx) begin
            btb_bj_type_54 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == feedback_idx) begin
            btb_bj_type_55 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == feedback_idx) begin
            btb_bj_type_56 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == feedback_idx) begin
            btb_bj_type_57 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == feedback_idx) begin
            btb_bj_type_58 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == feedback_idx) begin
            btb_bj_type_59 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == feedback_idx) begin
            btb_bj_type_60 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == feedback_idx) begin
            btb_bj_type_61 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == feedback_idx) begin
            btb_bj_type_62 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_bj_type_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == feedback_idx) begin
            btb_bj_type_63 <= fb_reg_btb_type;
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= _T_2147;
              end
            end else begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h0 == feedback_idx) begin
                btb_h_count_0 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= _T_2147;
              end
            end else begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1 == feedback_idx) begin
                btb_h_count_1 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= _T_2147;
              end
            end else begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2 == feedback_idx) begin
                btb_h_count_2 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= _T_2147;
              end
            end else begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3 == feedback_idx) begin
                btb_h_count_3 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= _T_2147;
              end
            end else begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h4 == feedback_idx) begin
                btb_h_count_4 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= _T_2147;
              end
            end else begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h5 == feedback_idx) begin
                btb_h_count_5 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= _T_2147;
              end
            end else begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h6 == feedback_idx) begin
                btb_h_count_6 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= _T_2147;
              end
            end else begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h7 == feedback_idx) begin
                btb_h_count_7 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= _T_2147;
              end
            end else begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h8 == feedback_idx) begin
                btb_h_count_8 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= _T_2147;
              end
            end else begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h9 == feedback_idx) begin
                btb_h_count_9 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= _T_2147;
              end
            end else begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'ha == feedback_idx) begin
                btb_h_count_10 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= _T_2147;
              end
            end else begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hb == feedback_idx) begin
                btb_h_count_11 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= _T_2147;
              end
            end else begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hc == feedback_idx) begin
                btb_h_count_12 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= _T_2147;
              end
            end else begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hd == feedback_idx) begin
                btb_h_count_13 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= _T_2147;
              end
            end else begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'he == feedback_idx) begin
                btb_h_count_14 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= _T_2147;
              end
            end else begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hf == feedback_idx) begin
                btb_h_count_15 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= _T_2147;
              end
            end else begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h10 == feedback_idx) begin
                btb_h_count_16 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= _T_2147;
              end
            end else begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h11 == feedback_idx) begin
                btb_h_count_17 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= _T_2147;
              end
            end else begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h12 == feedback_idx) begin
                btb_h_count_18 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= _T_2147;
              end
            end else begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h13 == feedback_idx) begin
                btb_h_count_19 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= _T_2147;
              end
            end else begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h14 == feedback_idx) begin
                btb_h_count_20 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= _T_2147;
              end
            end else begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h15 == feedback_idx) begin
                btb_h_count_21 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= _T_2147;
              end
            end else begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h16 == feedback_idx) begin
                btb_h_count_22 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= _T_2147;
              end
            end else begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h17 == feedback_idx) begin
                btb_h_count_23 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= _T_2147;
              end
            end else begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h18 == feedback_idx) begin
                btb_h_count_24 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= _T_2147;
              end
            end else begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h19 == feedback_idx) begin
                btb_h_count_25 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= _T_2147;
              end
            end else begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1a == feedback_idx) begin
                btb_h_count_26 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= _T_2147;
              end
            end else begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1b == feedback_idx) begin
                btb_h_count_27 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= _T_2147;
              end
            end else begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1c == feedback_idx) begin
                btb_h_count_28 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= _T_2147;
              end
            end else begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1d == feedback_idx) begin
                btb_h_count_29 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= _T_2147;
              end
            end else begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1e == feedback_idx) begin
                btb_h_count_30 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= _T_2147;
              end
            end else begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1f == feedback_idx) begin
                btb_h_count_31 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= _T_2147;
              end
            end else begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h20 == feedback_idx) begin
                btb_h_count_32 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= _T_2147;
              end
            end else begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h21 == feedback_idx) begin
                btb_h_count_33 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= _T_2147;
              end
            end else begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h22 == feedback_idx) begin
                btb_h_count_34 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= _T_2147;
              end
            end else begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h23 == feedback_idx) begin
                btb_h_count_35 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= _T_2147;
              end
            end else begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h24 == feedback_idx) begin
                btb_h_count_36 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= _T_2147;
              end
            end else begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h25 == feedback_idx) begin
                btb_h_count_37 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= _T_2147;
              end
            end else begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h26 == feedback_idx) begin
                btb_h_count_38 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= _T_2147;
              end
            end else begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h27 == feedback_idx) begin
                btb_h_count_39 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= _T_2147;
              end
            end else begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h28 == feedback_idx) begin
                btb_h_count_40 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= _T_2147;
              end
            end else begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h29 == feedback_idx) begin
                btb_h_count_41 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= _T_2147;
              end
            end else begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2a == feedback_idx) begin
                btb_h_count_42 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= _T_2147;
              end
            end else begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2b == feedback_idx) begin
                btb_h_count_43 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= _T_2147;
              end
            end else begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2c == feedback_idx) begin
                btb_h_count_44 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= _T_2147;
              end
            end else begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2d == feedback_idx) begin
                btb_h_count_45 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= _T_2147;
              end
            end else begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2e == feedback_idx) begin
                btb_h_count_46 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= _T_2147;
              end
            end else begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2f == feedback_idx) begin
                btb_h_count_47 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= _T_2147;
              end
            end else begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h30 == feedback_idx) begin
                btb_h_count_48 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= _T_2147;
              end
            end else begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h31 == feedback_idx) begin
                btb_h_count_49 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= _T_2147;
              end
            end else begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h32 == feedback_idx) begin
                btb_h_count_50 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= _T_2147;
              end
            end else begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h33 == feedback_idx) begin
                btb_h_count_51 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= _T_2147;
              end
            end else begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h34 == feedback_idx) begin
                btb_h_count_52 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= _T_2147;
              end
            end else begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h35 == feedback_idx) begin
                btb_h_count_53 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= _T_2147;
              end
            end else begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h36 == feedback_idx) begin
                btb_h_count_54 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= _T_2147;
              end
            end else begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h37 == feedback_idx) begin
                btb_h_count_55 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= _T_2147;
              end
            end else begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h38 == feedback_idx) begin
                btb_h_count_56 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= _T_2147;
              end
            end else begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h39 == feedback_idx) begin
                btb_h_count_57 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= _T_2147;
              end
            end else begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3a == feedback_idx) begin
                btb_h_count_58 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= _T_2147;
              end
            end else begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3b == feedback_idx) begin
                btb_h_count_59 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= _T_2147;
              end
            end else begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3c == feedback_idx) begin
                btb_h_count_60 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= _T_2147;
              end
            end else begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3d == feedback_idx) begin
                btb_h_count_61 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= _T_2147;
              end
            end else begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3e == feedback_idx) begin
                btb_h_count_62 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_h_count_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2135) begin
          if (_T_1776) begin
            if (fb_reg_redirect) begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= _T_2147;
              end
            end else begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= _T_2165;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3f == feedback_idx) begin
                btb_h_count_63 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (!(io_fb_miss)) begin
      if (io_forward) begin
        shift_reg <= _T_1200;
      end
    end
    if (reset) begin
      fb_reg_valid <= 1'h0;
    end else begin
      fb_reg_valid <= io_feedBack_valid;
    end
    if (reset) begin
      fb_reg_miss <= 1'h0;
    end else begin
      fb_reg_miss <= io_fb_miss;
    end
    if (reset) begin
      fb_reg_redirect <= 1'h0;
    end else begin
      fb_reg_redirect <= io_feedBack_redirect;
    end
    if (reset) begin
      fb_reg_btb_type <= 2'h0;
    end else begin
      fb_reg_btb_type <= io_fb_type;
    end
    if (reset) begin
      fb_reg_pc <= 32'h0;
    end else begin
      fb_reg_pc <= io_fb_pc;
    end
    if (reset) begin
      fb_reg_tgt <= 32'h0;
    end else begin
      fb_reg_tgt <= io_feedBack_tgt;
    end
    if (reset) begin
      fb_reg_diff <= 1'h0;
    end else begin
      fb_reg_diff <= io_feedBack_diff;
    end
    if (reset) begin
      fb_reg_gshare <= 10'h0;
    end else begin
      fb_reg_gshare <= _T_1248;
    end
    if (reset) begin
      fb_reg_lfsr <= 6'h1;
    end else begin
      fb_reg_lfsr <= _T_1253;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"BTB: Cyc= %d pc %x redirect %x index %d select %d gshare %d hcount %d bht idx %d <",io_cyc,io_if_pc,io_predict_redirect,_T_2221,predict_select,predict_gshare,predict_h_count,gshare_xor); // @[BTB.scala 221:11:@2172.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2225); // @[BTB.scala 231:32:@2178.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2229); // @[BTB.scala 231:32:@2184.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2233); // @[BTB.scala 231:32:@2190.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2237); // @[BTB.scala 231:32:@2196.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2241); // @[BTB.scala 231:32:@2202.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2245); // @[BTB.scala 231:32:@2208.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2249); // @[BTB.scala 231:32:@2214.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2253); // @[BTB.scala 231:32:@2220.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d,",_T_2257); // @[BTB.scala 231:32:@2226.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1195 & _T_2224) begin
          $fwrite(32'h80000002,"%d>\n",_T_2261); // @[BTB.scala 232:11:@2232.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module MyMem( // @[:@2236.2]
  input         clock, // @[:@2237.4]
  input         io_wen, // @[:@2239.4]
  input  [5:0]  io_addr, // @[:@2239.4]
  input  [31:0] io_wdata, // @[:@2239.4]
  output [31:0] io_rdata // @[:@2239.4]
);
  reg [31:0] mem [0:63]; // @[CaheCore.scala 16:24:@2241.4]
  reg [31:0] _RAND_0;
  wire [31:0] mem__T_15_data; // @[CaheCore.scala 16:24:@2241.4]
  wire [5:0] mem__T_15_addr; // @[CaheCore.scala 16:24:@2241.4]
  wire [31:0] mem__T_16_data; // @[CaheCore.scala 16:24:@2241.4]
  wire [5:0] mem__T_16_addr; // @[CaheCore.scala 16:24:@2241.4]
  wire  mem__T_16_mask; // @[CaheCore.scala 16:24:@2241.4]
  wire  mem__T_16_en; // @[CaheCore.scala 16:24:@2241.4]
  wire  _GEN_3; // @[CaheCore.scala 18:17:@2244.4]
  reg [5:0] mem__T_15_addr_pipe_0;
  reg [31:0] _RAND_1;
  assign mem__T_15_addr = mem__T_15_addr_pipe_0;
  assign mem__T_15_data = mem[mem__T_15_addr]; // @[CaheCore.scala 16:24:@2241.4]
  assign mem__T_16_data = io_wdata;
  assign mem__T_16_addr = io_addr;
  assign mem__T_16_mask = 1'h1;
  assign mem__T_16_en = io_wen;
  assign _GEN_3 = 1'h1; // @[CaheCore.scala 18:17:@2244.4]
  assign io_rdata = mem__T_15_data; // @[CaheCore.scala 17:12:@2243.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    mem[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  mem__T_15_addr_pipe_0 = _RAND_1[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(mem__T_16_en & mem__T_16_mask) begin
      mem[mem__T_16_addr] <= mem__T_16_data; // @[CaheCore.scala 16:24:@2241.4]
    end
    if (_GEN_3) begin
      mem__T_15_addr_pipe_0 <= io_addr;
    end
  end
endmodule
module CaheCore( // @[:@2444.2]
  input         clock, // @[:@2445.4]
  input         reset, // @[:@2446.4]
  input         io_wen, // @[:@2447.4]
  input  [31:0] io_addr, // @[:@2447.4]
  input  [31:0] io_wdata_0, // @[:@2447.4]
  input  [31:0] io_wdata_1, // @[:@2447.4]
  input  [31:0] io_wdata_2, // @[:@2447.4]
  input  [31:0] io_wdata_3, // @[:@2447.4]
  input  [31:0] io_wdata_4, // @[:@2447.4]
  input  [31:0] io_wdata_5, // @[:@2447.4]
  input  [31:0] io_wdata_6, // @[:@2447.4]
  input  [31:0] io_wdata_7, // @[:@2447.4]
  input  [31:0] io_wdata_8, // @[:@2447.4]
  input  [31:0] io_wdata_9, // @[:@2447.4]
  input  [31:0] io_wdata_10, // @[:@2447.4]
  input  [31:0] io_wdata_11, // @[:@2447.4]
  input  [31:0] io_wdata_12, // @[:@2447.4]
  input  [31:0] io_wdata_13, // @[:@2447.4]
  input  [31:0] io_wdata_14, // @[:@2447.4]
  input  [31:0] io_wdata_15, // @[:@2447.4]
  input         io_wstatus, // @[:@2447.4]
  output [31:0] io_rdata, // @[:@2447.4]
  output        io_rvalid // @[:@2447.4]
);
  wire  MyMem_clock; // @[CaheCore.scala 34:43:@2449.4]
  wire  MyMem_io_wen; // @[CaheCore.scala 34:43:@2449.4]
  wire [5:0] MyMem_io_addr; // @[CaheCore.scala 34:43:@2449.4]
  wire [31:0] MyMem_io_wdata; // @[CaheCore.scala 34:43:@2449.4]
  wire [31:0] MyMem_io_rdata; // @[CaheCore.scala 34:43:@2449.4]
  wire  MyMem_1_clock; // @[CaheCore.scala 34:43:@2452.4]
  wire  MyMem_1_io_wen; // @[CaheCore.scala 34:43:@2452.4]
  wire [5:0] MyMem_1_io_addr; // @[CaheCore.scala 34:43:@2452.4]
  wire [31:0] MyMem_1_io_wdata; // @[CaheCore.scala 34:43:@2452.4]
  wire [31:0] MyMem_1_io_rdata; // @[CaheCore.scala 34:43:@2452.4]
  wire  MyMem_2_clock; // @[CaheCore.scala 34:43:@2455.4]
  wire  MyMem_2_io_wen; // @[CaheCore.scala 34:43:@2455.4]
  wire [5:0] MyMem_2_io_addr; // @[CaheCore.scala 34:43:@2455.4]
  wire [31:0] MyMem_2_io_wdata; // @[CaheCore.scala 34:43:@2455.4]
  wire [31:0] MyMem_2_io_rdata; // @[CaheCore.scala 34:43:@2455.4]
  wire  MyMem_3_clock; // @[CaheCore.scala 34:43:@2458.4]
  wire  MyMem_3_io_wen; // @[CaheCore.scala 34:43:@2458.4]
  wire [5:0] MyMem_3_io_addr; // @[CaheCore.scala 34:43:@2458.4]
  wire [31:0] MyMem_3_io_wdata; // @[CaheCore.scala 34:43:@2458.4]
  wire [31:0] MyMem_3_io_rdata; // @[CaheCore.scala 34:43:@2458.4]
  wire  MyMem_4_clock; // @[CaheCore.scala 34:43:@2461.4]
  wire  MyMem_4_io_wen; // @[CaheCore.scala 34:43:@2461.4]
  wire [5:0] MyMem_4_io_addr; // @[CaheCore.scala 34:43:@2461.4]
  wire [31:0] MyMem_4_io_wdata; // @[CaheCore.scala 34:43:@2461.4]
  wire [31:0] MyMem_4_io_rdata; // @[CaheCore.scala 34:43:@2461.4]
  wire  MyMem_5_clock; // @[CaheCore.scala 34:43:@2464.4]
  wire  MyMem_5_io_wen; // @[CaheCore.scala 34:43:@2464.4]
  wire [5:0] MyMem_5_io_addr; // @[CaheCore.scala 34:43:@2464.4]
  wire [31:0] MyMem_5_io_wdata; // @[CaheCore.scala 34:43:@2464.4]
  wire [31:0] MyMem_5_io_rdata; // @[CaheCore.scala 34:43:@2464.4]
  wire  MyMem_6_clock; // @[CaheCore.scala 34:43:@2467.4]
  wire  MyMem_6_io_wen; // @[CaheCore.scala 34:43:@2467.4]
  wire [5:0] MyMem_6_io_addr; // @[CaheCore.scala 34:43:@2467.4]
  wire [31:0] MyMem_6_io_wdata; // @[CaheCore.scala 34:43:@2467.4]
  wire [31:0] MyMem_6_io_rdata; // @[CaheCore.scala 34:43:@2467.4]
  wire  MyMem_7_clock; // @[CaheCore.scala 34:43:@2470.4]
  wire  MyMem_7_io_wen; // @[CaheCore.scala 34:43:@2470.4]
  wire [5:0] MyMem_7_io_addr; // @[CaheCore.scala 34:43:@2470.4]
  wire [31:0] MyMem_7_io_wdata; // @[CaheCore.scala 34:43:@2470.4]
  wire [31:0] MyMem_7_io_rdata; // @[CaheCore.scala 34:43:@2470.4]
  wire  MyMem_8_clock; // @[CaheCore.scala 34:43:@2473.4]
  wire  MyMem_8_io_wen; // @[CaheCore.scala 34:43:@2473.4]
  wire [5:0] MyMem_8_io_addr; // @[CaheCore.scala 34:43:@2473.4]
  wire [31:0] MyMem_8_io_wdata; // @[CaheCore.scala 34:43:@2473.4]
  wire [31:0] MyMem_8_io_rdata; // @[CaheCore.scala 34:43:@2473.4]
  wire  MyMem_9_clock; // @[CaheCore.scala 34:43:@2476.4]
  wire  MyMem_9_io_wen; // @[CaheCore.scala 34:43:@2476.4]
  wire [5:0] MyMem_9_io_addr; // @[CaheCore.scala 34:43:@2476.4]
  wire [31:0] MyMem_9_io_wdata; // @[CaheCore.scala 34:43:@2476.4]
  wire [31:0] MyMem_9_io_rdata; // @[CaheCore.scala 34:43:@2476.4]
  wire  MyMem_10_clock; // @[CaheCore.scala 34:43:@2479.4]
  wire  MyMem_10_io_wen; // @[CaheCore.scala 34:43:@2479.4]
  wire [5:0] MyMem_10_io_addr; // @[CaheCore.scala 34:43:@2479.4]
  wire [31:0] MyMem_10_io_wdata; // @[CaheCore.scala 34:43:@2479.4]
  wire [31:0] MyMem_10_io_rdata; // @[CaheCore.scala 34:43:@2479.4]
  wire  MyMem_11_clock; // @[CaheCore.scala 34:43:@2482.4]
  wire  MyMem_11_io_wen; // @[CaheCore.scala 34:43:@2482.4]
  wire [5:0] MyMem_11_io_addr; // @[CaheCore.scala 34:43:@2482.4]
  wire [31:0] MyMem_11_io_wdata; // @[CaheCore.scala 34:43:@2482.4]
  wire [31:0] MyMem_11_io_rdata; // @[CaheCore.scala 34:43:@2482.4]
  wire  MyMem_12_clock; // @[CaheCore.scala 34:43:@2485.4]
  wire  MyMem_12_io_wen; // @[CaheCore.scala 34:43:@2485.4]
  wire [5:0] MyMem_12_io_addr; // @[CaheCore.scala 34:43:@2485.4]
  wire [31:0] MyMem_12_io_wdata; // @[CaheCore.scala 34:43:@2485.4]
  wire [31:0] MyMem_12_io_rdata; // @[CaheCore.scala 34:43:@2485.4]
  wire  MyMem_13_clock; // @[CaheCore.scala 34:43:@2488.4]
  wire  MyMem_13_io_wen; // @[CaheCore.scala 34:43:@2488.4]
  wire [5:0] MyMem_13_io_addr; // @[CaheCore.scala 34:43:@2488.4]
  wire [31:0] MyMem_13_io_wdata; // @[CaheCore.scala 34:43:@2488.4]
  wire [31:0] MyMem_13_io_rdata; // @[CaheCore.scala 34:43:@2488.4]
  wire  MyMem_14_clock; // @[CaheCore.scala 34:43:@2491.4]
  wire  MyMem_14_io_wen; // @[CaheCore.scala 34:43:@2491.4]
  wire [5:0] MyMem_14_io_addr; // @[CaheCore.scala 34:43:@2491.4]
  wire [31:0] MyMem_14_io_wdata; // @[CaheCore.scala 34:43:@2491.4]
  wire [31:0] MyMem_14_io_rdata; // @[CaheCore.scala 34:43:@2491.4]
  wire  MyMem_15_clock; // @[CaheCore.scala 34:43:@2494.4]
  wire  MyMem_15_io_wen; // @[CaheCore.scala 34:43:@2494.4]
  wire [5:0] MyMem_15_io_addr; // @[CaheCore.scala 34:43:@2494.4]
  wire [31:0] MyMem_15_io_wdata; // @[CaheCore.scala 34:43:@2494.4]
  wire [31:0] MyMem_15_io_rdata; // @[CaheCore.scala 34:43:@2494.4]
  reg [19:0] tag_RAM [0:63]; // @[CaheCore.scala 35:30:@2497.4]
  reg [31:0] _RAND_0;
  wire [19:0] tag_RAM_rtag_data; // @[CaheCore.scala 35:30:@2497.4]
  wire [5:0] tag_RAM_rtag_addr; // @[CaheCore.scala 35:30:@2497.4]
  wire [19:0] tag_RAM__T_550_data; // @[CaheCore.scala 35:30:@2497.4]
  wire [5:0] tag_RAM__T_550_addr; // @[CaheCore.scala 35:30:@2497.4]
  wire  tag_RAM__T_550_mask; // @[CaheCore.scala 35:30:@2497.4]
  wire  tag_RAM__T_550_en; // @[CaheCore.scala 35:30:@2497.4]
  reg  statusVec_0; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_1;
  reg  statusVec_1; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_2;
  reg  statusVec_2; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_3;
  reg  statusVec_3; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_4;
  reg  statusVec_4; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_5;
  reg  statusVec_5; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_6;
  reg  statusVec_6; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_7;
  reg  statusVec_7; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_8;
  reg  statusVec_8; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_9;
  reg  statusVec_9; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_10;
  reg  statusVec_10; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_11;
  reg  statusVec_11; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_12;
  reg  statusVec_12; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_13;
  reg  statusVec_13; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_14;
  reg  statusVec_14; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_15;
  reg  statusVec_15; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_16;
  reg  statusVec_16; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_17;
  reg  statusVec_17; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_18;
  reg  statusVec_18; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_19;
  reg  statusVec_19; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_20;
  reg  statusVec_20; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_21;
  reg  statusVec_21; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_22;
  reg  statusVec_22; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_23;
  reg  statusVec_23; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_24;
  reg  statusVec_24; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_25;
  reg  statusVec_25; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_26;
  reg  statusVec_26; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_27;
  reg  statusVec_27; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_28;
  reg  statusVec_28; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_29;
  reg  statusVec_29; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_30;
  reg  statusVec_30; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_31;
  reg  statusVec_31; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_32;
  reg  statusVec_32; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_33;
  reg  statusVec_33; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_34;
  reg  statusVec_34; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_35;
  reg  statusVec_35; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_36;
  reg  statusVec_36; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_37;
  reg  statusVec_37; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_38;
  reg  statusVec_38; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_39;
  reg  statusVec_39; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_40;
  reg  statusVec_40; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_41;
  reg  statusVec_41; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_42;
  reg  statusVec_42; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_43;
  reg  statusVec_43; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_44;
  reg  statusVec_44; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_45;
  reg  statusVec_45; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_46;
  reg  statusVec_46; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_47;
  reg  statusVec_47; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_48;
  reg  statusVec_48; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_49;
  reg  statusVec_49; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_50;
  reg  statusVec_50; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_51;
  reg  statusVec_51; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_52;
  reg  statusVec_52; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_53;
  reg  statusVec_53; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_54;
  reg  statusVec_54; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_55;
  reg  statusVec_55; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_56;
  reg  statusVec_56; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_57;
  reg  statusVec_57; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_58;
  reg  statusVec_58; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_59;
  reg  statusVec_59; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_60;
  reg  statusVec_60; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_61;
  reg  statusVec_61; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_62;
  reg  statusVec_62; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_63;
  reg  statusVec_63; // @[CaheCore.scala 36:26:@2563.4]
  reg [31:0] _RAND_64;
  reg [3:0] line_idx; // @[CaheCore.scala 37:26:@2565.4]
  reg [31:0] _RAND_65;
  wire [5:0] off_idx; // @[CaheCore.scala 40:25:@2568.4]
  reg  rstatus; // @[CaheCore.scala 52:24:@2635.4]
  reg [31:0] _RAND_66;
  wire  _GEN_1; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_2; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_3; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_4; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_5; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_6; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_7; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_8; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_9; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_10; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_11; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_12; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_13; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_14; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_15; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_16; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_17; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_18; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_19; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_20; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_21; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_22; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_23; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_24; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_25; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_26; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_27; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_28; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_29; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_30; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_31; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_32; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_33; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_34; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_35; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_36; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_37; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_38; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_39; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_40; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_41; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_42; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_43; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_44; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_45; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_46; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_47; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_48; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_49; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_50; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_51; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_52; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_53; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_54; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_55; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_56; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_57; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_58; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_59; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_60; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_61; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_62; // @[CaheCore.scala 52:24:@2636.4]
  wire  _GEN_67; // @[CaheCore.scala 54:16:@2637.4]
  wire  _GEN_69; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_70; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_71; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_72; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_73; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_74; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_75; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_76; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_77; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_78; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_79; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_80; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_81; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_82; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_83; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_84; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_85; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_86; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_87; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_88; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_89; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_90; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_91; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_92; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_93; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_94; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_95; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_96; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_97; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_98; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_99; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_100; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_101; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_102; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_103; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_104; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_105; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_106; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_107; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_108; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_109; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_110; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_111; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_112; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_113; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_114; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_115; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_116; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_117; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_118; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_119; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_120; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_121; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_122; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_123; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_124; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_125; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_126; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_127; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_128; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_129; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_130; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_131; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_132; // @[CaheCore.scala 55:37:@2643.6]
  wire  _GEN_133; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_134; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_135; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_136; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_137; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_138; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_139; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_140; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_141; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_142; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_143; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_144; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_145; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_146; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_147; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_148; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_149; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_150; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_151; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_152; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_153; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_154; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_155; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_156; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_157; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_158; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_159; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_160; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_161; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_162; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_163; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_164; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_165; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_166; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_167; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_168; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_169; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_170; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_171; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_172; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_173; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_174; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_175; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_176; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_177; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_178; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_179; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_180; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_181; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_182; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_183; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_184; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_185; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_186; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_187; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_188; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_189; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_190; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_191; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_192; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_193; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_194; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_195; // @[CaheCore.scala 55:16:@2642.4]
  wire  _GEN_196; // @[CaheCore.scala 55:16:@2642.4]
  reg [19:0] tag; // @[CaheCore.scala 57:23:@2645.4]
  reg [31:0] _RAND_67;
  wire [31:0] rdata_0; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2573.4]
  wire [31:0] rdata_1; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2577.4]
  wire [31:0] _GEN_198; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_2; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2581.4]
  wire [31:0] _GEN_199; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_3; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2585.4]
  wire [31:0] _GEN_200; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_4; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2589.4]
  wire [31:0] _GEN_201; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_5; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2593.4]
  wire [31:0] _GEN_202; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_6; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2597.4]
  wire [31:0] _GEN_203; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_7; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2601.4]
  wire [31:0] _GEN_204; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_8; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2605.4]
  wire [31:0] _GEN_205; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_9; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2609.4]
  wire [31:0] _GEN_206; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_10; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2613.4]
  wire [31:0] _GEN_207; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_11; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2617.4]
  wire [31:0] _GEN_208; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_12; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2621.4]
  wire [31:0] _GEN_209; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_13; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2625.4]
  wire [31:0] _GEN_210; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_14; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2629.4]
  wire [31:0] _GEN_211; // @[CaheCore.scala 58:13:@2649.4]
  wire [31:0] rdata_15; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2633.4]
  wire  _T_560; // @[CaheCore.scala 59:21:@2650.4]
  reg [5:0] tag_RAM_rtag_addr_pipe_0;
  reg [31:0] _RAND_68;
  MyMem MyMem ( // @[CaheCore.scala 34:43:@2449.4]
    .clock(MyMem_clock),
    .io_wen(MyMem_io_wen),
    .io_addr(MyMem_io_addr),
    .io_wdata(MyMem_io_wdata),
    .io_rdata(MyMem_io_rdata)
  );
  MyMem MyMem_1 ( // @[CaheCore.scala 34:43:@2452.4]
    .clock(MyMem_1_clock),
    .io_wen(MyMem_1_io_wen),
    .io_addr(MyMem_1_io_addr),
    .io_wdata(MyMem_1_io_wdata),
    .io_rdata(MyMem_1_io_rdata)
  );
  MyMem MyMem_2 ( // @[CaheCore.scala 34:43:@2455.4]
    .clock(MyMem_2_clock),
    .io_wen(MyMem_2_io_wen),
    .io_addr(MyMem_2_io_addr),
    .io_wdata(MyMem_2_io_wdata),
    .io_rdata(MyMem_2_io_rdata)
  );
  MyMem MyMem_3 ( // @[CaheCore.scala 34:43:@2458.4]
    .clock(MyMem_3_clock),
    .io_wen(MyMem_3_io_wen),
    .io_addr(MyMem_3_io_addr),
    .io_wdata(MyMem_3_io_wdata),
    .io_rdata(MyMem_3_io_rdata)
  );
  MyMem MyMem_4 ( // @[CaheCore.scala 34:43:@2461.4]
    .clock(MyMem_4_clock),
    .io_wen(MyMem_4_io_wen),
    .io_addr(MyMem_4_io_addr),
    .io_wdata(MyMem_4_io_wdata),
    .io_rdata(MyMem_4_io_rdata)
  );
  MyMem MyMem_5 ( // @[CaheCore.scala 34:43:@2464.4]
    .clock(MyMem_5_clock),
    .io_wen(MyMem_5_io_wen),
    .io_addr(MyMem_5_io_addr),
    .io_wdata(MyMem_5_io_wdata),
    .io_rdata(MyMem_5_io_rdata)
  );
  MyMem MyMem_6 ( // @[CaheCore.scala 34:43:@2467.4]
    .clock(MyMem_6_clock),
    .io_wen(MyMem_6_io_wen),
    .io_addr(MyMem_6_io_addr),
    .io_wdata(MyMem_6_io_wdata),
    .io_rdata(MyMem_6_io_rdata)
  );
  MyMem MyMem_7 ( // @[CaheCore.scala 34:43:@2470.4]
    .clock(MyMem_7_clock),
    .io_wen(MyMem_7_io_wen),
    .io_addr(MyMem_7_io_addr),
    .io_wdata(MyMem_7_io_wdata),
    .io_rdata(MyMem_7_io_rdata)
  );
  MyMem MyMem_8 ( // @[CaheCore.scala 34:43:@2473.4]
    .clock(MyMem_8_clock),
    .io_wen(MyMem_8_io_wen),
    .io_addr(MyMem_8_io_addr),
    .io_wdata(MyMem_8_io_wdata),
    .io_rdata(MyMem_8_io_rdata)
  );
  MyMem MyMem_9 ( // @[CaheCore.scala 34:43:@2476.4]
    .clock(MyMem_9_clock),
    .io_wen(MyMem_9_io_wen),
    .io_addr(MyMem_9_io_addr),
    .io_wdata(MyMem_9_io_wdata),
    .io_rdata(MyMem_9_io_rdata)
  );
  MyMem MyMem_10 ( // @[CaheCore.scala 34:43:@2479.4]
    .clock(MyMem_10_clock),
    .io_wen(MyMem_10_io_wen),
    .io_addr(MyMem_10_io_addr),
    .io_wdata(MyMem_10_io_wdata),
    .io_rdata(MyMem_10_io_rdata)
  );
  MyMem MyMem_11 ( // @[CaheCore.scala 34:43:@2482.4]
    .clock(MyMem_11_clock),
    .io_wen(MyMem_11_io_wen),
    .io_addr(MyMem_11_io_addr),
    .io_wdata(MyMem_11_io_wdata),
    .io_rdata(MyMem_11_io_rdata)
  );
  MyMem MyMem_12 ( // @[CaheCore.scala 34:43:@2485.4]
    .clock(MyMem_12_clock),
    .io_wen(MyMem_12_io_wen),
    .io_addr(MyMem_12_io_addr),
    .io_wdata(MyMem_12_io_wdata),
    .io_rdata(MyMem_12_io_rdata)
  );
  MyMem MyMem_13 ( // @[CaheCore.scala 34:43:@2488.4]
    .clock(MyMem_13_clock),
    .io_wen(MyMem_13_io_wen),
    .io_addr(MyMem_13_io_addr),
    .io_wdata(MyMem_13_io_wdata),
    .io_rdata(MyMem_13_io_rdata)
  );
  MyMem MyMem_14 ( // @[CaheCore.scala 34:43:@2491.4]
    .clock(MyMem_14_clock),
    .io_wen(MyMem_14_io_wen),
    .io_addr(MyMem_14_io_addr),
    .io_wdata(MyMem_14_io_wdata),
    .io_rdata(MyMem_14_io_rdata)
  );
  MyMem MyMem_15 ( // @[CaheCore.scala 34:43:@2494.4]
    .clock(MyMem_15_clock),
    .io_wen(MyMem_15_io_wen),
    .io_addr(MyMem_15_io_addr),
    .io_wdata(MyMem_15_io_wdata),
    .io_rdata(MyMem_15_io_rdata)
  );
  assign tag_RAM_rtag_addr = tag_RAM_rtag_addr_pipe_0;
  assign tag_RAM_rtag_data = tag_RAM[tag_RAM_rtag_addr]; // @[CaheCore.scala 35:30:@2497.4]
  assign tag_RAM__T_550_data = io_addr[31:12];
  assign tag_RAM__T_550_addr = io_addr[11:6];
  assign tag_RAM__T_550_mask = 1'h1;
  assign tag_RAM__T_550_en = io_wen;
  assign off_idx = io_addr[11:6]; // @[CaheCore.scala 40:25:@2568.4]
  assign _GEN_1 = 6'h1 == off_idx ? statusVec_1 : statusVec_0; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_2 = 6'h2 == off_idx ? statusVec_2 : _GEN_1; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_3 = 6'h3 == off_idx ? statusVec_3 : _GEN_2; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_4 = 6'h4 == off_idx ? statusVec_4 : _GEN_3; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_5 = 6'h5 == off_idx ? statusVec_5 : _GEN_4; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_6 = 6'h6 == off_idx ? statusVec_6 : _GEN_5; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_7 = 6'h7 == off_idx ? statusVec_7 : _GEN_6; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_8 = 6'h8 == off_idx ? statusVec_8 : _GEN_7; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_9 = 6'h9 == off_idx ? statusVec_9 : _GEN_8; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_10 = 6'ha == off_idx ? statusVec_10 : _GEN_9; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_11 = 6'hb == off_idx ? statusVec_11 : _GEN_10; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_12 = 6'hc == off_idx ? statusVec_12 : _GEN_11; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_13 = 6'hd == off_idx ? statusVec_13 : _GEN_12; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_14 = 6'he == off_idx ? statusVec_14 : _GEN_13; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_15 = 6'hf == off_idx ? statusVec_15 : _GEN_14; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_16 = 6'h10 == off_idx ? statusVec_16 : _GEN_15; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_17 = 6'h11 == off_idx ? statusVec_17 : _GEN_16; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_18 = 6'h12 == off_idx ? statusVec_18 : _GEN_17; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_19 = 6'h13 == off_idx ? statusVec_19 : _GEN_18; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_20 = 6'h14 == off_idx ? statusVec_20 : _GEN_19; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_21 = 6'h15 == off_idx ? statusVec_21 : _GEN_20; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_22 = 6'h16 == off_idx ? statusVec_22 : _GEN_21; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_23 = 6'h17 == off_idx ? statusVec_23 : _GEN_22; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_24 = 6'h18 == off_idx ? statusVec_24 : _GEN_23; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_25 = 6'h19 == off_idx ? statusVec_25 : _GEN_24; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_26 = 6'h1a == off_idx ? statusVec_26 : _GEN_25; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_27 = 6'h1b == off_idx ? statusVec_27 : _GEN_26; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_28 = 6'h1c == off_idx ? statusVec_28 : _GEN_27; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_29 = 6'h1d == off_idx ? statusVec_29 : _GEN_28; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_30 = 6'h1e == off_idx ? statusVec_30 : _GEN_29; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_31 = 6'h1f == off_idx ? statusVec_31 : _GEN_30; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_32 = 6'h20 == off_idx ? statusVec_32 : _GEN_31; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_33 = 6'h21 == off_idx ? statusVec_33 : _GEN_32; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_34 = 6'h22 == off_idx ? statusVec_34 : _GEN_33; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_35 = 6'h23 == off_idx ? statusVec_35 : _GEN_34; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_36 = 6'h24 == off_idx ? statusVec_36 : _GEN_35; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_37 = 6'h25 == off_idx ? statusVec_37 : _GEN_36; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_38 = 6'h26 == off_idx ? statusVec_38 : _GEN_37; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_39 = 6'h27 == off_idx ? statusVec_39 : _GEN_38; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_40 = 6'h28 == off_idx ? statusVec_40 : _GEN_39; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_41 = 6'h29 == off_idx ? statusVec_41 : _GEN_40; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_42 = 6'h2a == off_idx ? statusVec_42 : _GEN_41; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_43 = 6'h2b == off_idx ? statusVec_43 : _GEN_42; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_44 = 6'h2c == off_idx ? statusVec_44 : _GEN_43; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_45 = 6'h2d == off_idx ? statusVec_45 : _GEN_44; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_46 = 6'h2e == off_idx ? statusVec_46 : _GEN_45; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_47 = 6'h2f == off_idx ? statusVec_47 : _GEN_46; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_48 = 6'h30 == off_idx ? statusVec_48 : _GEN_47; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_49 = 6'h31 == off_idx ? statusVec_49 : _GEN_48; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_50 = 6'h32 == off_idx ? statusVec_50 : _GEN_49; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_51 = 6'h33 == off_idx ? statusVec_51 : _GEN_50; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_52 = 6'h34 == off_idx ? statusVec_52 : _GEN_51; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_53 = 6'h35 == off_idx ? statusVec_53 : _GEN_52; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_54 = 6'h36 == off_idx ? statusVec_54 : _GEN_53; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_55 = 6'h37 == off_idx ? statusVec_55 : _GEN_54; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_56 = 6'h38 == off_idx ? statusVec_56 : _GEN_55; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_57 = 6'h39 == off_idx ? statusVec_57 : _GEN_56; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_58 = 6'h3a == off_idx ? statusVec_58 : _GEN_57; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_59 = 6'h3b == off_idx ? statusVec_59 : _GEN_58; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_60 = 6'h3c == off_idx ? statusVec_60 : _GEN_59; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_61 = 6'h3d == off_idx ? statusVec_61 : _GEN_60; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_62 = 6'h3e == off_idx ? statusVec_62 : _GEN_61; // @[CaheCore.scala 52:24:@2636.4]
  assign _GEN_67 = 1'h1; // @[CaheCore.scala 54:16:@2637.4]
  assign _GEN_69 = 6'h0 == off_idx ? io_wstatus : statusVec_0; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_70 = 6'h1 == off_idx ? io_wstatus : statusVec_1; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_71 = 6'h2 == off_idx ? io_wstatus : statusVec_2; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_72 = 6'h3 == off_idx ? io_wstatus : statusVec_3; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_73 = 6'h4 == off_idx ? io_wstatus : statusVec_4; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_74 = 6'h5 == off_idx ? io_wstatus : statusVec_5; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_75 = 6'h6 == off_idx ? io_wstatus : statusVec_6; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_76 = 6'h7 == off_idx ? io_wstatus : statusVec_7; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_77 = 6'h8 == off_idx ? io_wstatus : statusVec_8; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_78 = 6'h9 == off_idx ? io_wstatus : statusVec_9; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_79 = 6'ha == off_idx ? io_wstatus : statusVec_10; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_80 = 6'hb == off_idx ? io_wstatus : statusVec_11; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_81 = 6'hc == off_idx ? io_wstatus : statusVec_12; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_82 = 6'hd == off_idx ? io_wstatus : statusVec_13; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_83 = 6'he == off_idx ? io_wstatus : statusVec_14; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_84 = 6'hf == off_idx ? io_wstatus : statusVec_15; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_85 = 6'h10 == off_idx ? io_wstatus : statusVec_16; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_86 = 6'h11 == off_idx ? io_wstatus : statusVec_17; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_87 = 6'h12 == off_idx ? io_wstatus : statusVec_18; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_88 = 6'h13 == off_idx ? io_wstatus : statusVec_19; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_89 = 6'h14 == off_idx ? io_wstatus : statusVec_20; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_90 = 6'h15 == off_idx ? io_wstatus : statusVec_21; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_91 = 6'h16 == off_idx ? io_wstatus : statusVec_22; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_92 = 6'h17 == off_idx ? io_wstatus : statusVec_23; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_93 = 6'h18 == off_idx ? io_wstatus : statusVec_24; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_94 = 6'h19 == off_idx ? io_wstatus : statusVec_25; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_95 = 6'h1a == off_idx ? io_wstatus : statusVec_26; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_96 = 6'h1b == off_idx ? io_wstatus : statusVec_27; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_97 = 6'h1c == off_idx ? io_wstatus : statusVec_28; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_98 = 6'h1d == off_idx ? io_wstatus : statusVec_29; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_99 = 6'h1e == off_idx ? io_wstatus : statusVec_30; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_100 = 6'h1f == off_idx ? io_wstatus : statusVec_31; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_101 = 6'h20 == off_idx ? io_wstatus : statusVec_32; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_102 = 6'h21 == off_idx ? io_wstatus : statusVec_33; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_103 = 6'h22 == off_idx ? io_wstatus : statusVec_34; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_104 = 6'h23 == off_idx ? io_wstatus : statusVec_35; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_105 = 6'h24 == off_idx ? io_wstatus : statusVec_36; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_106 = 6'h25 == off_idx ? io_wstatus : statusVec_37; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_107 = 6'h26 == off_idx ? io_wstatus : statusVec_38; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_108 = 6'h27 == off_idx ? io_wstatus : statusVec_39; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_109 = 6'h28 == off_idx ? io_wstatus : statusVec_40; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_110 = 6'h29 == off_idx ? io_wstatus : statusVec_41; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_111 = 6'h2a == off_idx ? io_wstatus : statusVec_42; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_112 = 6'h2b == off_idx ? io_wstatus : statusVec_43; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_113 = 6'h2c == off_idx ? io_wstatus : statusVec_44; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_114 = 6'h2d == off_idx ? io_wstatus : statusVec_45; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_115 = 6'h2e == off_idx ? io_wstatus : statusVec_46; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_116 = 6'h2f == off_idx ? io_wstatus : statusVec_47; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_117 = 6'h30 == off_idx ? io_wstatus : statusVec_48; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_118 = 6'h31 == off_idx ? io_wstatus : statusVec_49; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_119 = 6'h32 == off_idx ? io_wstatus : statusVec_50; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_120 = 6'h33 == off_idx ? io_wstatus : statusVec_51; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_121 = 6'h34 == off_idx ? io_wstatus : statusVec_52; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_122 = 6'h35 == off_idx ? io_wstatus : statusVec_53; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_123 = 6'h36 == off_idx ? io_wstatus : statusVec_54; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_124 = 6'h37 == off_idx ? io_wstatus : statusVec_55; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_125 = 6'h38 == off_idx ? io_wstatus : statusVec_56; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_126 = 6'h39 == off_idx ? io_wstatus : statusVec_57; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_127 = 6'h3a == off_idx ? io_wstatus : statusVec_58; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_128 = 6'h3b == off_idx ? io_wstatus : statusVec_59; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_129 = 6'h3c == off_idx ? io_wstatus : statusVec_60; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_130 = 6'h3d == off_idx ? io_wstatus : statusVec_61; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_131 = 6'h3e == off_idx ? io_wstatus : statusVec_62; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_132 = 6'h3f == off_idx ? io_wstatus : statusVec_63; // @[CaheCore.scala 55:37:@2643.6]
  assign _GEN_133 = io_wen ? _GEN_69 : statusVec_0; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_134 = io_wen ? _GEN_70 : statusVec_1; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_135 = io_wen ? _GEN_71 : statusVec_2; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_136 = io_wen ? _GEN_72 : statusVec_3; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_137 = io_wen ? _GEN_73 : statusVec_4; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_138 = io_wen ? _GEN_74 : statusVec_5; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_139 = io_wen ? _GEN_75 : statusVec_6; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_140 = io_wen ? _GEN_76 : statusVec_7; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_141 = io_wen ? _GEN_77 : statusVec_8; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_142 = io_wen ? _GEN_78 : statusVec_9; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_143 = io_wen ? _GEN_79 : statusVec_10; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_144 = io_wen ? _GEN_80 : statusVec_11; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_145 = io_wen ? _GEN_81 : statusVec_12; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_146 = io_wen ? _GEN_82 : statusVec_13; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_147 = io_wen ? _GEN_83 : statusVec_14; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_148 = io_wen ? _GEN_84 : statusVec_15; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_149 = io_wen ? _GEN_85 : statusVec_16; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_150 = io_wen ? _GEN_86 : statusVec_17; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_151 = io_wen ? _GEN_87 : statusVec_18; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_152 = io_wen ? _GEN_88 : statusVec_19; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_153 = io_wen ? _GEN_89 : statusVec_20; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_154 = io_wen ? _GEN_90 : statusVec_21; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_155 = io_wen ? _GEN_91 : statusVec_22; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_156 = io_wen ? _GEN_92 : statusVec_23; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_157 = io_wen ? _GEN_93 : statusVec_24; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_158 = io_wen ? _GEN_94 : statusVec_25; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_159 = io_wen ? _GEN_95 : statusVec_26; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_160 = io_wen ? _GEN_96 : statusVec_27; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_161 = io_wen ? _GEN_97 : statusVec_28; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_162 = io_wen ? _GEN_98 : statusVec_29; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_163 = io_wen ? _GEN_99 : statusVec_30; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_164 = io_wen ? _GEN_100 : statusVec_31; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_165 = io_wen ? _GEN_101 : statusVec_32; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_166 = io_wen ? _GEN_102 : statusVec_33; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_167 = io_wen ? _GEN_103 : statusVec_34; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_168 = io_wen ? _GEN_104 : statusVec_35; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_169 = io_wen ? _GEN_105 : statusVec_36; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_170 = io_wen ? _GEN_106 : statusVec_37; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_171 = io_wen ? _GEN_107 : statusVec_38; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_172 = io_wen ? _GEN_108 : statusVec_39; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_173 = io_wen ? _GEN_109 : statusVec_40; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_174 = io_wen ? _GEN_110 : statusVec_41; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_175 = io_wen ? _GEN_111 : statusVec_42; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_176 = io_wen ? _GEN_112 : statusVec_43; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_177 = io_wen ? _GEN_113 : statusVec_44; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_178 = io_wen ? _GEN_114 : statusVec_45; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_179 = io_wen ? _GEN_115 : statusVec_46; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_180 = io_wen ? _GEN_116 : statusVec_47; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_181 = io_wen ? _GEN_117 : statusVec_48; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_182 = io_wen ? _GEN_118 : statusVec_49; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_183 = io_wen ? _GEN_119 : statusVec_50; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_184 = io_wen ? _GEN_120 : statusVec_51; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_185 = io_wen ? _GEN_121 : statusVec_52; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_186 = io_wen ? _GEN_122 : statusVec_53; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_187 = io_wen ? _GEN_123 : statusVec_54; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_188 = io_wen ? _GEN_124 : statusVec_55; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_189 = io_wen ? _GEN_125 : statusVec_56; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_190 = io_wen ? _GEN_126 : statusVec_57; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_191 = io_wen ? _GEN_127 : statusVec_58; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_192 = io_wen ? _GEN_128 : statusVec_59; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_193 = io_wen ? _GEN_129 : statusVec_60; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_194 = io_wen ? _GEN_130 : statusVec_61; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_195 = io_wen ? _GEN_131 : statusVec_62; // @[CaheCore.scala 55:16:@2642.4]
  assign _GEN_196 = io_wen ? _GEN_132 : statusVec_63; // @[CaheCore.scala 55:16:@2642.4]
  assign rdata_0 = MyMem_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2573.4]
  assign rdata_1 = MyMem_1_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2577.4]
  assign _GEN_198 = 4'h1 == line_idx ? rdata_1 : rdata_0; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_2 = MyMem_2_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2581.4]
  assign _GEN_199 = 4'h2 == line_idx ? rdata_2 : _GEN_198; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_3 = MyMem_3_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2585.4]
  assign _GEN_200 = 4'h3 == line_idx ? rdata_3 : _GEN_199; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_4 = MyMem_4_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2589.4]
  assign _GEN_201 = 4'h4 == line_idx ? rdata_4 : _GEN_200; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_5 = MyMem_5_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2593.4]
  assign _GEN_202 = 4'h5 == line_idx ? rdata_5 : _GEN_201; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_6 = MyMem_6_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2597.4]
  assign _GEN_203 = 4'h6 == line_idx ? rdata_6 : _GEN_202; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_7 = MyMem_7_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2601.4]
  assign _GEN_204 = 4'h7 == line_idx ? rdata_7 : _GEN_203; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_8 = MyMem_8_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2605.4]
  assign _GEN_205 = 4'h8 == line_idx ? rdata_8 : _GEN_204; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_9 = MyMem_9_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2609.4]
  assign _GEN_206 = 4'h9 == line_idx ? rdata_9 : _GEN_205; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_10 = MyMem_10_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2613.4]
  assign _GEN_207 = 4'ha == line_idx ? rdata_10 : _GEN_206; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_11 = MyMem_11_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2617.4]
  assign _GEN_208 = 4'hb == line_idx ? rdata_11 : _GEN_207; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_12 = MyMem_12_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2621.4]
  assign _GEN_209 = 4'hc == line_idx ? rdata_12 : _GEN_208; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_13 = MyMem_13_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2625.4]
  assign _GEN_210 = 4'hd == line_idx ? rdata_13 : _GEN_209; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_14 = MyMem_14_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2629.4]
  assign _GEN_211 = 4'he == line_idx ? rdata_14 : _GEN_210; // @[CaheCore.scala 58:13:@2649.4]
  assign rdata_15 = MyMem_15_io_rdata; // @[CaheCore.scala 42:19:@2569.4 CaheCore.scala 48:14:@2633.4]
  assign _T_560 = tag_RAM_rtag_data == tag; // @[CaheCore.scala 59:21:@2650.4]
  assign io_rdata = 4'hf == line_idx ? rdata_15 : _GEN_211; // @[CaheCore.scala 58:13:@2649.4]
  assign io_rvalid = _T_560 & rstatus; // @[CaheCore.scala 59:13:@2652.4]
  assign MyMem_clock = clock; // @[:@2450.4]
  assign MyMem_io_wen = io_wen; // @[CaheCore.scala 46:24:@2571.4]
  assign MyMem_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2570.4]
  assign MyMem_io_wdata = io_wdata_0; // @[CaheCore.scala 47:24:@2572.4]
  assign MyMem_1_clock = clock; // @[:@2453.4]
  assign MyMem_1_io_wen = io_wen; // @[CaheCore.scala 46:24:@2575.4]
  assign MyMem_1_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2574.4]
  assign MyMem_1_io_wdata = io_wdata_1; // @[CaheCore.scala 47:24:@2576.4]
  assign MyMem_2_clock = clock; // @[:@2456.4]
  assign MyMem_2_io_wen = io_wen; // @[CaheCore.scala 46:24:@2579.4]
  assign MyMem_2_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2578.4]
  assign MyMem_2_io_wdata = io_wdata_2; // @[CaheCore.scala 47:24:@2580.4]
  assign MyMem_3_clock = clock; // @[:@2459.4]
  assign MyMem_3_io_wen = io_wen; // @[CaheCore.scala 46:24:@2583.4]
  assign MyMem_3_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2582.4]
  assign MyMem_3_io_wdata = io_wdata_3; // @[CaheCore.scala 47:24:@2584.4]
  assign MyMem_4_clock = clock; // @[:@2462.4]
  assign MyMem_4_io_wen = io_wen; // @[CaheCore.scala 46:24:@2587.4]
  assign MyMem_4_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2586.4]
  assign MyMem_4_io_wdata = io_wdata_4; // @[CaheCore.scala 47:24:@2588.4]
  assign MyMem_5_clock = clock; // @[:@2465.4]
  assign MyMem_5_io_wen = io_wen; // @[CaheCore.scala 46:24:@2591.4]
  assign MyMem_5_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2590.4]
  assign MyMem_5_io_wdata = io_wdata_5; // @[CaheCore.scala 47:24:@2592.4]
  assign MyMem_6_clock = clock; // @[:@2468.4]
  assign MyMem_6_io_wen = io_wen; // @[CaheCore.scala 46:24:@2595.4]
  assign MyMem_6_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2594.4]
  assign MyMem_6_io_wdata = io_wdata_6; // @[CaheCore.scala 47:24:@2596.4]
  assign MyMem_7_clock = clock; // @[:@2471.4]
  assign MyMem_7_io_wen = io_wen; // @[CaheCore.scala 46:24:@2599.4]
  assign MyMem_7_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2598.4]
  assign MyMem_7_io_wdata = io_wdata_7; // @[CaheCore.scala 47:24:@2600.4]
  assign MyMem_8_clock = clock; // @[:@2474.4]
  assign MyMem_8_io_wen = io_wen; // @[CaheCore.scala 46:24:@2603.4]
  assign MyMem_8_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2602.4]
  assign MyMem_8_io_wdata = io_wdata_8; // @[CaheCore.scala 47:24:@2604.4]
  assign MyMem_9_clock = clock; // @[:@2477.4]
  assign MyMem_9_io_wen = io_wen; // @[CaheCore.scala 46:24:@2607.4]
  assign MyMem_9_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2606.4]
  assign MyMem_9_io_wdata = io_wdata_9; // @[CaheCore.scala 47:24:@2608.4]
  assign MyMem_10_clock = clock; // @[:@2480.4]
  assign MyMem_10_io_wen = io_wen; // @[CaheCore.scala 46:24:@2611.4]
  assign MyMem_10_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2610.4]
  assign MyMem_10_io_wdata = io_wdata_10; // @[CaheCore.scala 47:24:@2612.4]
  assign MyMem_11_clock = clock; // @[:@2483.4]
  assign MyMem_11_io_wen = io_wen; // @[CaheCore.scala 46:24:@2615.4]
  assign MyMem_11_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2614.4]
  assign MyMem_11_io_wdata = io_wdata_11; // @[CaheCore.scala 47:24:@2616.4]
  assign MyMem_12_clock = clock; // @[:@2486.4]
  assign MyMem_12_io_wen = io_wen; // @[CaheCore.scala 46:24:@2619.4]
  assign MyMem_12_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2618.4]
  assign MyMem_12_io_wdata = io_wdata_12; // @[CaheCore.scala 47:24:@2620.4]
  assign MyMem_13_clock = clock; // @[:@2489.4]
  assign MyMem_13_io_wen = io_wen; // @[CaheCore.scala 46:24:@2623.4]
  assign MyMem_13_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2622.4]
  assign MyMem_13_io_wdata = io_wdata_13; // @[CaheCore.scala 47:24:@2624.4]
  assign MyMem_14_clock = clock; // @[:@2492.4]
  assign MyMem_14_io_wen = io_wen; // @[CaheCore.scala 46:24:@2627.4]
  assign MyMem_14_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2626.4]
  assign MyMem_14_io_wdata = io_wdata_14; // @[CaheCore.scala 47:24:@2628.4]
  assign MyMem_15_clock = clock; // @[:@2495.4]
  assign MyMem_15_io_wen = io_wen; // @[CaheCore.scala 46:24:@2631.4]
  assign MyMem_15_io_addr = io_addr[11:6]; // @[CaheCore.scala 45:24:@2630.4]
  assign MyMem_15_io_wdata = io_wdata_15; // @[CaheCore.scala 47:24:@2632.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 64; initvar = initvar+1)
    tag_RAM[initvar] = _RAND_0[19:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  statusVec_0 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  statusVec_1 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  statusVec_2 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  statusVec_3 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  statusVec_4 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  statusVec_5 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  statusVec_6 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  statusVec_7 = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  statusVec_8 = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  statusVec_9 = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  statusVec_10 = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  statusVec_11 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  statusVec_12 = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  statusVec_13 = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  statusVec_14 = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  statusVec_15 = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  statusVec_16 = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  statusVec_17 = _RAND_18[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  statusVec_18 = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  statusVec_19 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  statusVec_20 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  statusVec_21 = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  statusVec_22 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  statusVec_23 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  statusVec_24 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  statusVec_25 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  statusVec_26 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  statusVec_27 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  statusVec_28 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  statusVec_29 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  statusVec_30 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  statusVec_31 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  statusVec_32 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  statusVec_33 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  statusVec_34 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  statusVec_35 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  statusVec_36 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  statusVec_37 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  statusVec_38 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  statusVec_39 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  statusVec_40 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  statusVec_41 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  statusVec_42 = _RAND_43[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  statusVec_43 = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  statusVec_44 = _RAND_45[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  statusVec_45 = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  statusVec_46 = _RAND_47[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  statusVec_47 = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  statusVec_48 = _RAND_49[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  statusVec_49 = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  statusVec_50 = _RAND_51[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  statusVec_51 = _RAND_52[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  statusVec_52 = _RAND_53[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  statusVec_53 = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  statusVec_54 = _RAND_55[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  statusVec_55 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  statusVec_56 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  statusVec_57 = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  statusVec_58 = _RAND_59[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  statusVec_59 = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  statusVec_60 = _RAND_61[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  statusVec_61 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  statusVec_62 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  statusVec_63 = _RAND_64[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  line_idx = _RAND_65[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  rstatus = _RAND_66[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  tag = _RAND_67[19:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  tag_RAM_rtag_addr_pipe_0 = _RAND_68[5:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(tag_RAM__T_550_en & tag_RAM__T_550_mask) begin
      tag_RAM[tag_RAM__T_550_addr] <= tag_RAM__T_550_data; // @[CaheCore.scala 35:30:@2497.4]
    end
    if (reset) begin
      statusVec_0 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h0 == off_idx) begin
          statusVec_0 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_1 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1 == off_idx) begin
          statusVec_1 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_2 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2 == off_idx) begin
          statusVec_2 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_3 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3 == off_idx) begin
          statusVec_3 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_4 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h4 == off_idx) begin
          statusVec_4 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_5 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h5 == off_idx) begin
          statusVec_5 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_6 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h6 == off_idx) begin
          statusVec_6 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_7 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h7 == off_idx) begin
          statusVec_7 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_8 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h8 == off_idx) begin
          statusVec_8 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_9 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h9 == off_idx) begin
          statusVec_9 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_10 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'ha == off_idx) begin
          statusVec_10 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_11 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hb == off_idx) begin
          statusVec_11 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_12 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hc == off_idx) begin
          statusVec_12 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_13 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hd == off_idx) begin
          statusVec_13 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_14 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'he == off_idx) begin
          statusVec_14 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_15 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'hf == off_idx) begin
          statusVec_15 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_16 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h10 == off_idx) begin
          statusVec_16 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_17 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h11 == off_idx) begin
          statusVec_17 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_18 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h12 == off_idx) begin
          statusVec_18 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_19 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h13 == off_idx) begin
          statusVec_19 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_20 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h14 == off_idx) begin
          statusVec_20 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_21 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h15 == off_idx) begin
          statusVec_21 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_22 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h16 == off_idx) begin
          statusVec_22 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_23 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h17 == off_idx) begin
          statusVec_23 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_24 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h18 == off_idx) begin
          statusVec_24 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_25 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h19 == off_idx) begin
          statusVec_25 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_26 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1a == off_idx) begin
          statusVec_26 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_27 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1b == off_idx) begin
          statusVec_27 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_28 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1c == off_idx) begin
          statusVec_28 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_29 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1d == off_idx) begin
          statusVec_29 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_30 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1e == off_idx) begin
          statusVec_30 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_31 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h1f == off_idx) begin
          statusVec_31 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_32 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h20 == off_idx) begin
          statusVec_32 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_33 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h21 == off_idx) begin
          statusVec_33 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_34 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h22 == off_idx) begin
          statusVec_34 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_35 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h23 == off_idx) begin
          statusVec_35 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_36 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h24 == off_idx) begin
          statusVec_36 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_37 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h25 == off_idx) begin
          statusVec_37 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_38 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h26 == off_idx) begin
          statusVec_38 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_39 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h27 == off_idx) begin
          statusVec_39 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_40 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h28 == off_idx) begin
          statusVec_40 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_41 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h29 == off_idx) begin
          statusVec_41 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_42 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2a == off_idx) begin
          statusVec_42 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_43 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2b == off_idx) begin
          statusVec_43 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_44 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2c == off_idx) begin
          statusVec_44 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_45 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2d == off_idx) begin
          statusVec_45 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_46 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2e == off_idx) begin
          statusVec_46 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_47 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h2f == off_idx) begin
          statusVec_47 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_48 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h30 == off_idx) begin
          statusVec_48 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_49 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h31 == off_idx) begin
          statusVec_49 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_50 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h32 == off_idx) begin
          statusVec_50 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_51 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h33 == off_idx) begin
          statusVec_51 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_52 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h34 == off_idx) begin
          statusVec_52 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_53 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h35 == off_idx) begin
          statusVec_53 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_54 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h36 == off_idx) begin
          statusVec_54 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_55 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h37 == off_idx) begin
          statusVec_55 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_56 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h38 == off_idx) begin
          statusVec_56 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_57 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h39 == off_idx) begin
          statusVec_57 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_58 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3a == off_idx) begin
          statusVec_58 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_59 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3b == off_idx) begin
          statusVec_59 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_60 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3c == off_idx) begin
          statusVec_60 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_61 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3d == off_idx) begin
          statusVec_61 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_62 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3e == off_idx) begin
          statusVec_62 <= io_wstatus;
        end
      end
    end
    if (reset) begin
      statusVec_63 <= 1'h0;
    end else begin
      if (io_wen) begin
        if (6'h3f == off_idx) begin
          statusVec_63 <= io_wstatus;
        end
      end
    end
    line_idx <= io_addr[5:2];
    if (6'h3f == off_idx) begin
      rstatus <= statusVec_63;
    end else begin
      if (6'h3e == off_idx) begin
        rstatus <= statusVec_62;
      end else begin
        if (6'h3d == off_idx) begin
          rstatus <= statusVec_61;
        end else begin
          if (6'h3c == off_idx) begin
            rstatus <= statusVec_60;
          end else begin
            if (6'h3b == off_idx) begin
              rstatus <= statusVec_59;
            end else begin
              if (6'h3a == off_idx) begin
                rstatus <= statusVec_58;
              end else begin
                if (6'h39 == off_idx) begin
                  rstatus <= statusVec_57;
                end else begin
                  if (6'h38 == off_idx) begin
                    rstatus <= statusVec_56;
                  end else begin
                    if (6'h37 == off_idx) begin
                      rstatus <= statusVec_55;
                    end else begin
                      if (6'h36 == off_idx) begin
                        rstatus <= statusVec_54;
                      end else begin
                        if (6'h35 == off_idx) begin
                          rstatus <= statusVec_53;
                        end else begin
                          if (6'h34 == off_idx) begin
                            rstatus <= statusVec_52;
                          end else begin
                            if (6'h33 == off_idx) begin
                              rstatus <= statusVec_51;
                            end else begin
                              if (6'h32 == off_idx) begin
                                rstatus <= statusVec_50;
                              end else begin
                                if (6'h31 == off_idx) begin
                                  rstatus <= statusVec_49;
                                end else begin
                                  if (6'h30 == off_idx) begin
                                    rstatus <= statusVec_48;
                                  end else begin
                                    if (6'h2f == off_idx) begin
                                      rstatus <= statusVec_47;
                                    end else begin
                                      if (6'h2e == off_idx) begin
                                        rstatus <= statusVec_46;
                                      end else begin
                                        if (6'h2d == off_idx) begin
                                          rstatus <= statusVec_45;
                                        end else begin
                                          if (6'h2c == off_idx) begin
                                            rstatus <= statusVec_44;
                                          end else begin
                                            if (6'h2b == off_idx) begin
                                              rstatus <= statusVec_43;
                                            end else begin
                                              if (6'h2a == off_idx) begin
                                                rstatus <= statusVec_42;
                                              end else begin
                                                if (6'h29 == off_idx) begin
                                                  rstatus <= statusVec_41;
                                                end else begin
                                                  if (6'h28 == off_idx) begin
                                                    rstatus <= statusVec_40;
                                                  end else begin
                                                    if (6'h27 == off_idx) begin
                                                      rstatus <= statusVec_39;
                                                    end else begin
                                                      if (6'h26 == off_idx) begin
                                                        rstatus <= statusVec_38;
                                                      end else begin
                                                        if (6'h25 == off_idx) begin
                                                          rstatus <= statusVec_37;
                                                        end else begin
                                                          if (6'h24 == off_idx) begin
                                                            rstatus <= statusVec_36;
                                                          end else begin
                                                            if (6'h23 == off_idx) begin
                                                              rstatus <= statusVec_35;
                                                            end else begin
                                                              if (6'h22 == off_idx) begin
                                                                rstatus <= statusVec_34;
                                                              end else begin
                                                                if (6'h21 == off_idx) begin
                                                                  rstatus <= statusVec_33;
                                                                end else begin
                                                                  if (6'h20 == off_idx) begin
                                                                    rstatus <= statusVec_32;
                                                                  end else begin
                                                                    if (6'h1f == off_idx) begin
                                                                      rstatus <= statusVec_31;
                                                                    end else begin
                                                                      if (6'h1e == off_idx) begin
                                                                        rstatus <= statusVec_30;
                                                                      end else begin
                                                                        if (6'h1d == off_idx) begin
                                                                          rstatus <= statusVec_29;
                                                                        end else begin
                                                                          if (6'h1c == off_idx) begin
                                                                            rstatus <= statusVec_28;
                                                                          end else begin
                                                                            if (6'h1b == off_idx) begin
                                                                              rstatus <= statusVec_27;
                                                                            end else begin
                                                                              if (6'h1a == off_idx) begin
                                                                                rstatus <= statusVec_26;
                                                                              end else begin
                                                                                if (6'h19 == off_idx) begin
                                                                                  rstatus <= statusVec_25;
                                                                                end else begin
                                                                                  if (6'h18 == off_idx) begin
                                                                                    rstatus <= statusVec_24;
                                                                                  end else begin
                                                                                    if (6'h17 == off_idx) begin
                                                                                      rstatus <= statusVec_23;
                                                                                    end else begin
                                                                                      if (6'h16 == off_idx) begin
                                                                                        rstatus <= statusVec_22;
                                                                                      end else begin
                                                                                        if (6'h15 == off_idx) begin
                                                                                          rstatus <= statusVec_21;
                                                                                        end else begin
                                                                                          if (6'h14 == off_idx) begin
                                                                                            rstatus <= statusVec_20;
                                                                                          end else begin
                                                                                            if (6'h13 == off_idx) begin
                                                                                              rstatus <= statusVec_19;
                                                                                            end else begin
                                                                                              if (6'h12 == off_idx) begin
                                                                                                rstatus <= statusVec_18;
                                                                                              end else begin
                                                                                                if (6'h11 == off_idx) begin
                                                                                                  rstatus <= statusVec_17;
                                                                                                end else begin
                                                                                                  if (6'h10 == off_idx) begin
                                                                                                    rstatus <= statusVec_16;
                                                                                                  end else begin
                                                                                                    if (6'hf == off_idx) begin
                                                                                                      rstatus <= statusVec_15;
                                                                                                    end else begin
                                                                                                      if (6'he == off_idx) begin
                                                                                                        rstatus <= statusVec_14;
                                                                                                      end else begin
                                                                                                        if (6'hd == off_idx) begin
                                                                                                          rstatus <= statusVec_13;
                                                                                                        end else begin
                                                                                                          if (6'hc == off_idx) begin
                                                                                                            rstatus <= statusVec_12;
                                                                                                          end else begin
                                                                                                            if (6'hb == off_idx) begin
                                                                                                              rstatus <= statusVec_11;
                                                                                                            end else begin
                                                                                                              if (6'ha == off_idx) begin
                                                                                                                rstatus <= statusVec_10;
                                                                                                              end else begin
                                                                                                                if (6'h9 == off_idx) begin
                                                                                                                  rstatus <= statusVec_9;
                                                                                                                end else begin
                                                                                                                  if (6'h8 == off_idx) begin
                                                                                                                    rstatus <= statusVec_8;
                                                                                                                  end else begin
                                                                                                                    if (6'h7 == off_idx) begin
                                                                                                                      rstatus <= statusVec_7;
                                                                                                                    end else begin
                                                                                                                      if (6'h6 == off_idx) begin
                                                                                                                        rstatus <= statusVec_6;
                                                                                                                      end else begin
                                                                                                                        if (6'h5 == off_idx) begin
                                                                                                                          rstatus <= statusVec_5;
                                                                                                                        end else begin
                                                                                                                          if (6'h4 == off_idx) begin
                                                                                                                            rstatus <= statusVec_4;
                                                                                                                          end else begin
                                                                                                                            if (6'h3 == off_idx) begin
                                                                                                                              rstatus <= statusVec_3;
                                                                                                                            end else begin
                                                                                                                              if (6'h2 == off_idx) begin
                                                                                                                                rstatus <= statusVec_2;
                                                                                                                              end else begin
                                                                                                                                if (6'h1 == off_idx) begin
                                                                                                                                  rstatus <= statusVec_1;
                                                                                                                                end else begin
                                                                                                                                  rstatus <= statusVec_0;
                                                                                                                                end
                                                                                                                              end
                                                                                                                            end
                                                                                                                          end
                                                                                                                        end
                                                                                                                      end
                                                                                                                    end
                                                                                                                  end
                                                                                                                end
                                                                                                              end
                                                                                                            end
                                                                                                          end
                                                                                                        end
                                                                                                      end
                                                                                                    end
                                                                                                  end
                                                                                                end
                                                                                              end
                                                                                            end
                                                                                          end
                                                                                        end
                                                                                      end
                                                                                    end
                                                                                  end
                                                                                end
                                                                              end
                                                                            end
                                                                          end
                                                                        end
                                                                      end
                                                                    end
                                                                  end
                                                                end
                                                              end
                                                            end
                                                          end
                                                        end
                                                      end
                                                    end
                                                  end
                                                end
                                              end
                                            end
                                          end
                                        end
                                      end
                                    end
                                  end
                                end
                              end
                            end
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    tag <= io_addr[31:12];
    if (_GEN_67) begin
      tag_RAM_rtag_addr_pipe_0 <= off_idx;
    end
  end
endmodule
module Icache( // @[:@2654.2]
  input         clock, // @[:@2655.4]
  input         reset, // @[:@2656.4]
  input         io_core_pc_valid, // @[:@2657.4]
  input  [31:0] io_core_pc_bits, // @[:@2657.4]
  output        io_core_inst_valid, // @[:@2657.4]
  output [31:0] io_core_inst_bits, // @[:@2657.4]
  output        io_core_ready, // @[:@2657.4]
  input  [31:0] io_axi_r_data, // @[:@2657.4]
  input         io_axi_r_valid, // @[:@2657.4]
  input         io_axi_r_last, // @[:@2657.4]
  input         io_axi_ar_ready, // @[:@2657.4]
  output        io_axi_ar_valid, // @[:@2657.4]
  output [31:0] io_axi_ar_addr // @[:@2657.4]
);
  wire  icache_clock; // @[Icache.scala 66:22:@2677.4]
  wire  icache_reset; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_wen; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_addr; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_0; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_1; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_2; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_3; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_4; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_5; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_6; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_7; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_8; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_9; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_10; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_11; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_12; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_13; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_14; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_wdata_15; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_wstatus; // @[Icache.scala 66:22:@2677.4]
  wire [31:0] icache_io_rdata; // @[Icache.scala 66:22:@2677.4]
  wire  icache_io_rvalid; // @[Icache.scala 66:22:@2677.4]
  reg  pc_valid; // @[Icache.scala 56:25:@2667.4]
  reg [31:0] _RAND_0;
  reg [31:0] pc; // @[Icache.scala 57:15:@2668.4]
  reg [31:0] _RAND_1;
  wire  pc_accept; // @[Icache.scala 58:39:@2669.4]
  reg [1:0] state; // @[Icache.scala 62:22:@2674.4]
  reg [31:0] _RAND_2;
  reg [31:0] wb_buffer_0; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_3;
  reg [31:0] wb_buffer_1; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_4;
  reg [31:0] wb_buffer_2; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_5;
  reg [31:0] wb_buffer_3; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_6;
  reg [31:0] wb_buffer_4; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_7;
  reg [31:0] wb_buffer_5; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_8;
  reg [31:0] wb_buffer_6; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_9;
  reg [31:0] wb_buffer_7; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_10;
  reg [31:0] wb_buffer_8; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_11;
  reg [31:0] wb_buffer_9; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_12;
  reg [31:0] wb_buffer_10; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_13;
  reg [31:0] wb_buffer_11; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_14;
  reg [31:0] wb_buffer_12; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_15;
  reg [31:0] wb_buffer_13; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_16;
  reg [31:0] wb_buffer_14; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_17;
  reg [31:0] wb_buffer_15; // @[Icache.scala 64:22:@2675.4]
  reg [31:0] _RAND_18;
  reg [25:0] wb_addr; // @[Icache.scala 65:20:@2676.4]
  reg [31:0] _RAND_19;
  wire  _T_78; // @[Icache.scala 67:30:@2680.4]
  wire [31:0] _T_81; // @[Cat.scala 30:58:@2683.4]
  wire  cache_hit; // @[Icache.scala 73:33:@2705.4]
  wire [25:0] _T_84; // @[Icache.scala 74:26:@2706.4]
  wire  line_hit; // @[Icache.scala 74:59:@2707.4]
  wire  _T_86; // @[Icache.scala 75:36:@2708.4]
  wire  miss; // @[Icache.scala 75:33:@2709.4]
  wire  _T_87; // @[Icache.scala 76:39:@2710.4]
  wire  _T_89; // @[Icache.scala 76:54:@2711.4]
  wire  _T_90; // @[Icache.scala 76:51:@2712.4]
  wire  pc_miss; // @[Icache.scala 76:29:@2713.4]
  wire  _T_91; // @[Icache.scala 79:50:@2714.4]
  wire  _T_92; // @[Icache.scala 79:41:@2715.4]
  wire  _T_95; // @[Icache.scala 79:62:@2717.4]
  reg  _T_99; // @[Icache.scala 27:27:@2719.4]
  reg [31:0] _RAND_20;
  wire  _GEN_1; // @[Icache.scala 29:20:@2724.6]
  wire  _GEN_2; // @[Icache.scala 28:17:@2720.4]
  wire  pc_double_miss; // @[Icache.scala 30:8:@2727.4]
  reg  _T_104; // @[Icache.scala 27:27:@2728.4]
  reg [31:0] _RAND_21;
  wire  _GEN_3; // @[Icache.scala 29:20:@2733.6]
  wire  _GEN_4; // @[Icache.scala 28:17:@2729.4]
  wire  _T_112; // @[Conditional.scala 37:30:@2743.4]
  wire [1:0] _GEN_5; // @[Icache.scala 86:22:@2745.6]
  wire  _T_113; // @[Conditional.scala 37:30:@2753.6]
  wire  _T_114; // @[Icache.scala 90:19:@2755.8]
  wire [1:0] _GEN_6; // @[Icache.scala 90:30:@2756.8]
  wire  _T_115; // @[Conditional.scala 37:30:@2764.8]
  wire [1:0] _GEN_7; // @[Icache.scala 94:29:@2766.10]
  wire [1:0] _GEN_8; // @[Conditional.scala 39:67:@2765.8]
  wire [1:0] _GEN_9; // @[Conditional.scala 39:67:@2754.6]
  wire [1:0] _GEN_10; // @[Conditional.scala 40:58:@2744.4]
  wire  _T_117; // @[Icache.scala 99:31:@2774.4]
  wire  _T_119; // @[Icache.scala 100:31:@2776.4]
  wire  _T_120; // @[Icache.scala 99:43:@2777.4]
  reg [3:0] cnt; // @[Icache.scala 103:20:@2782.4]
  reg [31:0] _RAND_22;
  reg  wb_buf_valid_0; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_23;
  reg  wb_buf_valid_1; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_24;
  reg  wb_buf_valid_2; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_25;
  reg  wb_buf_valid_3; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_26;
  reg  wb_buf_valid_4; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_27;
  reg  wb_buf_valid_5; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_28;
  reg  wb_buf_valid_6; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_29;
  reg  wb_buf_valid_7; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_30;
  reg  wb_buf_valid_8; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_31;
  reg  wb_buf_valid_9; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_32;
  reg  wb_buf_valid_10; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_33;
  reg  wb_buf_valid_11; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_34;
  reg  wb_buf_valid_12; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_35;
  reg  wb_buf_valid_13; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_36;
  reg  wb_buf_valid_14; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_37;
  reg  wb_buf_valid_15; // @[Icache.scala 104:29:@2800.4]
  reg [31:0] _RAND_38;
  wire [4:0] _T_268; // @[Icache.scala 110:18:@2820.8]
  wire [3:0] _T_269; // @[Icache.scala 110:18:@2821.8]
  wire  _GEN_12; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_13; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_14; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_15; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_16; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_17; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_18; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_19; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_20; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_21; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_22; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_23; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_24; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_25; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_26; // @[Icache.scala 111:25:@2823.8]
  wire  _GEN_27; // @[Icache.scala 111:25:@2823.8]
  wire [3:0] _GEN_28; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_29; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_30; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_31; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_32; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_33; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_34; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_35; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_36; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_37; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_38; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_39; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_40; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_41; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_42; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_43; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_44; // @[Icache.scala 109:19:@2819.6]
  wire  _GEN_45; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_46; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_47; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_48; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_49; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_50; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_51; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_52; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_53; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_54; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_55; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_56; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_57; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_58; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_59; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_60; // @[Icache.scala 115:23:@2831.8]
  wire  _GEN_62; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_63; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_64; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_65; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_66; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_67; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_68; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_69; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_70; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_71; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_72; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_73; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_74; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_75; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_76; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_77; // @[Icache.scala 113:22:@2827.6]
  wire  _GEN_78; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_79; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_80; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_81; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_82; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_83; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_84; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_85; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_86; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_87; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_88; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_89; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_90; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_91; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_92; // @[Icache.scala 105:31:@2802.4]
  wire  _GEN_93; // @[Icache.scala 105:31:@2802.4]
  wire [3:0] _GEN_94; // @[Icache.scala 105:31:@2802.4]
  wire [31:0] _GEN_95; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_96; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_97; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_98; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_99; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_100; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_101; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_102; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_103; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_104; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_105; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_106; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_107; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_108; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_109; // @[Icache.scala 118:34:@2834.6]
  wire [31:0] _GEN_110; // @[Icache.scala 118:34:@2834.6]
  wire  _T_283; // @[Icache.scala 121:27:@2837.4]
  wire  _T_284; // @[Icache.scala 121:39:@2838.4]
  wire  _T_287; // @[Icache.scala 121:52:@2841.4]
  wire  wait_inst_back; // @[Icache.scala 122:39:@2844.4]
  wire [3:0] line_idx; // @[Icache.scala 125:23:@2845.4]
  wire [31:0] _GEN_128; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_129; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_130; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_131; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_132; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_133; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_134; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_135; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_136; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_137; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_138; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_139; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_140; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_141; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] _GEN_142; // @[Icache.scala 126:24:@2846.4]
  wire [31:0] buffer_inst; // @[Icache.scala 126:24:@2846.4]
  wire  _GEN_144; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_145; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_146; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_147; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_148; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_149; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_150; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_151; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_152; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_153; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_154; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_155; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_156; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_157; // @[Icache.scala 127:78:@2847.4]
  wire  _GEN_158; // @[Icache.scala 127:78:@2847.4]
  wire  _T_294; // @[Icache.scala 127:78:@2847.4]
  reg  _T_297; // @[Icache.scala 36:27:@2848.4]
  reg [31:0] _RAND_39;
  wire  _GEN_159; // @[Icache.scala 38:20:@2853.6]
  wire  _GEN_160; // @[Icache.scala 37:17:@2849.4]
  wire  _T_300; // @[Icache.scala 39:9:@2856.4]
  wire  _T_301; // @[Icache.scala 39:22:@2857.4]
  wire  buf_inst_valid; // @[Icache.scala 127:91:@2858.4]
  CaheCore icache ( // @[Icache.scala 66:22:@2677.4]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_wen(icache_io_wen),
    .io_addr(icache_io_addr),
    .io_wdata_0(icache_io_wdata_0),
    .io_wdata_1(icache_io_wdata_1),
    .io_wdata_2(icache_io_wdata_2),
    .io_wdata_3(icache_io_wdata_3),
    .io_wdata_4(icache_io_wdata_4),
    .io_wdata_5(icache_io_wdata_5),
    .io_wdata_6(icache_io_wdata_6),
    .io_wdata_7(icache_io_wdata_7),
    .io_wdata_8(icache_io_wdata_8),
    .io_wdata_9(icache_io_wdata_9),
    .io_wdata_10(icache_io_wdata_10),
    .io_wdata_11(icache_io_wdata_11),
    .io_wdata_12(icache_io_wdata_12),
    .io_wdata_13(icache_io_wdata_13),
    .io_wdata_14(icache_io_wdata_14),
    .io_wdata_15(icache_io_wdata_15),
    .io_wstatus(icache_io_wstatus),
    .io_rdata(icache_io_rdata),
    .io_rvalid(icache_io_rvalid)
  );
  assign pc_accept = io_core_ready & io_core_pc_valid; // @[Icache.scala 58:39:@2669.4]
  assign _T_78 = state == 2'h2; // @[Icache.scala 67:30:@2680.4]
  assign _T_81 = {wb_addr,6'h0}; // @[Cat.scala 30:58:@2683.4]
  assign cache_hit = pc_valid & icache_io_rvalid; // @[Icache.scala 73:33:@2705.4]
  assign _T_84 = pc[31:6]; // @[Icache.scala 74:26:@2706.4]
  assign line_hit = _T_84 == wb_addr; // @[Icache.scala 74:59:@2707.4]
  assign _T_86 = icache_io_rvalid == 1'h0; // @[Icache.scala 75:36:@2708.4]
  assign miss = pc_valid & _T_86; // @[Icache.scala 75:33:@2709.4]
  assign _T_87 = state == 2'h0; // @[Icache.scala 76:39:@2710.4]
  assign _T_89 = line_hit == 1'h0; // @[Icache.scala 76:54:@2711.4]
  assign _T_90 = _T_87 | _T_89; // @[Icache.scala 76:51:@2712.4]
  assign pc_miss = miss & _T_90; // @[Icache.scala 76:29:@2713.4]
  assign _T_91 = state != 2'h0; // @[Icache.scala 79:50:@2714.4]
  assign _T_92 = miss & _T_91; // @[Icache.scala 79:41:@2715.4]
  assign _T_95 = _T_92 & _T_89; // @[Icache.scala 79:62:@2717.4]
  assign _GEN_1 = _T_95 ? 1'h1 : _T_99; // @[Icache.scala 29:20:@2724.6]
  assign _GEN_2 = _T_78 ? 1'h0 : _GEN_1; // @[Icache.scala 28:17:@2720.4]
  assign pc_double_miss = _T_95 | _T_99; // @[Icache.scala 30:8:@2727.4]
  assign _GEN_3 = pc_miss ? 1'h1 : _T_104; // @[Icache.scala 29:20:@2733.6]
  assign _GEN_4 = io_axi_ar_ready ? 1'h0 : _GEN_3; // @[Icache.scala 28:17:@2729.4]
  assign _T_112 = 2'h0 == state; // @[Conditional.scala 37:30:@2743.4]
  assign _GEN_5 = pc_miss ? 2'h1 : 2'h0; // @[Icache.scala 86:22:@2745.6]
  assign _T_113 = 2'h1 == state; // @[Conditional.scala 37:30:@2753.6]
  assign _T_114 = io_axi_r_last & io_axi_r_valid; // @[Icache.scala 90:19:@2755.8]
  assign _GEN_6 = _T_114 ? 2'h2 : 2'h1; // @[Icache.scala 90:30:@2756.8]
  assign _T_115 = 2'h2 == state; // @[Conditional.scala 37:30:@2764.8]
  assign _GEN_7 = pc_double_miss ? 2'h1 : 2'h0; // @[Icache.scala 94:29:@2766.10]
  assign _GEN_8 = _T_115 ? _GEN_7 : state; // @[Conditional.scala 39:67:@2765.8]
  assign _GEN_9 = _T_113 ? _GEN_6 : _GEN_8; // @[Conditional.scala 39:67:@2754.6]
  assign _GEN_10 = _T_112 ? _GEN_5 : _GEN_9; // @[Conditional.scala 40:58:@2744.4]
  assign _T_117 = _T_87 & pc_miss; // @[Icache.scala 99:31:@2774.4]
  assign _T_119 = _T_78 & pc_double_miss; // @[Icache.scala 100:31:@2776.4]
  assign _T_120 = _T_117 | _T_119; // @[Icache.scala 99:43:@2777.4]
  assign _T_268 = cnt + 4'h1; // @[Icache.scala 110:18:@2820.8]
  assign _T_269 = cnt + 4'h1; // @[Icache.scala 110:18:@2821.8]
  assign _GEN_12 = 4'h0 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_13 = 4'h1 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_14 = 4'h2 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_15 = 4'h3 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_16 = 4'h4 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_17 = 4'h5 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_18 = 4'h6 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_19 = 4'h7 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_20 = 4'h8 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_21 = 4'h9 == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_22 = 4'ha == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_23 = 4'hb == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_24 = 4'hc == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_25 = 4'hd == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_26 = 4'he == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_27 = 4'hf == cnt; // @[Icache.scala 111:25:@2823.8]
  assign _GEN_28 = io_axi_r_valid ? _T_269 : cnt; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_29 = io_axi_r_valid ? _GEN_12 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_30 = io_axi_r_valid ? _GEN_13 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_31 = io_axi_r_valid ? _GEN_14 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_32 = io_axi_r_valid ? _GEN_15 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_33 = io_axi_r_valid ? _GEN_16 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_34 = io_axi_r_valid ? _GEN_17 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_35 = io_axi_r_valid ? _GEN_18 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_36 = io_axi_r_valid ? _GEN_19 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_37 = io_axi_r_valid ? _GEN_20 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_38 = io_axi_r_valid ? _GEN_21 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_39 = io_axi_r_valid ? _GEN_22 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_40 = io_axi_r_valid ? _GEN_23 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_41 = io_axi_r_valid ? _GEN_24 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_42 = io_axi_r_valid ? _GEN_25 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_43 = io_axi_r_valid ? _GEN_26 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_44 = io_axi_r_valid ? _GEN_27 : 1'h0; // @[Icache.scala 109:19:@2819.6]
  assign _GEN_45 = 4'h0 == cnt ? 1'h1 : wb_buf_valid_0; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_46 = 4'h1 == cnt ? 1'h1 : wb_buf_valid_1; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_47 = 4'h2 == cnt ? 1'h1 : wb_buf_valid_2; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_48 = 4'h3 == cnt ? 1'h1 : wb_buf_valid_3; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_49 = 4'h4 == cnt ? 1'h1 : wb_buf_valid_4; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_50 = 4'h5 == cnt ? 1'h1 : wb_buf_valid_5; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_51 = 4'h6 == cnt ? 1'h1 : wb_buf_valid_6; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_52 = 4'h7 == cnt ? 1'h1 : wb_buf_valid_7; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_53 = 4'h8 == cnt ? 1'h1 : wb_buf_valid_8; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_54 = 4'h9 == cnt ? 1'h1 : wb_buf_valid_9; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_55 = 4'ha == cnt ? 1'h1 : wb_buf_valid_10; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_56 = 4'hb == cnt ? 1'h1 : wb_buf_valid_11; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_57 = 4'hc == cnt ? 1'h1 : wb_buf_valid_12; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_58 = 4'hd == cnt ? 1'h1 : wb_buf_valid_13; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_59 = 4'he == cnt ? 1'h1 : wb_buf_valid_14; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_60 = 4'hf == cnt ? 1'h1 : wb_buf_valid_15; // @[Icache.scala 115:23:@2831.8]
  assign _GEN_62 = io_axi_r_valid ? _GEN_45 : wb_buf_valid_0; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_63 = io_axi_r_valid ? _GEN_46 : wb_buf_valid_1; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_64 = io_axi_r_valid ? _GEN_47 : wb_buf_valid_2; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_65 = io_axi_r_valid ? _GEN_48 : wb_buf_valid_3; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_66 = io_axi_r_valid ? _GEN_49 : wb_buf_valid_4; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_67 = io_axi_r_valid ? _GEN_50 : wb_buf_valid_5; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_68 = io_axi_r_valid ? _GEN_51 : wb_buf_valid_6; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_69 = io_axi_r_valid ? _GEN_52 : wb_buf_valid_7; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_70 = io_axi_r_valid ? _GEN_53 : wb_buf_valid_8; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_71 = io_axi_r_valid ? _GEN_54 : wb_buf_valid_9; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_72 = io_axi_r_valid ? _GEN_55 : wb_buf_valid_10; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_73 = io_axi_r_valid ? _GEN_56 : wb_buf_valid_11; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_74 = io_axi_r_valid ? _GEN_57 : wb_buf_valid_12; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_75 = io_axi_r_valid ? _GEN_58 : wb_buf_valid_13; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_76 = io_axi_r_valid ? _GEN_59 : wb_buf_valid_14; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_77 = io_axi_r_valid ? _GEN_60 : wb_buf_valid_15; // @[Icache.scala 113:22:@2827.6]
  assign _GEN_78 = _T_78 ? _GEN_29 : _GEN_62; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_79 = _T_78 ? _GEN_30 : _GEN_63; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_80 = _T_78 ? _GEN_31 : _GEN_64; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_81 = _T_78 ? _GEN_32 : _GEN_65; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_82 = _T_78 ? _GEN_33 : _GEN_66; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_83 = _T_78 ? _GEN_34 : _GEN_67; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_84 = _T_78 ? _GEN_35 : _GEN_68; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_85 = _T_78 ? _GEN_36 : _GEN_69; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_86 = _T_78 ? _GEN_37 : _GEN_70; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_87 = _T_78 ? _GEN_38 : _GEN_71; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_88 = _T_78 ? _GEN_39 : _GEN_72; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_89 = _T_78 ? _GEN_40 : _GEN_73; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_90 = _T_78 ? _GEN_41 : _GEN_74; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_91 = _T_78 ? _GEN_42 : _GEN_75; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_92 = _T_78 ? _GEN_43 : _GEN_76; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_93 = _T_78 ? _GEN_44 : _GEN_77; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_94 = _T_78 ? _GEN_28 : _GEN_28; // @[Icache.scala 105:31:@2802.4]
  assign _GEN_95 = 4'h0 == cnt ? io_axi_r_data : wb_buffer_0; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_96 = 4'h1 == cnt ? io_axi_r_data : wb_buffer_1; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_97 = 4'h2 == cnt ? io_axi_r_data : wb_buffer_2; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_98 = 4'h3 == cnt ? io_axi_r_data : wb_buffer_3; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_99 = 4'h4 == cnt ? io_axi_r_data : wb_buffer_4; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_100 = 4'h5 == cnt ? io_axi_r_data : wb_buffer_5; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_101 = 4'h6 == cnt ? io_axi_r_data : wb_buffer_6; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_102 = 4'h7 == cnt ? io_axi_r_data : wb_buffer_7; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_103 = 4'h8 == cnt ? io_axi_r_data : wb_buffer_8; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_104 = 4'h9 == cnt ? io_axi_r_data : wb_buffer_9; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_105 = 4'ha == cnt ? io_axi_r_data : wb_buffer_10; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_106 = 4'hb == cnt ? io_axi_r_data : wb_buffer_11; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_107 = 4'hc == cnt ? io_axi_r_data : wb_buffer_12; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_108 = 4'hd == cnt ? io_axi_r_data : wb_buffer_13; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_109 = 4'he == cnt ? io_axi_r_data : wb_buffer_14; // @[Icache.scala 118:34:@2834.6]
  assign _GEN_110 = 4'hf == cnt ? io_axi_r_data : wb_buffer_15; // @[Icache.scala 118:34:@2834.6]
  assign _T_283 = _T_91 & pc_valid; // @[Icache.scala 121:27:@2837.4]
  assign _T_284 = _T_283 & line_hit; // @[Icache.scala 121:39:@2838.4]
  assign _T_287 = _T_284 | _T_117; // @[Icache.scala 121:52:@2841.4]
  assign wait_inst_back = _T_287 | _T_119; // @[Icache.scala 122:39:@2844.4]
  assign line_idx = pc[5:2]; // @[Icache.scala 125:23:@2845.4]
  assign _GEN_128 = 4'h1 == line_idx ? wb_buffer_1 : wb_buffer_0; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_129 = 4'h2 == line_idx ? wb_buffer_2 : _GEN_128; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_130 = 4'h3 == line_idx ? wb_buffer_3 : _GEN_129; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_131 = 4'h4 == line_idx ? wb_buffer_4 : _GEN_130; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_132 = 4'h5 == line_idx ? wb_buffer_5 : _GEN_131; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_133 = 4'h6 == line_idx ? wb_buffer_6 : _GEN_132; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_134 = 4'h7 == line_idx ? wb_buffer_7 : _GEN_133; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_135 = 4'h8 == line_idx ? wb_buffer_8 : _GEN_134; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_136 = 4'h9 == line_idx ? wb_buffer_9 : _GEN_135; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_137 = 4'ha == line_idx ? wb_buffer_10 : _GEN_136; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_138 = 4'hb == line_idx ? wb_buffer_11 : _GEN_137; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_139 = 4'hc == line_idx ? wb_buffer_12 : _GEN_138; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_140 = 4'hd == line_idx ? wb_buffer_13 : _GEN_139; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_141 = 4'he == line_idx ? wb_buffer_14 : _GEN_140; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_142 = 4'hf == line_idx ? wb_buffer_15 : _GEN_141; // @[Icache.scala 126:24:@2846.4]
  assign buffer_inst = line_hit ? _GEN_142 : icache_io_rdata; // @[Icache.scala 126:24:@2846.4]
  assign _GEN_144 = 4'h1 == line_idx ? wb_buf_valid_1 : wb_buf_valid_0; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_145 = 4'h2 == line_idx ? wb_buf_valid_2 : _GEN_144; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_146 = 4'h3 == line_idx ? wb_buf_valid_3 : _GEN_145; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_147 = 4'h4 == line_idx ? wb_buf_valid_4 : _GEN_146; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_148 = 4'h5 == line_idx ? wb_buf_valid_5 : _GEN_147; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_149 = 4'h6 == line_idx ? wb_buf_valid_6 : _GEN_148; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_150 = 4'h7 == line_idx ? wb_buf_valid_7 : _GEN_149; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_151 = 4'h8 == line_idx ? wb_buf_valid_8 : _GEN_150; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_152 = 4'h9 == line_idx ? wb_buf_valid_9 : _GEN_151; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_153 = 4'ha == line_idx ? wb_buf_valid_10 : _GEN_152; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_154 = 4'hb == line_idx ? wb_buf_valid_11 : _GEN_153; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_155 = 4'hc == line_idx ? wb_buf_valid_12 : _GEN_154; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_156 = 4'hd == line_idx ? wb_buf_valid_13 : _GEN_155; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_157 = 4'he == line_idx ? wb_buf_valid_14 : _GEN_156; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_158 = 4'hf == line_idx ? wb_buf_valid_15 : _GEN_157; // @[Icache.scala 127:78:@2847.4]
  assign _T_294 = _GEN_158 & line_hit; // @[Icache.scala 127:78:@2847.4]
  assign _GEN_159 = wait_inst_back ? 1'h1 : _T_297; // @[Icache.scala 38:20:@2853.6]
  assign _GEN_160 = _T_294 ? 1'h0 : _GEN_159; // @[Icache.scala 37:17:@2849.4]
  assign _T_300 = wait_inst_back | _T_297; // @[Icache.scala 39:9:@2856.4]
  assign _T_301 = _T_300 & _T_294; // @[Icache.scala 39:22:@2857.4]
  assign buf_inst_valid = _T_301 | cache_hit; // @[Icache.scala 127:91:@2858.4]
  assign io_core_inst_valid = _T_87 ? cache_hit : buf_inst_valid; // @[Icache.scala 128:22:@2861.4]
  assign io_core_inst_bits = _T_87 ? icache_io_rdata : buffer_inst; // @[Icache.scala 129:22:@2864.4]
  assign io_core_ready = state != 2'h2; // @[Icache.scala 82:19:@2742.4]
  assign io_axi_ar_valid = pc_miss | _T_104; // @[Icache.scala 80:19:@2737.4]
  assign io_axi_ar_addr = {_T_84,6'h0}; // @[Icache.scala 81:19:@2740.4]
  assign icache_clock = clock; // @[:@2678.4]
  assign icache_reset = reset; // @[:@2679.4]
  assign icache_io_wen = state == 2'h2; // @[Icache.scala 67:21:@2681.4]
  assign icache_io_addr = _T_78 ? _T_81 : io_core_pc_bits; // @[Icache.scala 68:21:@2685.4]
  assign icache_io_wdata_0 = wb_buffer_0; // @[Icache.scala 69:21:@2686.4]
  assign icache_io_wdata_1 = wb_buffer_1; // @[Icache.scala 69:21:@2687.4]
  assign icache_io_wdata_2 = wb_buffer_2; // @[Icache.scala 69:21:@2688.4]
  assign icache_io_wdata_3 = wb_buffer_3; // @[Icache.scala 69:21:@2689.4]
  assign icache_io_wdata_4 = wb_buffer_4; // @[Icache.scala 69:21:@2690.4]
  assign icache_io_wdata_5 = wb_buffer_5; // @[Icache.scala 69:21:@2691.4]
  assign icache_io_wdata_6 = wb_buffer_6; // @[Icache.scala 69:21:@2692.4]
  assign icache_io_wdata_7 = wb_buffer_7; // @[Icache.scala 69:21:@2693.4]
  assign icache_io_wdata_8 = wb_buffer_8; // @[Icache.scala 69:21:@2694.4]
  assign icache_io_wdata_9 = wb_buffer_9; // @[Icache.scala 69:21:@2695.4]
  assign icache_io_wdata_10 = wb_buffer_10; // @[Icache.scala 69:21:@2696.4]
  assign icache_io_wdata_11 = wb_buffer_11; // @[Icache.scala 69:21:@2697.4]
  assign icache_io_wdata_12 = wb_buffer_12; // @[Icache.scala 69:21:@2698.4]
  assign icache_io_wdata_13 = wb_buffer_13; // @[Icache.scala 69:21:@2699.4]
  assign icache_io_wdata_14 = wb_buffer_14; // @[Icache.scala 69:21:@2700.4]
  assign icache_io_wdata_15 = wb_buffer_15; // @[Icache.scala 69:21:@2701.4]
  assign icache_io_wstatus = state == 2'h2; // @[Icache.scala 70:21:@2703.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_valid = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  wb_buffer_0 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  wb_buffer_1 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  wb_buffer_2 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  wb_buffer_3 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  wb_buffer_4 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  wb_buffer_5 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  wb_buffer_6 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  wb_buffer_7 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  wb_buffer_8 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  wb_buffer_9 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  wb_buffer_10 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  wb_buffer_11 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  wb_buffer_12 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  wb_buffer_13 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  wb_buffer_14 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  wb_buffer_15 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  wb_addr = _RAND_19[25:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  _T_99 = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  _T_104 = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  cnt = _RAND_22[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  wb_buf_valid_0 = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  wb_buf_valid_1 = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  wb_buf_valid_2 = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  wb_buf_valid_3 = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  wb_buf_valid_4 = _RAND_27[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  wb_buf_valid_5 = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  wb_buf_valid_6 = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  wb_buf_valid_7 = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  wb_buf_valid_8 = _RAND_31[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  wb_buf_valid_9 = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_buf_valid_10 = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wb_buf_valid_11 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wb_buf_valid_12 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wb_buf_valid_13 = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  wb_buf_valid_14 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  wb_buf_valid_15 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_297 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc_valid <= 1'h0;
    end else begin
      pc_valid <= pc_accept;
    end
    if (pc_accept) begin
      pc <= io_core_pc_bits;
    end
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_112) begin
        if (pc_miss) begin
          state <= 2'h1;
        end else begin
          state <= 2'h0;
        end
      end else begin
        if (_T_113) begin
          if (_T_114) begin
            state <= 2'h2;
          end else begin
            state <= 2'h1;
          end
        end else begin
          if (_T_115) begin
            if (pc_double_miss) begin
              state <= 2'h1;
            end else begin
              state <= 2'h0;
            end
          end
        end
      end
    end
    if (io_axi_r_valid) begin
      if (4'h0 == cnt) begin
        wb_buffer_0 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h1 == cnt) begin
        wb_buffer_1 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h2 == cnt) begin
        wb_buffer_2 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h3 == cnt) begin
        wb_buffer_3 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h4 == cnt) begin
        wb_buffer_4 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h5 == cnt) begin
        wb_buffer_5 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h6 == cnt) begin
        wb_buffer_6 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h7 == cnt) begin
        wb_buffer_7 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h8 == cnt) begin
        wb_buffer_8 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'h9 == cnt) begin
        wb_buffer_9 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'ha == cnt) begin
        wb_buffer_10 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hb == cnt) begin
        wb_buffer_11 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hc == cnt) begin
        wb_buffer_12 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hd == cnt) begin
        wb_buffer_13 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'he == cnt) begin
        wb_buffer_14 <= io_axi_r_data;
      end
    end
    if (io_axi_r_valid) begin
      if (4'hf == cnt) begin
        wb_buffer_15 <= io_axi_r_data;
      end
    end
    if (_T_120) begin
      wb_addr <= _T_84;
    end
    if (reset) begin
      _T_99 <= 1'h0;
    end else begin
      if (_T_78) begin
        _T_99 <= 1'h0;
      end else begin
        if (_T_95) begin
          _T_99 <= 1'h1;
        end
      end
    end
    if (reset) begin
      _T_104 <= 1'h0;
    end else begin
      if (io_axi_ar_ready) begin
        _T_104 <= 1'h0;
      end else begin
        if (pc_miss) begin
          _T_104 <= 1'h1;
        end
      end
    end
    if (reset) begin
      cnt <= 4'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          cnt <= _T_269;
        end
      end else begin
        if (io_axi_r_valid) begin
          cnt <= _T_269;
        end
      end
    end
    if (reset) begin
      wb_buf_valid_0 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_0 <= _GEN_12;
        end else begin
          wb_buf_valid_0 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h0 == cnt) begin
            wb_buf_valid_0 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_1 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_1 <= _GEN_13;
        end else begin
          wb_buf_valid_1 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h1 == cnt) begin
            wb_buf_valid_1 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_2 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_2 <= _GEN_14;
        end else begin
          wb_buf_valid_2 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h2 == cnt) begin
            wb_buf_valid_2 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_3 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_3 <= _GEN_15;
        end else begin
          wb_buf_valid_3 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h3 == cnt) begin
            wb_buf_valid_3 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_4 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_4 <= _GEN_16;
        end else begin
          wb_buf_valid_4 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h4 == cnt) begin
            wb_buf_valid_4 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_5 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_5 <= _GEN_17;
        end else begin
          wb_buf_valid_5 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h5 == cnt) begin
            wb_buf_valid_5 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_6 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_6 <= _GEN_18;
        end else begin
          wb_buf_valid_6 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h6 == cnt) begin
            wb_buf_valid_6 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_7 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_7 <= _GEN_19;
        end else begin
          wb_buf_valid_7 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h7 == cnt) begin
            wb_buf_valid_7 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_8 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_8 <= _GEN_20;
        end else begin
          wb_buf_valid_8 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h8 == cnt) begin
            wb_buf_valid_8 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_9 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_9 <= _GEN_21;
        end else begin
          wb_buf_valid_9 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'h9 == cnt) begin
            wb_buf_valid_9 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_10 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_10 <= _GEN_22;
        end else begin
          wb_buf_valid_10 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'ha == cnt) begin
            wb_buf_valid_10 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_11 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_11 <= _GEN_23;
        end else begin
          wb_buf_valid_11 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hb == cnt) begin
            wb_buf_valid_11 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_12 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_12 <= _GEN_24;
        end else begin
          wb_buf_valid_12 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hc == cnt) begin
            wb_buf_valid_12 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_13 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_13 <= _GEN_25;
        end else begin
          wb_buf_valid_13 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hd == cnt) begin
            wb_buf_valid_13 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_14 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_14 <= _GEN_26;
        end else begin
          wb_buf_valid_14 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'he == cnt) begin
            wb_buf_valid_14 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      wb_buf_valid_15 <= 1'h0;
    end else begin
      if (_T_78) begin
        if (io_axi_r_valid) begin
          wb_buf_valid_15 <= _GEN_27;
        end else begin
          wb_buf_valid_15 <= 1'h0;
        end
      end else begin
        if (io_axi_r_valid) begin
          if (4'hf == cnt) begin
            wb_buf_valid_15 <= 1'h1;
          end
        end
      end
    end
    if (reset) begin
      _T_297 <= 1'h0;
    end else begin
      if (_T_294) begin
        _T_297 <= 1'h0;
      end else begin
        if (wait_inst_back) begin
          _T_297 <= 1'h1;
        end
      end
    end
  end
endmodule
module FetchInst( // @[:@2866.2]
  input         clock, // @[:@2867.4]
  input         reset, // @[:@2868.4]
  input  [31:0] io_mem_r_data, // @[:@2869.4]
  input         io_mem_r_valid, // @[:@2869.4]
  input         io_mem_r_last, // @[:@2869.4]
  input         io_mem_ar_ready, // @[:@2869.4]
  output        io_mem_ar_valid, // @[:@2869.4]
  output [31:0] io_mem_ar_addr, // @[:@2869.4]
  input  [9:0]  io_if_btb_history, // @[:@2869.4]
  input         io_if_btb_diff, // @[:@2869.4]
  input  [31:0] io_if_btb_tgt, // @[:@2869.4]
  output [9:0]  io_dec_btb_history, // @[:@2869.4]
  output        io_dec_btb_diff, // @[:@2869.4]
  output [31:0] io_dec_btb_tgt, // @[:@2869.4]
  input  [31:0] io_if_pc, // @[:@2869.4]
  output [31:0] io_dec_pc, // @[:@2869.4]
  input         io_if_kill, // @[:@2869.4]
  input         io_dec_kill, // @[:@2869.4]
  output        io_pc_forward, // @[:@2869.4]
  input         io_forward, // @[:@2869.4]
  output        io_inst_valid, // @[:@2869.4]
  output [31:0] io_inst_bits // @[:@2869.4]
);
  wire  icache_clock; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_reset; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_core_pc_valid; // @[FetchInst.scala 35:22:@2873.4]
  wire [31:0] icache_io_core_pc_bits; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_core_inst_valid; // @[FetchInst.scala 35:22:@2873.4]
  wire [31:0] icache_io_core_inst_bits; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_core_ready; // @[FetchInst.scala 35:22:@2873.4]
  wire [31:0] icache_io_axi_r_data; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_axi_r_valid; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_axi_r_last; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_axi_ar_ready; // @[FetchInst.scala 35:22:@2873.4]
  wire  icache_io_axi_ar_valid; // @[FetchInst.scala 35:22:@2873.4]
  wire [31:0] icache_io_axi_ar_addr; // @[FetchInst.scala 35:22:@2873.4]
  reg [1:0] state; // @[FetchInst.scala 33:22:@2871.4]
  reg [31:0] _RAND_0;
  wire  _T_101; // @[FetchInst.scala 81:21:@2962.4]
  wire  inst_valid; // @[FetchInst.scala 49:20:@2902.4]
  reg  inst_kill; // @[FetchInst.scala 53:26:@2907.4]
  reg [31:0] _RAND_1;
  wire  _T_102; // @[FetchInst.scala 82:32:@2963.4]
  wire  _T_103; // @[FetchInst.scala 82:17:@2964.4]
  wire  _T_104; // @[FetchInst.scala 81:35:@2965.4]
  wire  _T_105; // @[FetchInst.scala 83:12:@2966.4]
  wire  _T_106; // @[FetchInst.scala 83:27:@2967.4]
  wire  pc_valid; // @[FetchInst.scala 82:47:@2968.4]
  wire  addr_ready; // @[FetchInst.scala 47:29:@2899.4]
  wire [31:0] inst_bits; // @[FetchInst.scala 50:20:@2905.4]
  wire  _T_86; // @[Conditional.scala 37:30:@2908.4]
  wire [1:0] _GEN_0; // @[FetchInst.scala 56:24:@2910.6]
  wire  _T_87; // @[Conditional.scala 37:30:@2915.6]
  wire [1:0] _T_89; // @[FetchInst.scala 61:23:@2920.12]
  wire [1:0] _GEN_1; // @[FetchInst.scala 62:33:@2924.12]
  wire [1:0] _GEN_2; // @[FetchInst.scala 60:39:@2919.10]
  wire [1:0] _GEN_3; // @[FetchInst.scala 59:24:@2917.8]
  wire  _T_90; // @[Conditional.scala 37:30:@2933.8]
  wire [1:0] _GEN_4; // @[FetchInst.scala 69:31:@2940.12]
  wire [1:0] _GEN_5; // @[FetchInst.scala 67:24:@2935.10]
  wire [1:0] _GEN_6; // @[Conditional.scala 39:67:@2934.8]
  wire [1:0] _GEN_7; // @[Conditional.scala 39:67:@2916.6]
  wire [1:0] _GEN_8; // @[Conditional.scala 40:58:@2909.4]
  wire  _T_93; // @[FetchInst.scala 76:35:@2952.8]
  wire  _T_94; // @[FetchInst.scala 76:26:@2953.8]
  wire  _GEN_9; // @[FetchInst.scala 76:50:@2954.8]
  wire  _GEN_10; // @[FetchInst.scala 74:26:@2948.6]
  wire  _GEN_11; // @[FetchInst.scala 72:19:@2944.4]
  wire  _T_97; // @[FetchInst.scala 80:35:@2957.4]
  wire  _T_98; // @[FetchInst.scala 80:32:@2958.4]
  wire  _T_108; // @[FetchInst.scala 84:46:@2970.4]
  reg [9:0] reg_pred_history; // @[FetchInst.scala 86:21:@2973.4]
  reg [31:0] _RAND_2;
  reg  reg_pred_diff; // @[FetchInst.scala 86:21:@2973.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_pred_tgt; // @[FetchInst.scala 86:21:@2973.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_pc; // @[FetchInst.scala 87:21:@2974.4]
  reg [31:0] _RAND_5;
  reg [31:0] _T_113; // @[FetchInst.scala 9:25:@2982.4]
  reg [31:0] _RAND_6;
  Icache icache ( // @[FetchInst.scala 35:22:@2873.4]
    .clock(icache_clock),
    .reset(icache_reset),
    .io_core_pc_valid(icache_io_core_pc_valid),
    .io_core_pc_bits(icache_io_core_pc_bits),
    .io_core_inst_valid(icache_io_core_inst_valid),
    .io_core_inst_bits(icache_io_core_inst_bits),
    .io_core_ready(icache_io_core_ready),
    .io_axi_r_data(icache_io_axi_r_data),
    .io_axi_r_valid(icache_io_axi_r_valid),
    .io_axi_r_last(icache_io_axi_r_last),
    .io_axi_ar_ready(icache_io_axi_ar_ready),
    .io_axi_ar_valid(icache_io_axi_ar_valid),
    .io_axi_ar_addr(icache_io_axi_ar_addr)
  );
  assign _T_101 = state == 2'h0; // @[FetchInst.scala 81:21:@2962.4]
  assign inst_valid = icache_io_core_inst_valid; // @[FetchInst.scala 49:20:@2902.4]
  assign _T_102 = io_forward | inst_kill; // @[FetchInst.scala 82:32:@2963.4]
  assign _T_103 = inst_valid & _T_102; // @[FetchInst.scala 82:17:@2964.4]
  assign _T_104 = _T_101 | _T_103; // @[FetchInst.scala 81:35:@2965.4]
  assign _T_105 = state == 2'h2; // @[FetchInst.scala 83:12:@2966.4]
  assign _T_106 = _T_105 & io_forward; // @[FetchInst.scala 83:27:@2967.4]
  assign pc_valid = _T_104 | _T_106; // @[FetchInst.scala 82:47:@2968.4]
  assign addr_ready = icache_io_core_ready; // @[FetchInst.scala 47:29:@2899.4]
  assign inst_bits = icache_io_core_inst_bits; // @[FetchInst.scala 50:20:@2905.4]
  assign _T_86 = 2'h0 == state; // @[Conditional.scala 37:30:@2908.4]
  assign _GEN_0 = addr_ready ? 2'h1 : state; // @[FetchInst.scala 56:24:@2910.6]
  assign _T_87 = 2'h1 == state; // @[Conditional.scala 37:30:@2915.6]
  assign _T_89 = addr_ready ? 2'h1 : 2'h0; // @[FetchInst.scala 61:23:@2920.12]
  assign _GEN_1 = io_dec_kill ? 2'h0 : 2'h2; // @[FetchInst.scala 62:33:@2924.12]
  assign _GEN_2 = _T_102 ? _T_89 : _GEN_1; // @[FetchInst.scala 60:39:@2919.10]
  assign _GEN_3 = inst_valid ? _GEN_2 : state; // @[FetchInst.scala 59:24:@2917.8]
  assign _T_90 = 2'h2 == state; // @[Conditional.scala 37:30:@2933.8]
  assign _GEN_4 = io_dec_kill ? 2'h0 : state; // @[FetchInst.scala 69:31:@2940.12]
  assign _GEN_5 = io_forward ? _T_89 : _GEN_4; // @[FetchInst.scala 67:24:@2935.10]
  assign _GEN_6 = _T_90 ? _GEN_5 : state; // @[Conditional.scala 39:67:@2934.8]
  assign _GEN_7 = _T_87 ? _GEN_3 : _GEN_6; // @[Conditional.scala 39:67:@2916.6]
  assign _GEN_8 = _T_86 ? _GEN_0 : _GEN_7; // @[Conditional.scala 40:58:@2909.4]
  assign _T_93 = state == 2'h1; // @[FetchInst.scala 76:35:@2952.8]
  assign _T_94 = io_dec_kill & _T_93; // @[FetchInst.scala 76:26:@2953.8]
  assign _GEN_9 = _T_94 ? 1'h1 : inst_kill; // @[FetchInst.scala 76:50:@2954.8]
  assign _GEN_10 = inst_valid ? 1'h0 : _GEN_9; // @[FetchInst.scala 74:26:@2948.6]
  assign _GEN_11 = pc_valid ? io_if_kill : _GEN_10; // @[FetchInst.scala 72:19:@2944.4]
  assign _T_97 = inst_kill == 1'h0; // @[FetchInst.scala 80:35:@2957.4]
  assign _T_98 = inst_valid & _T_97; // @[FetchInst.scala 80:32:@2958.4]
  assign _T_108 = addr_ready & pc_valid; // @[FetchInst.scala 84:46:@2970.4]
  assign io_mem_ar_valid = icache_io_axi_ar_valid; // @[FetchInst.scala 42:19:@2888.4]
  assign io_mem_ar_addr = icache_io_axi_ar_addr; // @[FetchInst.scala 43:19:@2890.4]
  assign io_dec_btb_history = reg_pred_history; // @[FetchInst.scala 95:14:@2990.4]
  assign io_dec_btb_diff = reg_pred_diff; // @[FetchInst.scala 95:14:@2989.4]
  assign io_dec_btb_tgt = reg_pred_tgt; // @[FetchInst.scala 95:14:@2988.4]
  assign io_dec_pc = reg_pc; // @[FetchInst.scala 96:14:@2992.4]
  assign io_pc_forward = io_if_kill | _T_108; // @[FetchInst.scala 84:17:@2972.4]
  assign io_inst_valid = _T_98 | _T_105; // @[FetchInst.scala 80:17:@2961.4]
  assign io_inst_bits = inst_valid ? inst_bits : _T_113; // @[FetchInst.scala 94:16:@2987.4]
  assign icache_clock = clock; // @[:@2874.4]
  assign icache_reset = reset; // @[:@2875.4]
  assign icache_io_core_pc_valid = _T_104 | _T_106; // @[FetchInst.scala 40:27:@2884.4]
  assign icache_io_core_pc_bits = io_if_pc; // @[FetchInst.scala 39:26:@2882.4]
  assign icache_io_axi_r_data = io_mem_r_data; // @[FetchInst.scala 37:19:@2880.4]
  assign icache_io_axi_r_valid = io_mem_r_valid; // @[FetchInst.scala 37:19:@2879.4]
  assign icache_io_axi_r_last = io_mem_r_last; // @[FetchInst.scala 37:19:@2878.4]
  assign icache_io_axi_ar_ready = io_mem_ar_ready; // @[FetchInst.scala 38:26:@2881.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  state = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inst_kill = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_pred_history = _RAND_2[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_pred_diff = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_pred_tgt = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  _T_113 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      state <= 2'h0;
    end else begin
      if (_T_86) begin
        if (addr_ready) begin
          state <= 2'h1;
        end
      end else begin
        if (_T_87) begin
          if (inst_valid) begin
            if (_T_102) begin
              if (addr_ready) begin
                state <= 2'h1;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (io_dec_kill) begin
                state <= 2'h0;
              end else begin
                state <= 2'h2;
              end
            end
          end
        end else begin
          if (_T_90) begin
            if (io_forward) begin
              if (addr_ready) begin
                state <= 2'h1;
              end else begin
                state <= 2'h0;
              end
            end else begin
              if (io_dec_kill) begin
                state <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      inst_kill <= 1'h0;
    end else begin
      if (pc_valid) begin
        inst_kill <= io_if_kill;
      end else begin
        if (inst_valid) begin
          inst_kill <= 1'h0;
        end else begin
          if (_T_94) begin
            inst_kill <= 1'h1;
          end
        end
      end
    end
    if (pc_valid) begin
      reg_pred_history <= io_if_btb_history;
    end
    if (pc_valid) begin
      reg_pred_diff <= io_if_btb_diff;
    end
    if (pc_valid) begin
      reg_pred_tgt <= io_if_btb_tgt;
    end
    if (pc_valid) begin
      reg_pc <= io_if_pc;
    end
    if (inst_valid) begin
      _T_113 <= inst_bits;
    end
  end
endmodule
module MicroDecoder( // @[:@2994.2]
  input  [31:0] io_inst, // @[:@2997.4]
  output        io_isbrnch // @[:@2997.4]
);
  wire [4:0] func; // @[MicroDecoder.scala 21:22:@2999.4]
  assign func = io_inst[6:2]; // @[MicroDecoder.scala 21:22:@2999.4]
  assign io_isbrnch = func == 5'h18; // @[MicroDecoder.scala 34:14:@3012.4]
endmodule
module FrontEnd( // @[:@3085.2]
  input         clock, // @[:@3086.4]
  input         reset, // @[:@3087.4]
  input  [31:0] io_cyc, // @[:@3088.4]
  input  [31:0] io_mem_r_data, // @[:@3088.4]
  input         io_mem_r_valid, // @[:@3088.4]
  input         io_mem_r_last, // @[:@3088.4]
  input         io_mem_ar_ready, // @[:@3088.4]
  output        io_mem_ar_valid, // @[:@3088.4]
  output [31:0] io_mem_ar_addr, // @[:@3088.4]
  input         io_back_xcpt_valid, // @[:@3088.4]
  input  [31:0] io_back_xcpt_bits, // @[:@3088.4]
  input         io_back_kill, // @[:@3088.4]
  input         io_back_forward, // @[:@3088.4]
  output        io_back_inst_valid, // @[:@3088.4]
  output [31:0] io_back_inst_bits, // @[:@3088.4]
  output [31:0] io_back_pc, // @[:@3088.4]
  output [9:0]  io_back_pred_history, // @[:@3088.4]
  output        io_back_pred_diff, // @[:@3088.4]
  output [31:0] io_back_pred_tgt, // @[:@3088.4]
  input         io_back_ras_pop, // @[:@3088.4]
  input         io_back_ras_push_valid, // @[:@3088.4]
  input  [31:0] io_back_ras_push_bits, // @[:@3088.4]
  input  [31:0] io_back_fb_pc, // @[:@3088.4]
  input  [1:0]  io_back_fb_type, // @[:@3088.4]
  input         io_back_feedBack_redirect, // @[:@3088.4]
  input  [9:0]  io_back_feedBack_history, // @[:@3088.4]
  input         io_back_feedBack_diff, // @[:@3088.4]
  input  [31:0] io_back_feedBack_tgt, // @[:@3088.4]
  input         io_back_feedBack_valid // @[:@3088.4]
);
  wire  BTB_clock; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_reset; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_if_pc; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_predict_redirect; // @[FrontEnd.scala 12:24:@3090.4]
  wire [9:0] BTB_io_predict_history; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_predict_diff; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_predict_tgt; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_branch; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_forward; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_ras_pop; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_ras_push_valid; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_ras_push_bits; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_fb_pc; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_fb_miss; // @[FrontEnd.scala 12:24:@3090.4]
  wire [1:0] BTB_io_fb_type; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_feedBack_redirect; // @[FrontEnd.scala 12:24:@3090.4]
  wire [9:0] BTB_io_feedBack_history; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_feedBack_diff; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_feedBack_tgt; // @[FrontEnd.scala 12:24:@3090.4]
  wire  BTB_io_feedBack_valid; // @[FrontEnd.scala 12:24:@3090.4]
  wire [31:0] BTB_io_cyc; // @[FrontEnd.scala 12:24:@3090.4]
  wire  FetchInst_clock; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_reset; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_mem_r_data; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_mem_r_valid; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_mem_r_last; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_mem_ar_ready; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_mem_ar_valid; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_mem_ar_addr; // @[FrontEnd.scala 13:24:@3093.4]
  wire [9:0] FetchInst_io_if_btb_history; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_if_btb_diff; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_if_btb_tgt; // @[FrontEnd.scala 13:24:@3093.4]
  wire [9:0] FetchInst_io_dec_btb_history; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_dec_btb_diff; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_dec_btb_tgt; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_if_pc; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_dec_pc; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_if_kill; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_dec_kill; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_pc_forward; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_forward; // @[FrontEnd.scala 13:24:@3093.4]
  wire  FetchInst_io_inst_valid; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] FetchInst_io_inst_bits; // @[FrontEnd.scala 13:24:@3093.4]
  wire [31:0] MicroDecoder_io_inst; // @[FrontEnd.scala 14:24:@3096.4]
  wire  MicroDecoder_io_isbrnch; // @[FrontEnd.scala 14:24:@3096.4]
  reg [31:0] if_reg_pc; // @[FrontEnd.scala 15:27:@3099.4]
  reg [31:0] _RAND_0;
  wire [31:0] _T_74; // @[FrontEnd.scala 53:10:@3147.4]
  wire [31:0] if_pc_next; // @[FrontEnd.scala 52:10:@3148.4]
  wire [31:0] _GEN_0; // @[FrontEnd.scala 62:28:@3150.4]
  wire  _T_77; // @[FrontEnd.scala 63:9:@3153.4]
  wire  _T_78; // @[FrontEnd.scala 63:26:@3154.4]
  wire  _T_81; // @[FrontEnd.scala 64:11:@3157.6]
  BTB BTB ( // @[FrontEnd.scala 12:24:@3090.4]
    .clock(BTB_clock),
    .reset(BTB_reset),
    .io_if_pc(BTB_io_if_pc),
    .io_predict_redirect(BTB_io_predict_redirect),
    .io_predict_history(BTB_io_predict_history),
    .io_predict_diff(BTB_io_predict_diff),
    .io_predict_tgt(BTB_io_predict_tgt),
    .io_branch(BTB_io_branch),
    .io_forward(BTB_io_forward),
    .io_ras_pop(BTB_io_ras_pop),
    .io_ras_push_valid(BTB_io_ras_push_valid),
    .io_ras_push_bits(BTB_io_ras_push_bits),
    .io_fb_pc(BTB_io_fb_pc),
    .io_fb_miss(BTB_io_fb_miss),
    .io_fb_type(BTB_io_fb_type),
    .io_feedBack_redirect(BTB_io_feedBack_redirect),
    .io_feedBack_history(BTB_io_feedBack_history),
    .io_feedBack_diff(BTB_io_feedBack_diff),
    .io_feedBack_tgt(BTB_io_feedBack_tgt),
    .io_feedBack_valid(BTB_io_feedBack_valid),
    .io_cyc(BTB_io_cyc)
  );
  FetchInst FetchInst ( // @[FrontEnd.scala 13:24:@3093.4]
    .clock(FetchInst_clock),
    .reset(FetchInst_reset),
    .io_mem_r_data(FetchInst_io_mem_r_data),
    .io_mem_r_valid(FetchInst_io_mem_r_valid),
    .io_mem_r_last(FetchInst_io_mem_r_last),
    .io_mem_ar_ready(FetchInst_io_mem_ar_ready),
    .io_mem_ar_valid(FetchInst_io_mem_ar_valid),
    .io_mem_ar_addr(FetchInst_io_mem_ar_addr),
    .io_if_btb_history(FetchInst_io_if_btb_history),
    .io_if_btb_diff(FetchInst_io_if_btb_diff),
    .io_if_btb_tgt(FetchInst_io_if_btb_tgt),
    .io_dec_btb_history(FetchInst_io_dec_btb_history),
    .io_dec_btb_diff(FetchInst_io_dec_btb_diff),
    .io_dec_btb_tgt(FetchInst_io_dec_btb_tgt),
    .io_if_pc(FetchInst_io_if_pc),
    .io_dec_pc(FetchInst_io_dec_pc),
    .io_if_kill(FetchInst_io_if_kill),
    .io_dec_kill(FetchInst_io_dec_kill),
    .io_pc_forward(FetchInst_io_pc_forward),
    .io_forward(FetchInst_io_forward),
    .io_inst_valid(FetchInst_io_inst_valid),
    .io_inst_bits(FetchInst_io_inst_bits)
  );
  MicroDecoder MicroDecoder ( // @[FrontEnd.scala 14:24:@3096.4]
    .io_inst(MicroDecoder_io_inst),
    .io_isbrnch(MicroDecoder_io_isbrnch)
  );
  assign _T_74 = io_back_kill ? io_back_feedBack_tgt : BTB_io_predict_tgt; // @[FrontEnd.scala 53:10:@3147.4]
  assign if_pc_next = io_back_xcpt_valid ? io_back_xcpt_bits : _T_74; // @[FrontEnd.scala 52:10:@3148.4]
  assign _GEN_0 = FetchInst_io_pc_forward ? if_pc_next : if_reg_pc; // @[FrontEnd.scala 62:28:@3150.4]
  assign _T_77 = io_back_forward == 1'h0; // @[FrontEnd.scala 63:9:@3153.4]
  assign _T_78 = _T_77 & io_back_inst_valid; // @[FrontEnd.scala 63:26:@3154.4]
  assign _T_81 = reset == 1'h0; // @[FrontEnd.scala 64:11:@3157.6]
  assign io_mem_ar_valid = FetchInst_io_mem_ar_valid; // @[FrontEnd.scala 18:19:@3107.4]
  assign io_mem_ar_addr = FetchInst_io_mem_ar_addr; // @[FrontEnd.scala 18:19:@3105.4]
  assign io_back_inst_valid = FetchInst_io_inst_valid; // @[FrontEnd.scala 29:16:@3125.4]
  assign io_back_inst_bits = FetchInst_io_inst_bits; // @[FrontEnd.scala 29:16:@3124.4]
  assign io_back_pc = FetchInst_io_dec_pc; // @[FrontEnd.scala 30:16:@3126.4]
  assign io_back_pred_history = FetchInst_io_dec_btb_history; // @[FrontEnd.scala 31:16:@3129.4]
  assign io_back_pred_diff = FetchInst_io_dec_btb_diff; // @[FrontEnd.scala 31:16:@3128.4]
  assign io_back_pred_tgt = FetchInst_io_dec_btb_tgt; // @[FrontEnd.scala 31:16:@3127.4]
  assign BTB_clock = clock; // @[:@3091.4]
  assign BTB_reset = reset; // @[:@3092.4]
  assign BTB_io_if_pc = if_reg_pc; // @[FrontEnd.scala 39:13:@3131.4]
  assign BTB_io_branch = FetchInst_io_inst_valid & MicroDecoder_io_isbrnch; // @[FrontEnd.scala 41:16:@3134.4]
  assign BTB_io_forward = FetchInst_io_pc_forward; // @[FrontEnd.scala 40:16:@3132.4]
  assign BTB_io_ras_pop = io_back_ras_pop; // @[FrontEnd.scala 43:16:@3137.4]
  assign BTB_io_ras_push_valid = io_back_ras_push_valid; // @[FrontEnd.scala 42:16:@3136.4]
  assign BTB_io_ras_push_bits = io_back_ras_push_bits; // @[FrontEnd.scala 42:16:@3135.4]
  assign BTB_io_fb_pc = io_back_fb_pc; // @[FrontEnd.scala 45:16:@3139.4]
  assign BTB_io_fb_miss = io_back_kill; // @[FrontEnd.scala 44:16:@3138.4]
  assign BTB_io_fb_type = io_back_fb_type; // @[FrontEnd.scala 46:16:@3140.4]
  assign BTB_io_feedBack_redirect = io_back_feedBack_redirect; // @[FrontEnd.scala 47:16:@3145.4]
  assign BTB_io_feedBack_history = io_back_feedBack_history; // @[FrontEnd.scala 47:16:@3144.4]
  assign BTB_io_feedBack_diff = io_back_feedBack_diff; // @[FrontEnd.scala 47:16:@3143.4]
  assign BTB_io_feedBack_tgt = io_back_feedBack_tgt; // @[FrontEnd.scala 47:16:@3142.4]
  assign BTB_io_feedBack_valid = io_back_feedBack_valid; // @[FrontEnd.scala 47:16:@3141.4]
  assign BTB_io_cyc = io_cyc; // @[FrontEnd.scala 16:14:@3100.4]
  assign FetchInst_clock = clock; // @[:@3094.4]
  assign FetchInst_reset = reset; // @[:@3095.4]
  assign FetchInst_io_mem_r_data = io_mem_r_data; // @[FrontEnd.scala 18:19:@3112.4]
  assign FetchInst_io_mem_r_valid = io_mem_r_valid; // @[FrontEnd.scala 18:19:@3111.4]
  assign FetchInst_io_mem_r_last = io_mem_r_last; // @[FrontEnd.scala 18:19:@3110.4]
  assign FetchInst_io_mem_ar_ready = io_mem_ar_ready; // @[FrontEnd.scala 18:19:@3108.4]
  assign FetchInst_io_if_btb_history = BTB_io_predict_history; // @[FrontEnd.scala 20:19:@3116.4]
  assign FetchInst_io_if_btb_diff = BTB_io_predict_diff; // @[FrontEnd.scala 20:19:@3115.4]
  assign FetchInst_io_if_btb_tgt = BTB_io_predict_tgt; // @[FrontEnd.scala 20:19:@3114.4]
  assign FetchInst_io_if_pc = if_reg_pc; // @[FrontEnd.scala 19:19:@3113.4]
  assign FetchInst_io_if_kill = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 21:19:@3119.4]
  assign FetchInst_io_dec_kill = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 22:19:@3121.4]
  assign FetchInst_io_forward = io_back_forward; // @[FrontEnd.scala 23:19:@3122.4]
  assign MicroDecoder_io_inst = FetchInst_io_inst_bits; // @[FrontEnd.scala 24:19:@3123.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_reg_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      if_reg_pc <= 32'h80000000;
    end else begin
      if (FetchInst_io_pc_forward) begin
        if (io_back_xcpt_valid) begin
          if_reg_pc <= io_back_xcpt_bits;
        end else begin
          if (io_back_kill) begin
            if_reg_pc <= io_back_feedBack_tgt;
          end else begin
            if_reg_pc <= BTB_io_predict_tgt;
          end
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_78 & _T_81) begin
          $fwrite(32'h80000002,"STALL\n"); // @[FrontEnd.scala 64:11:@3159.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSRFile( // @[:@3163.2]
  input         clock, // @[:@3164.4]
  input         reset, // @[:@3165.4]
  input  [2:0]  io_rw_cmd, // @[:@3166.4]
  input  [11:0] io_rw_addr, // @[:@3166.4]
  output [31:0] io_rw_rdata, // @[:@3166.4]
  input  [31:0] io_rw_wdata, // @[:@3166.4]
  output        io_eret, // @[:@3166.4]
  output [1:0]  io_status_prv, // @[:@3166.4]
  output [13:0] io_status_unimp5, // @[:@3166.4]
  output        io_status_mprv, // @[:@3166.4]
  output [1:0]  io_status_unimp4, // @[:@3166.4]
  output [1:0]  io_status_mpp, // @[:@3166.4]
  output [2:0]  io_status_unimp3, // @[:@3166.4]
  output        io_status_mpie, // @[:@3166.4]
  output [2:0]  io_status_unimp2, // @[:@3166.4]
  output        io_status_mie, // @[:@3166.4]
  output [2:0]  io_status_unimp1, // @[:@3166.4]
  input         io_xcpt, // @[:@3166.4]
  input  [31:0] io_cause, // @[:@3166.4]
  input  [31:0] io_tval, // @[:@3166.4]
  output [31:0] io_evec, // @[:@3166.4]
  input         io_illegal, // @[:@3166.4]
  input  [1:0]  io_retire, // @[:@3166.4]
  input  [31:0] io_pc, // @[:@3166.4]
  output [31:0] io_time // @[:@3166.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 112:28:@3293.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 112:28:@3293.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 112:28:@3293.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[CSR.scala 113:21:@3294.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[CSR.scala 114:23:@3295.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[CSR.scala 115:22:@3296.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[CSR.scala 116:25:@3297.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[CSR.scala 118:24:@3299.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[CSR.scala 120:24:@3317.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[CSR.scala 120:24:@3317.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[CSR.scala 121:24:@3335.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[CSR.scala 121:24:@3335.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_240; // @[Util.scala 112:41:@3338.4]
  reg [31:0] _RAND_12;
  wire [6:0] _T_241; // @[Util.scala 113:33:@3339.4]
  reg [57:0] _T_244; // @[Util.scala 117:31:@3341.4]
  reg [63:0] _RAND_13;
  wire  _T_245; // @[Util.scala 118:20:@3342.4]
  wire [58:0] _T_247; // @[Util.scala 118:43:@3344.6]
  wire [57:0] _T_248; // @[Util.scala 118:43:@3345.6]
  wire [57:0] _GEN_0; // @[Util.scala 118:34:@3343.4]
  wire [63:0] _T_249; // @[Cat.scala 30:58:@3348.4]
  reg [5:0] _T_252; // @[Util.scala 112:41:@3349.4]
  reg [31:0] _RAND_14;
  wire [5:0] _GEN_147; // @[Util.scala 113:33:@3350.4]
  wire [6:0] _T_253; // @[Util.scala 113:33:@3350.4]
  reg [57:0] _T_256; // @[Util.scala 117:31:@3352.4]
  reg [63:0] _RAND_15;
  wire  _T_257; // @[Util.scala 118:20:@3353.4]
  wire [58:0] _T_259; // @[Util.scala 118:43:@3355.6]
  wire [57:0] _T_260; // @[Util.scala 118:43:@3356.6]
  wire [57:0] _GEN_1; // @[Util.scala 118:34:@3354.4]
  wire [63:0] _T_261; // @[Cat.scala 30:58:@3359.4]
  reg [39:0] _T_264; // @[Util.scala 112:74:@3361.4]
  reg [63:0] _RAND_16;
  wire [40:0] _T_265; // @[Util.scala 113:33:@3362.4]
  reg [39:0] _T_267; // @[Util.scala 112:74:@3364.4]
  reg [63:0] _RAND_17;
  wire [40:0] _T_268; // @[Util.scala 113:33:@3365.4]
  reg [39:0] _T_270; // @[Util.scala 112:74:@3367.4]
  reg [63:0] _RAND_18;
  wire [40:0] _T_271; // @[Util.scala 113:33:@3368.4]
  reg [39:0] _T_273; // @[Util.scala 112:74:@3370.4]
  reg [63:0] _RAND_19;
  wire [40:0] _T_274; // @[Util.scala 113:33:@3371.4]
  reg [39:0] _T_276; // @[Util.scala 112:74:@3373.4]
  reg [63:0] _RAND_20;
  wire [40:0] _T_277; // @[Util.scala 113:33:@3374.4]
  reg [39:0] _T_279; // @[Util.scala 112:74:@3376.4]
  reg [63:0] _RAND_21;
  wire [40:0] _T_280; // @[Util.scala 113:33:@3377.4]
  reg [39:0] _T_282; // @[Util.scala 112:74:@3379.4]
  reg [63:0] _RAND_22;
  wire [40:0] _T_283; // @[Util.scala 113:33:@3380.4]
  reg [39:0] _T_285; // @[Util.scala 112:74:@3382.4]
  reg [63:0] _RAND_23;
  wire [40:0] _T_286; // @[Util.scala 113:33:@3383.4]
  reg [39:0] _T_288; // @[Util.scala 112:74:@3385.4]
  reg [63:0] _RAND_24;
  wire [40:0] _T_289; // @[Util.scala 113:33:@3386.4]
  reg [39:0] _T_291; // @[Util.scala 112:74:@3388.4]
  reg [63:0] _RAND_25;
  wire [40:0] _T_292; // @[Util.scala 113:33:@3389.4]
  reg [39:0] _T_294; // @[Util.scala 112:74:@3391.4]
  reg [63:0] _RAND_26;
  wire [40:0] _T_295; // @[Util.scala 113:33:@3392.4]
  reg [39:0] _T_297; // @[Util.scala 112:74:@3394.4]
  reg [63:0] _RAND_27;
  wire [40:0] _T_298; // @[Util.scala 113:33:@3395.4]
  reg [39:0] _T_300; // @[Util.scala 112:74:@3397.4]
  reg [63:0] _RAND_28;
  wire [40:0] _T_301; // @[Util.scala 113:33:@3398.4]
  reg [39:0] _T_303; // @[Util.scala 112:74:@3400.4]
  reg [63:0] _RAND_29;
  wire [40:0] _T_304; // @[Util.scala 113:33:@3401.4]
  reg [39:0] _T_306; // @[Util.scala 112:74:@3403.4]
  reg [63:0] _RAND_30;
  wire [40:0] _T_307; // @[Util.scala 113:33:@3404.4]
  reg [39:0] _T_309; // @[Util.scala 112:74:@3406.4]
  reg [63:0] _RAND_31;
  wire [40:0] _T_310; // @[Util.scala 113:33:@3407.4]
  reg [39:0] _T_312; // @[Util.scala 112:74:@3409.4]
  reg [63:0] _RAND_32;
  wire [40:0] _T_313; // @[Util.scala 113:33:@3410.4]
  reg [39:0] _T_315; // @[Util.scala 112:74:@3412.4]
  reg [63:0] _RAND_33;
  wire [40:0] _T_316; // @[Util.scala 113:33:@3413.4]
  reg [39:0] _T_318; // @[Util.scala 112:74:@3415.4]
  reg [63:0] _RAND_34;
  wire [40:0] _T_319; // @[Util.scala 113:33:@3416.4]
  reg [39:0] _T_321; // @[Util.scala 112:74:@3418.4]
  reg [63:0] _RAND_35;
  wire [40:0] _T_322; // @[Util.scala 113:33:@3419.4]
  reg [39:0] _T_324; // @[Util.scala 112:74:@3421.4]
  reg [63:0] _RAND_36;
  wire [40:0] _T_325; // @[Util.scala 113:33:@3422.4]
  reg [39:0] _T_327; // @[Util.scala 112:74:@3424.4]
  reg [63:0] _RAND_37;
  wire [40:0] _T_328; // @[Util.scala 113:33:@3425.4]
  reg [39:0] _T_330; // @[Util.scala 112:74:@3427.4]
  reg [63:0] _RAND_38;
  wire [40:0] _T_331; // @[Util.scala 113:33:@3428.4]
  reg [39:0] _T_333; // @[Util.scala 112:74:@3430.4]
  reg [63:0] _RAND_39;
  wire [40:0] _T_334; // @[Util.scala 113:33:@3431.4]
  reg [39:0] _T_336; // @[Util.scala 112:74:@3433.4]
  reg [63:0] _RAND_40;
  wire [40:0] _T_337; // @[Util.scala 113:33:@3434.4]
  reg [39:0] _T_339; // @[Util.scala 112:74:@3436.4]
  reg [63:0] _RAND_41;
  wire [40:0] _T_340; // @[Util.scala 113:33:@3437.4]
  reg [39:0] _T_342; // @[Util.scala 112:74:@3439.4]
  reg [63:0] _RAND_42;
  wire [40:0] _T_343; // @[Util.scala 113:33:@3440.4]
  reg [39:0] _T_345; // @[Util.scala 112:74:@3442.4]
  reg [63:0] _RAND_43;
  wire [40:0] _T_346; // @[Util.scala 113:33:@3443.4]
  reg [39:0] _T_348; // @[Util.scala 112:74:@3445.4]
  reg [63:0] _RAND_44;
  wire [40:0] _T_349; // @[Util.scala 113:33:@3446.4]
  reg [39:0] _T_351; // @[Util.scala 112:74:@3448.4]
  reg [63:0] _RAND_45;
  wire [40:0] _T_352; // @[Util.scala 113:33:@3449.4]
  reg [39:0] _T_354; // @[Util.scala 112:74:@3451.4]
  reg [63:0] _RAND_46;
  wire [40:0] _T_355; // @[Util.scala 113:33:@3452.4]
  reg [39:0] _T_357; // @[Util.scala 112:74:@3454.4]
  reg [63:0] _RAND_47;
  wire [40:0] _T_358; // @[Util.scala 113:33:@3455.4]
  reg [31:0] reg_dscratch; // @[CSR.scala 134:25:@3544.4]
  reg [31:0] _RAND_48;
  wire  system_insn; // @[CSR.scala 137:31:@3546.4]
  wire  _T_446; // @[CSR.scala 138:27:@3547.4]
  wire  _T_448; // @[CSR.scala 138:40:@3548.4]
  wire  cpu_ren; // @[CSR.scala 138:37:@3549.4]
  wire [31:0] read_mstatus; // @[CSR.scala 140:32:@3558.4]
  wire [15:0] _T_468; // @[CSR.scala 156:25:@3564.4]
  wire [15:0] _T_474; // @[CSR.scala 157:25:@3570.4]
  wire  _T_478; // @[CSR.scala 177:73:@3571.4]
  wire  _T_480; // @[CSR.scala 177:73:@3572.4]
  wire  _T_482; // @[CSR.scala 177:73:@3573.4]
  wire  _T_488; // @[CSR.scala 177:73:@3576.4]
  wire  _T_490; // @[CSR.scala 177:73:@3577.4]
  wire  _T_492; // @[CSR.scala 177:73:@3578.4]
  wire  _T_494; // @[CSR.scala 177:73:@3579.4]
  wire  _T_496; // @[CSR.scala 177:73:@3580.4]
  wire  _T_498; // @[CSR.scala 177:73:@3581.4]
  wire  _T_500; // @[CSR.scala 177:73:@3582.4]
  wire  _T_502; // @[CSR.scala 177:73:@3583.4]
  wire  _T_504; // @[CSR.scala 177:73:@3584.4]
  wire  _T_508; // @[CSR.scala 177:73:@3586.4]
  wire  _T_510; // @[CSR.scala 177:73:@3587.4]
  wire  _T_512; // @[CSR.scala 177:73:@3588.4]
  wire  _T_514; // @[CSR.scala 177:73:@3589.4]
  wire  _T_516; // @[CSR.scala 177:73:@3590.4]
  wire  _T_518; // @[CSR.scala 177:73:@3591.4]
  wire  _T_520; // @[CSR.scala 177:73:@3592.4]
  wire  _T_522; // @[CSR.scala 177:73:@3593.4]
  wire  _T_524; // @[CSR.scala 177:73:@3594.4]
  wire  _T_526; // @[CSR.scala 177:73:@3595.4]
  wire  _T_528; // @[CSR.scala 177:73:@3596.4]
  wire  _T_530; // @[CSR.scala 177:73:@3597.4]
  wire  _T_532; // @[CSR.scala 177:73:@3598.4]
  wire  _T_534; // @[CSR.scala 177:73:@3599.4]
  wire  _T_536; // @[CSR.scala 177:73:@3600.4]
  wire  _T_538; // @[CSR.scala 177:73:@3601.4]
  wire  _T_540; // @[CSR.scala 177:73:@3602.4]
  wire  _T_542; // @[CSR.scala 177:73:@3603.4]
  wire  _T_544; // @[CSR.scala 177:73:@3604.4]
  wire  _T_546; // @[CSR.scala 177:73:@3605.4]
  wire  _T_548; // @[CSR.scala 177:73:@3606.4]
  wire  _T_550; // @[CSR.scala 177:73:@3607.4]
  wire  _T_552; // @[CSR.scala 177:73:@3608.4]
  wire  _T_554; // @[CSR.scala 177:73:@3609.4]
  wire  _T_556; // @[CSR.scala 177:73:@3610.4]
  wire  _T_558; // @[CSR.scala 177:73:@3611.4]
  wire  _T_560; // @[CSR.scala 177:73:@3612.4]
  wire  _T_562; // @[CSR.scala 177:73:@3613.4]
  wire  _T_564; // @[CSR.scala 177:73:@3614.4]
  wire  _T_566; // @[CSR.scala 177:73:@3615.4]
  wire  _T_568; // @[CSR.scala 177:73:@3616.4]
  wire  _T_570; // @[CSR.scala 177:73:@3617.4]
  wire  _T_572; // @[CSR.scala 177:73:@3618.4]
  wire  _T_574; // @[CSR.scala 177:73:@3619.4]
  wire  _T_576; // @[CSR.scala 177:73:@3620.4]
  wire  _T_578; // @[CSR.scala 177:73:@3621.4]
  wire  _T_580; // @[CSR.scala 177:73:@3622.4]
  wire  _T_582; // @[CSR.scala 177:73:@3623.4]
  wire  _T_584; // @[CSR.scala 177:73:@3624.4]
  wire  _T_586; // @[CSR.scala 177:73:@3625.4]
  wire  _T_588; // @[CSR.scala 177:73:@3626.4]
  wire  _T_590; // @[CSR.scala 177:73:@3627.4]
  wire  _T_592; // @[CSR.scala 177:73:@3628.4]
  wire  _T_594; // @[CSR.scala 177:73:@3629.4]
  wire  _T_596; // @[CSR.scala 177:73:@3630.4]
  wire  _T_598; // @[CSR.scala 177:73:@3631.4]
  wire  _T_600; // @[CSR.scala 177:73:@3632.4]
  wire  _T_602; // @[CSR.scala 177:73:@3633.4]
  wire  _T_604; // @[CSR.scala 177:73:@3634.4]
  wire  _T_606; // @[CSR.scala 177:73:@3635.4]
  wire  _T_608; // @[CSR.scala 177:73:@3636.4]
  wire  _T_610; // @[CSR.scala 177:73:@3637.4]
  wire  _T_612; // @[CSR.scala 177:73:@3638.4]
  wire  _T_614; // @[CSR.scala 177:73:@3639.4]
  wire  _T_616; // @[CSR.scala 177:73:@3640.4]
  wire  _T_618; // @[CSR.scala 177:73:@3641.4]
  wire  _T_620; // @[CSR.scala 177:73:@3642.4]
  wire  _T_622; // @[CSR.scala 177:73:@3643.4]
  wire  _T_624; // @[CSR.scala 177:73:@3644.4]
  wire  _T_626; // @[CSR.scala 177:73:@3645.4]
  wire  _T_628; // @[CSR.scala 177:73:@3646.4]
  wire  _T_630; // @[CSR.scala 177:73:@3647.4]
  wire  _T_632; // @[CSR.scala 177:73:@3648.4]
  wire  _T_634; // @[CSR.scala 177:73:@3649.4]
  wire  _T_636; // @[CSR.scala 177:73:@3650.4]
  wire  _T_638; // @[CSR.scala 177:73:@3651.4]
  wire  _T_640; // @[CSR.scala 177:73:@3652.4]
  wire  _T_642; // @[CSR.scala 177:73:@3653.4]
  wire [1:0] _T_643; // @[CSR.scala 179:54:@3654.4]
  wire  priv_sufficient; // @[CSR.scala 179:41:@3655.4]
  wire [1:0] _T_644; // @[CSR.scala 180:29:@3656.4]
  wire [1:0] _T_645; // @[CSR.scala 180:37:@3657.4]
  wire  read_only; // @[CSR.scala 180:37:@3658.4]
  wire  _T_647; // @[CSR.scala 181:38:@3659.4]
  wire  _T_648; // @[CSR.scala 181:25:@3660.4]
  wire  cpu_wen; // @[CSR.scala 181:48:@3661.4]
  wire  _T_650; // @[CSR.scala 182:24:@3662.4]
  wire  wen; // @[CSR.scala 182:21:@3663.4]
  wire  _T_651; // @[Util.scala 23:47:@3664.4]
  wire  _T_652; // @[Util.scala 23:47:@3665.4]
  wire  _T_653; // @[Util.scala 23:62:@3666.4]
  wire [31:0] _T_655; // @[CSR.scala 281:9:@3667.4]
  wire [31:0] _T_656; // @[CSR.scala 281:49:@3668.4]
  wire [31:0] _T_659; // @[CSR.scala 281:64:@3670.4]
  wire [31:0] _T_660; // @[CSR.scala 281:60:@3671.4]
  wire [31:0] wdata; // @[CSR.scala 281:58:@3672.4]
  wire [2:0] _T_662; // @[CSR.scala 185:33:@3673.4]
  wire [7:0] opcode; // @[CSR.scala 185:20:@3674.4]
  wire  _T_663; // @[CSR.scala 186:40:@3675.4]
  wire  insn_call; // @[CSR.scala 186:31:@3676.4]
  wire  _T_664; // @[CSR.scala 187:41:@3677.4]
  wire  insn_break; // @[CSR.scala 187:32:@3678.4]
  wire  _T_665; // @[CSR.scala 188:39:@3679.4]
  wire  _T_666; // @[CSR.scala 188:30:@3680.4]
  wire  insn_ret; // @[CSR.scala 188:43:@3681.4]
  wire  _T_940; // @[CSR.scala 199:24:@3880.4]
  wire [1:0] _T_942; // @[Bitwise.scala 48:55:@3883.4]
  wire  _T_944; // @[CSR.scala 201:50:@3884.4]
  wire  _T_946; // @[CSR.scala 201:9:@3886.4]
  wire  _T_948; // @[CSR.scala 201:9:@3887.4]
  wire  _T_951; // @[CSR.scala 208:32:@3896.4]
  wire  _T_953; // @[CSR.scala 208:21:@3897.4]
  wire  _T_954; // @[CSR.scala 208:18:@3898.4]
  wire  _GEN_3; // @[CSR.scala 208:38:@3899.4]
  wire  _GEN_4; // @[CSR.scala 208:38:@3899.4]
  wire [1:0] new_prv; // @[CSR.scala 208:38:@3899.4]
  wire [3:0] _GEN_148; // @[CSR.scala 218:35:@3907.6]
  wire [4:0] _T_958; // @[CSR.scala 218:35:@3907.6]
  wire [3:0] _T_959; // @[CSR.scala 218:35:@3908.6]
  wire [31:0] _GEN_7; // @[CSR.scala 216:18:@3905.4]
  wire [31:0] _GEN_8; // @[CSR.scala 216:18:@3905.4]
  wire [31:0] _GEN_9; // @[CSR.scala 216:18:@3905.4]
  wire [31:0] _GEN_10; // @[CSR.scala 223:19:@3912.4]
  wire [31:0] _GEN_11; // @[CSR.scala 223:19:@3912.4]
  wire [31:0] _GEN_12; // @[CSR.scala 223:19:@3912.4]
  wire [31:0] _GEN_14; // @[CSR.scala 229:17:@3917.4]
  wire [31:0] _GEN_15; // @[CSR.scala 229:17:@3917.4]
  wire [31:0] _GEN_16; // @[CSR.scala 229:17:@3917.4]
  wire [63:0] _T_965; // @[Mux.scala 19:72:@3925.4]
  wire [63:0] _T_967; // @[Mux.scala 19:72:@3926.4]
  wire [15:0] _T_969; // @[Mux.scala 19:72:@3927.4]
  wire [30:0] _T_975; // @[Mux.scala 19:72:@3930.4]
  wire [31:0] _T_977; // @[Mux.scala 19:72:@3931.4]
  wire [8:0] _T_979; // @[Mux.scala 19:72:@3932.4]
  wire [15:0] _T_981; // @[Mux.scala 19:72:@3933.4]
  wire [15:0] _T_983; // @[Mux.scala 19:72:@3934.4]
  wire [31:0] _T_985; // @[Mux.scala 19:72:@3935.4]
  wire [31:0] _T_987; // @[Mux.scala 19:72:@3936.4]
  wire [31:0] _T_989; // @[Mux.scala 19:72:@3937.4]
  wire [31:0] _T_991; // @[Mux.scala 19:72:@3938.4]
  wire [31:0] _T_995; // @[Mux.scala 19:72:@3940.4]
  wire [31:0] _T_997; // @[Mux.scala 19:72:@3941.4]
  wire [39:0] _T_999; // @[Mux.scala 19:72:@3942.4]
  wire [39:0] _T_1001; // @[Mux.scala 19:72:@3943.4]
  wire [39:0] _T_1003; // @[Mux.scala 19:72:@3944.4]
  wire [39:0] _T_1005; // @[Mux.scala 19:72:@3945.4]
  wire [39:0] _T_1007; // @[Mux.scala 19:72:@3946.4]
  wire [39:0] _T_1009; // @[Mux.scala 19:72:@3947.4]
  wire [39:0] _T_1011; // @[Mux.scala 19:72:@3948.4]
  wire [39:0] _T_1013; // @[Mux.scala 19:72:@3949.4]
  wire [39:0] _T_1015; // @[Mux.scala 19:72:@3950.4]
  wire [39:0] _T_1017; // @[Mux.scala 19:72:@3951.4]
  wire [39:0] _T_1019; // @[Mux.scala 19:72:@3952.4]
  wire [39:0] _T_1021; // @[Mux.scala 19:72:@3953.4]
  wire [39:0] _T_1023; // @[Mux.scala 19:72:@3954.4]
  wire [39:0] _T_1025; // @[Mux.scala 19:72:@3955.4]
  wire [39:0] _T_1027; // @[Mux.scala 19:72:@3956.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:@3957.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:@3958.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:@3959.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:@3960.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:@3961.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:@3962.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:@3963.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:@3964.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:@3965.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:@3966.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:@3967.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:@3968.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:@3969.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:@3970.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:@3971.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:@3972.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:@3973.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:@3974.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:@3975.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:@3976.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:@3977.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:@3978.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:@3979.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:@3980.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:@3981.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:@3982.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:@3983.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:@3984.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:@3985.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:@3986.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:@3987.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:@3988.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:@3989.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:@3990.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:@3991.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:@3992.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:@3993.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:@3994.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:@3995.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:@3996.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:@3997.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:@3998.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:@3999.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:@4000.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:@4001.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:@4002.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:@4003.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:@4004.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:@4005.4]
  wire [63:0] _T_1130; // @[Mux.scala 19:72:@4008.4]
  wire [63:0] _GEN_149; // @[Mux.scala 19:72:@4009.4]
  wire [63:0] _T_1131; // @[Mux.scala 19:72:@4009.4]
  wire [63:0] _GEN_150; // @[Mux.scala 19:72:@4012.4]
  wire [63:0] _T_1134; // @[Mux.scala 19:72:@4012.4]
  wire [63:0] _GEN_151; // @[Mux.scala 19:72:@4013.4]
  wire [63:0] _T_1135; // @[Mux.scala 19:72:@4013.4]
  wire [63:0] _GEN_152; // @[Mux.scala 19:72:@4014.4]
  wire [63:0] _T_1136; // @[Mux.scala 19:72:@4014.4]
  wire [63:0] _GEN_153; // @[Mux.scala 19:72:@4015.4]
  wire [63:0] _T_1137; // @[Mux.scala 19:72:@4015.4]
  wire [63:0] _GEN_154; // @[Mux.scala 19:72:@4016.4]
  wire [63:0] _T_1138; // @[Mux.scala 19:72:@4016.4]
  wire [63:0] _GEN_155; // @[Mux.scala 19:72:@4017.4]
  wire [63:0] _T_1139; // @[Mux.scala 19:72:@4017.4]
  wire [63:0] _GEN_156; // @[Mux.scala 19:72:@4018.4]
  wire [63:0] _T_1140; // @[Mux.scala 19:72:@4018.4]
  wire [63:0] _GEN_157; // @[Mux.scala 19:72:@4019.4]
  wire [63:0] _T_1141; // @[Mux.scala 19:72:@4019.4]
  wire [63:0] _GEN_158; // @[Mux.scala 19:72:@4020.4]
  wire [63:0] _T_1142; // @[Mux.scala 19:72:@4020.4]
  wire [63:0] _GEN_159; // @[Mux.scala 19:72:@4022.4]
  wire [63:0] _T_1144; // @[Mux.scala 19:72:@4022.4]
  wire [63:0] _GEN_160; // @[Mux.scala 19:72:@4023.4]
  wire [63:0] _T_1145; // @[Mux.scala 19:72:@4023.4]
  wire [63:0] _GEN_161; // @[Mux.scala 19:72:@4024.4]
  wire [63:0] _T_1146; // @[Mux.scala 19:72:@4024.4]
  wire [63:0] _GEN_162; // @[Mux.scala 19:72:@4025.4]
  wire [63:0] _T_1147; // @[Mux.scala 19:72:@4025.4]
  wire [63:0] _GEN_163; // @[Mux.scala 19:72:@4026.4]
  wire [63:0] _T_1148; // @[Mux.scala 19:72:@4026.4]
  wire [63:0] _GEN_164; // @[Mux.scala 19:72:@4027.4]
  wire [63:0] _T_1149; // @[Mux.scala 19:72:@4027.4]
  wire [63:0] _GEN_165; // @[Mux.scala 19:72:@4028.4]
  wire [63:0] _T_1150; // @[Mux.scala 19:72:@4028.4]
  wire [63:0] _GEN_166; // @[Mux.scala 19:72:@4029.4]
  wire [63:0] _T_1151; // @[Mux.scala 19:72:@4029.4]
  wire [63:0] _GEN_167; // @[Mux.scala 19:72:@4030.4]
  wire [63:0] _T_1152; // @[Mux.scala 19:72:@4030.4]
  wire [63:0] _GEN_168; // @[Mux.scala 19:72:@4031.4]
  wire [63:0] _T_1153; // @[Mux.scala 19:72:@4031.4]
  wire [63:0] _GEN_169; // @[Mux.scala 19:72:@4032.4]
  wire [63:0] _T_1154; // @[Mux.scala 19:72:@4032.4]
  wire [63:0] _GEN_170; // @[Mux.scala 19:72:@4033.4]
  wire [63:0] _T_1155; // @[Mux.scala 19:72:@4033.4]
  wire [63:0] _GEN_171; // @[Mux.scala 19:72:@4034.4]
  wire [63:0] _T_1156; // @[Mux.scala 19:72:@4034.4]
  wire [63:0] _GEN_172; // @[Mux.scala 19:72:@4035.4]
  wire [63:0] _T_1157; // @[Mux.scala 19:72:@4035.4]
  wire [63:0] _GEN_173; // @[Mux.scala 19:72:@4036.4]
  wire [63:0] _T_1158; // @[Mux.scala 19:72:@4036.4]
  wire [63:0] _GEN_174; // @[Mux.scala 19:72:@4037.4]
  wire [63:0] _T_1159; // @[Mux.scala 19:72:@4037.4]
  wire [63:0] _GEN_175; // @[Mux.scala 19:72:@4038.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:@4038.4]
  wire [63:0] _GEN_176; // @[Mux.scala 19:72:@4039.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:@4039.4]
  wire [63:0] _GEN_177; // @[Mux.scala 19:72:@4040.4]
  wire [63:0] _T_1162; // @[Mux.scala 19:72:@4040.4]
  wire [63:0] _GEN_178; // @[Mux.scala 19:72:@4041.4]
  wire [63:0] _T_1163; // @[Mux.scala 19:72:@4041.4]
  wire [63:0] _GEN_179; // @[Mux.scala 19:72:@4042.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:@4042.4]
  wire [63:0] _GEN_180; // @[Mux.scala 19:72:@4043.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:@4043.4]
  wire [63:0] _GEN_181; // @[Mux.scala 19:72:@4044.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:@4044.4]
  wire [63:0] _GEN_182; // @[Mux.scala 19:72:@4045.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:@4045.4]
  wire [63:0] _GEN_183; // @[Mux.scala 19:72:@4046.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:@4046.4]
  wire [63:0] _GEN_184; // @[Mux.scala 19:72:@4047.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:@4047.4]
  wire [63:0] _GEN_185; // @[Mux.scala 19:72:@4048.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:@4048.4]
  wire [63:0] _GEN_186; // @[Mux.scala 19:72:@4049.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:@4049.4]
  wire [63:0] _GEN_187; // @[Mux.scala 19:72:@4050.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:@4050.4]
  wire [63:0] _GEN_188; // @[Mux.scala 19:72:@4051.4]
  wire [63:0] _T_1173; // @[Mux.scala 19:72:@4051.4]
  wire [63:0] _GEN_189; // @[Mux.scala 19:72:@4052.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:@4052.4]
  wire [63:0] _GEN_190; // @[Mux.scala 19:72:@4053.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:@4053.4]
  wire [63:0] _GEN_191; // @[Mux.scala 19:72:@4054.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:@4054.4]
  wire [63:0] _GEN_192; // @[Mux.scala 19:72:@4055.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:@4055.4]
  wire [63:0] _GEN_193; // @[Mux.scala 19:72:@4056.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:@4056.4]
  wire [63:0] _GEN_194; // @[Mux.scala 19:72:@4057.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:@4057.4]
  wire [63:0] _GEN_195; // @[Mux.scala 19:72:@4058.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:@4058.4]
  wire [63:0] _GEN_196; // @[Mux.scala 19:72:@4059.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:@4059.4]
  wire [63:0] _GEN_197; // @[Mux.scala 19:72:@4060.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:@4060.4]
  wire [63:0] _GEN_198; // @[Mux.scala 19:72:@4061.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:@4061.4]
  wire [63:0] _GEN_199; // @[Mux.scala 19:72:@4062.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:@4062.4]
  wire [63:0] _GEN_200; // @[Mux.scala 19:72:@4063.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:@4063.4]
  wire [63:0] _GEN_201; // @[Mux.scala 19:72:@4064.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:@4064.4]
  wire [63:0] _GEN_202; // @[Mux.scala 19:72:@4065.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:@4065.4]
  wire [63:0] _GEN_203; // @[Mux.scala 19:72:@4066.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:@4066.4]
  wire [63:0] _GEN_204; // @[Mux.scala 19:72:@4067.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:@4067.4]
  wire [63:0] _GEN_205; // @[Mux.scala 19:72:@4068.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:@4068.4]
  wire [63:0] _GEN_206; // @[Mux.scala 19:72:@4069.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:@4069.4]
  wire [63:0] _GEN_207; // @[Mux.scala 19:72:@4070.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:@4070.4]
  wire [63:0] _GEN_208; // @[Mux.scala 19:72:@4071.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:@4071.4]
  wire [63:0] _GEN_209; // @[Mux.scala 19:72:@4072.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:@4072.4]
  wire [63:0] _GEN_210; // @[Mux.scala 19:72:@4073.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:@4073.4]
  wire [63:0] _GEN_211; // @[Mux.scala 19:72:@4074.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:@4074.4]
  wire [63:0] _GEN_212; // @[Mux.scala 19:72:@4075.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:@4075.4]
  wire [63:0] _GEN_213; // @[Mux.scala 19:72:@4076.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:@4076.4]
  wire [63:0] _GEN_214; // @[Mux.scala 19:72:@4077.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:@4077.4]
  wire [63:0] _GEN_215; // @[Mux.scala 19:72:@4078.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:@4078.4]
  wire [63:0] _GEN_216; // @[Mux.scala 19:72:@4079.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:@4079.4]
  wire [63:0] _GEN_217; // @[Mux.scala 19:72:@4080.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:@4080.4]
  wire [63:0] _GEN_218; // @[Mux.scala 19:72:@4081.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:@4081.4]
  wire [63:0] _GEN_219; // @[Mux.scala 19:72:@4082.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:@4082.4]
  wire [63:0] _GEN_220; // @[Mux.scala 19:72:@4083.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:@4083.4]
  wire [63:0] _GEN_221; // @[Mux.scala 19:72:@4084.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:@4084.4]
  wire [63:0] _GEN_222; // @[Mux.scala 19:72:@4085.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:@4085.4]
  wire [63:0] _GEN_223; // @[Mux.scala 19:72:@4086.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:@4086.4]
  wire [63:0] _GEN_224; // @[Mux.scala 19:72:@4087.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:@4087.4]
  wire  _T_1220; // @[CSR.scala 245:39:@4100.8]
  wire  _T_1222; // @[CSR.scala 245:39:@4104.8]
  wire  _GEN_17; // @[CSR.scala 244:39:@4094.6]
  wire  _GEN_18; // @[CSR.scala 244:39:@4094.6]
  wire [15:0] _T_1233; // @[:@4123.8 :@4124.8]
  wire  _T_1235; // @[CSR.scala 250:35:@4127.8]
  wire  _T_1237; // @[CSR.scala 250:35:@4131.8]
  wire  _GEN_19; // @[CSR.scala 249:35:@4121.6]
  wire  _GEN_20; // @[CSR.scala 253:35:@4141.6]
  wire  _GEN_21; // @[CSR.scala 253:35:@4141.6]
  wire [7:0] _T_1253; // @[CSR.scala 277:47:@4163.8]
  wire [31:0] _T_1254; // @[CSR.scala 277:72:@4164.8]
  wire [39:0] _T_1255; // @[Cat.scala 30:58:@4165.8]
  wire [40:0] _GEN_22; // @[CSR.scala 277:29:@4162.6]
  wire [7:0] _T_1256; // @[CSR.scala 278:45:@4169.8]
  wire [39:0] _T_1257; // @[Cat.scala 30:58:@4170.8]
  wire [40:0] _GEN_23; // @[CSR.scala 278:29:@4168.6]
  wire [31:0] _T_1259; // @[CSR.scala 277:72:@4175.8]
  wire [39:0] _T_1260; // @[Cat.scala 30:58:@4176.8]
  wire [40:0] _GEN_24; // @[CSR.scala 277:29:@4173.6]
  wire [7:0] _T_1261; // @[CSR.scala 278:45:@4180.8]
  wire [39:0] _T_1262; // @[Cat.scala 30:58:@4181.8]
  wire [40:0] _GEN_25; // @[CSR.scala 278:29:@4179.6]
  wire [31:0] _T_1264; // @[CSR.scala 277:72:@4186.8]
  wire [39:0] _T_1265; // @[Cat.scala 30:58:@4187.8]
  wire [40:0] _GEN_26; // @[CSR.scala 277:29:@4184.6]
  wire [7:0] _T_1266; // @[CSR.scala 278:45:@4191.8]
  wire [39:0] _T_1267; // @[Cat.scala 30:58:@4192.8]
  wire [40:0] _GEN_27; // @[CSR.scala 278:29:@4190.6]
  wire [31:0] _T_1269; // @[CSR.scala 277:72:@4197.8]
  wire [39:0] _T_1270; // @[Cat.scala 30:58:@4198.8]
  wire [40:0] _GEN_28; // @[CSR.scala 277:29:@4195.6]
  wire [7:0] _T_1271; // @[CSR.scala 278:45:@4202.8]
  wire [39:0] _T_1272; // @[Cat.scala 30:58:@4203.8]
  wire [40:0] _GEN_29; // @[CSR.scala 278:29:@4201.6]
  wire [31:0] _T_1274; // @[CSR.scala 277:72:@4208.8]
  wire [39:0] _T_1275; // @[Cat.scala 30:58:@4209.8]
  wire [40:0] _GEN_30; // @[CSR.scala 277:29:@4206.6]
  wire [7:0] _T_1276; // @[CSR.scala 278:45:@4213.8]
  wire [39:0] _T_1277; // @[Cat.scala 30:58:@4214.8]
  wire [40:0] _GEN_31; // @[CSR.scala 278:29:@4212.6]
  wire [31:0] _T_1279; // @[CSR.scala 277:72:@4219.8]
  wire [39:0] _T_1280; // @[Cat.scala 30:58:@4220.8]
  wire [40:0] _GEN_32; // @[CSR.scala 277:29:@4217.6]
  wire [7:0] _T_1281; // @[CSR.scala 278:45:@4224.8]
  wire [39:0] _T_1282; // @[Cat.scala 30:58:@4225.8]
  wire [40:0] _GEN_33; // @[CSR.scala 278:29:@4223.6]
  wire [31:0] _T_1284; // @[CSR.scala 277:72:@4230.8]
  wire [39:0] _T_1285; // @[Cat.scala 30:58:@4231.8]
  wire [40:0] _GEN_34; // @[CSR.scala 277:29:@4228.6]
  wire [7:0] _T_1286; // @[CSR.scala 278:45:@4235.8]
  wire [39:0] _T_1287; // @[Cat.scala 30:58:@4236.8]
  wire [40:0] _GEN_35; // @[CSR.scala 278:29:@4234.6]
  wire [31:0] _T_1289; // @[CSR.scala 277:72:@4241.8]
  wire [39:0] _T_1290; // @[Cat.scala 30:58:@4242.8]
  wire [40:0] _GEN_36; // @[CSR.scala 277:29:@4239.6]
  wire [7:0] _T_1291; // @[CSR.scala 278:45:@4246.8]
  wire [39:0] _T_1292; // @[Cat.scala 30:58:@4247.8]
  wire [40:0] _GEN_37; // @[CSR.scala 278:29:@4245.6]
  wire [31:0] _T_1294; // @[CSR.scala 277:72:@4252.8]
  wire [39:0] _T_1295; // @[Cat.scala 30:58:@4253.8]
  wire [40:0] _GEN_38; // @[CSR.scala 277:29:@4250.6]
  wire [7:0] _T_1296; // @[CSR.scala 278:45:@4257.8]
  wire [39:0] _T_1297; // @[Cat.scala 30:58:@4258.8]
  wire [40:0] _GEN_39; // @[CSR.scala 278:29:@4256.6]
  wire [31:0] _T_1299; // @[CSR.scala 277:72:@4263.8]
  wire [39:0] _T_1300; // @[Cat.scala 30:58:@4264.8]
  wire [40:0] _GEN_40; // @[CSR.scala 277:29:@4261.6]
  wire [7:0] _T_1301; // @[CSR.scala 278:45:@4268.8]
  wire [39:0] _T_1302; // @[Cat.scala 30:58:@4269.8]
  wire [40:0] _GEN_41; // @[CSR.scala 278:29:@4267.6]
  wire [31:0] _T_1304; // @[CSR.scala 277:72:@4274.8]
  wire [39:0] _T_1305; // @[Cat.scala 30:58:@4275.8]
  wire [40:0] _GEN_42; // @[CSR.scala 277:29:@4272.6]
  wire [7:0] _T_1306; // @[CSR.scala 278:45:@4279.8]
  wire [39:0] _T_1307; // @[Cat.scala 30:58:@4280.8]
  wire [40:0] _GEN_43; // @[CSR.scala 278:29:@4278.6]
  wire [31:0] _T_1309; // @[CSR.scala 277:72:@4285.8]
  wire [39:0] _T_1310; // @[Cat.scala 30:58:@4286.8]
  wire [40:0] _GEN_44; // @[CSR.scala 277:29:@4283.6]
  wire [7:0] _T_1311; // @[CSR.scala 278:45:@4290.8]
  wire [39:0] _T_1312; // @[Cat.scala 30:58:@4291.8]
  wire [40:0] _GEN_45; // @[CSR.scala 278:29:@4289.6]
  wire [31:0] _T_1314; // @[CSR.scala 277:72:@4296.8]
  wire [39:0] _T_1315; // @[Cat.scala 30:58:@4297.8]
  wire [40:0] _GEN_46; // @[CSR.scala 277:29:@4294.6]
  wire [7:0] _T_1316; // @[CSR.scala 278:45:@4301.8]
  wire [39:0] _T_1317; // @[Cat.scala 30:58:@4302.8]
  wire [40:0] _GEN_47; // @[CSR.scala 278:29:@4300.6]
  wire [31:0] _T_1319; // @[CSR.scala 277:72:@4307.8]
  wire [39:0] _T_1320; // @[Cat.scala 30:58:@4308.8]
  wire [40:0] _GEN_48; // @[CSR.scala 277:29:@4305.6]
  wire [7:0] _T_1321; // @[CSR.scala 278:45:@4312.8]
  wire [39:0] _T_1322; // @[Cat.scala 30:58:@4313.8]
  wire [40:0] _GEN_49; // @[CSR.scala 278:29:@4311.6]
  wire [31:0] _T_1324; // @[CSR.scala 277:72:@4318.8]
  wire [39:0] _T_1325; // @[Cat.scala 30:58:@4319.8]
  wire [40:0] _GEN_50; // @[CSR.scala 277:29:@4316.6]
  wire [7:0] _T_1326; // @[CSR.scala 278:45:@4323.8]
  wire [39:0] _T_1327; // @[Cat.scala 30:58:@4324.8]
  wire [40:0] _GEN_51; // @[CSR.scala 278:29:@4322.6]
  wire [31:0] _T_1329; // @[CSR.scala 277:72:@4329.8]
  wire [39:0] _T_1330; // @[Cat.scala 30:58:@4330.8]
  wire [40:0] _GEN_52; // @[CSR.scala 277:29:@4327.6]
  wire [7:0] _T_1331; // @[CSR.scala 278:45:@4334.8]
  wire [39:0] _T_1332; // @[Cat.scala 30:58:@4335.8]
  wire [40:0] _GEN_53; // @[CSR.scala 278:29:@4333.6]
  wire [31:0] _T_1334; // @[CSR.scala 277:72:@4340.8]
  wire [39:0] _T_1335; // @[Cat.scala 30:58:@4341.8]
  wire [40:0] _GEN_54; // @[CSR.scala 277:29:@4338.6]
  wire [7:0] _T_1336; // @[CSR.scala 278:45:@4345.8]
  wire [39:0] _T_1337; // @[Cat.scala 30:58:@4346.8]
  wire [40:0] _GEN_55; // @[CSR.scala 278:29:@4344.6]
  wire [31:0] _T_1339; // @[CSR.scala 277:72:@4351.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:@4352.8]
  wire [40:0] _GEN_56; // @[CSR.scala 277:29:@4349.6]
  wire [7:0] _T_1341; // @[CSR.scala 278:45:@4356.8]
  wire [39:0] _T_1342; // @[Cat.scala 30:58:@4357.8]
  wire [40:0] _GEN_57; // @[CSR.scala 278:29:@4355.6]
  wire [31:0] _T_1344; // @[CSR.scala 277:72:@4362.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:@4363.8]
  wire [40:0] _GEN_58; // @[CSR.scala 277:29:@4360.6]
  wire [7:0] _T_1346; // @[CSR.scala 278:45:@4367.8]
  wire [39:0] _T_1347; // @[Cat.scala 30:58:@4368.8]
  wire [40:0] _GEN_59; // @[CSR.scala 278:29:@4366.6]
  wire [31:0] _T_1349; // @[CSR.scala 277:72:@4373.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:@4374.8]
  wire [40:0] _GEN_60; // @[CSR.scala 277:29:@4371.6]
  wire [7:0] _T_1351; // @[CSR.scala 278:45:@4378.8]
  wire [39:0] _T_1352; // @[Cat.scala 30:58:@4379.8]
  wire [40:0] _GEN_61; // @[CSR.scala 278:29:@4377.6]
  wire [31:0] _T_1354; // @[CSR.scala 277:72:@4384.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:@4385.8]
  wire [40:0] _GEN_62; // @[CSR.scala 277:29:@4382.6]
  wire [7:0] _T_1356; // @[CSR.scala 278:45:@4389.8]
  wire [39:0] _T_1357; // @[Cat.scala 30:58:@4390.8]
  wire [40:0] _GEN_63; // @[CSR.scala 278:29:@4388.6]
  wire [31:0] _T_1359; // @[CSR.scala 277:72:@4395.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:@4396.8]
  wire [40:0] _GEN_64; // @[CSR.scala 277:29:@4393.6]
  wire [7:0] _T_1361; // @[CSR.scala 278:45:@4400.8]
  wire [39:0] _T_1362; // @[Cat.scala 30:58:@4401.8]
  wire [40:0] _GEN_65; // @[CSR.scala 278:29:@4399.6]
  wire [31:0] _T_1364; // @[CSR.scala 277:72:@4406.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:@4407.8]
  wire [40:0] _GEN_66; // @[CSR.scala 277:29:@4404.6]
  wire [7:0] _T_1366; // @[CSR.scala 278:45:@4411.8]
  wire [39:0] _T_1367; // @[Cat.scala 30:58:@4412.8]
  wire [40:0] _GEN_67; // @[CSR.scala 278:29:@4410.6]
  wire [31:0] _T_1369; // @[CSR.scala 277:72:@4417.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:@4418.8]
  wire [40:0] _GEN_68; // @[CSR.scala 277:29:@4415.6]
  wire [7:0] _T_1371; // @[CSR.scala 278:45:@4422.8]
  wire [39:0] _T_1372; // @[Cat.scala 30:58:@4423.8]
  wire [40:0] _GEN_69; // @[CSR.scala 278:29:@4421.6]
  wire [31:0] _T_1374; // @[CSR.scala 277:72:@4428.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:@4429.8]
  wire [40:0] _GEN_70; // @[CSR.scala 277:29:@4426.6]
  wire [7:0] _T_1376; // @[CSR.scala 278:45:@4433.8]
  wire [39:0] _T_1377; // @[Cat.scala 30:58:@4434.8]
  wire [40:0] _GEN_71; // @[CSR.scala 278:29:@4432.6]
  wire [31:0] _T_1379; // @[CSR.scala 277:72:@4439.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:@4440.8]
  wire [40:0] _GEN_72; // @[CSR.scala 277:29:@4437.6]
  wire [7:0] _T_1381; // @[CSR.scala 278:45:@4444.8]
  wire [39:0] _T_1382; // @[Cat.scala 30:58:@4445.8]
  wire [40:0] _GEN_73; // @[CSR.scala 278:29:@4443.6]
  wire [31:0] _T_1384; // @[CSR.scala 277:72:@4450.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:@4451.8]
  wire [40:0] _GEN_74; // @[CSR.scala 277:29:@4448.6]
  wire [7:0] _T_1386; // @[CSR.scala 278:45:@4455.8]
  wire [39:0] _T_1387; // @[Cat.scala 30:58:@4456.8]
  wire [40:0] _GEN_75; // @[CSR.scala 278:29:@4454.6]
  wire [31:0] _T_1389; // @[CSR.scala 277:72:@4461.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:@4462.8]
  wire [40:0] _GEN_76; // @[CSR.scala 277:29:@4459.6]
  wire [7:0] _T_1391; // @[CSR.scala 278:45:@4466.8]
  wire [39:0] _T_1392; // @[Cat.scala 30:58:@4467.8]
  wire [40:0] _GEN_77; // @[CSR.scala 278:29:@4465.6]
  wire [31:0] _T_1394; // @[CSR.scala 277:72:@4472.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:@4473.8]
  wire [40:0] _GEN_78; // @[CSR.scala 277:29:@4470.6]
  wire [7:0] _T_1396; // @[CSR.scala 278:45:@4477.8]
  wire [39:0] _T_1397; // @[Cat.scala 30:58:@4478.8]
  wire [40:0] _GEN_79; // @[CSR.scala 278:29:@4476.6]
  wire [31:0] _T_1399; // @[CSR.scala 277:72:@4483.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:@4484.8]
  wire [40:0] _GEN_80; // @[CSR.scala 277:29:@4481.6]
  wire [7:0] _T_1401; // @[CSR.scala 278:45:@4488.8]
  wire [39:0] _T_1402; // @[Cat.scala 30:58:@4489.8]
  wire [40:0] _GEN_81; // @[CSR.scala 278:29:@4487.6]
  wire [31:0] _T_1404; // @[CSR.scala 277:72:@4494.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:@4495.8]
  wire [40:0] _GEN_82; // @[CSR.scala 277:29:@4492.6]
  wire [7:0] _T_1406; // @[CSR.scala 278:45:@4499.8]
  wire [39:0] _T_1407; // @[Cat.scala 30:58:@4500.8]
  wire [40:0] _GEN_83; // @[CSR.scala 278:29:@4498.6]
  wire [31:0] _T_1409; // @[CSR.scala 277:72:@4505.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:@4506.8]
  wire [40:0] _GEN_84; // @[CSR.scala 277:29:@4503.6]
  wire [7:0] _T_1411; // @[CSR.scala 278:45:@4510.8]
  wire [39:0] _T_1412; // @[Cat.scala 30:58:@4511.8]
  wire [40:0] _GEN_85; // @[CSR.scala 278:29:@4509.6]
  wire [31:0] _T_1414; // @[CSR.scala 277:72:@4516.8]
  wire [63:0] _T_1415; // @[Cat.scala 30:58:@4517.8]
  wire [57:0] _T_1416; // @[Util.scala 133:28:@4519.8]
  wire [63:0] _GEN_86; // @[CSR.scala 277:29:@4514.6]
  wire [57:0] _GEN_87; // @[CSR.scala 277:29:@4514.6]
  wire [31:0] _T_1417; // @[CSR.scala 278:45:@4523.8]
  wire [63:0] _T_1418; // @[Cat.scala 30:58:@4524.8]
  wire [57:0] _T_1419; // @[Util.scala 133:28:@4526.8]
  wire [63:0] _GEN_88; // @[CSR.scala 278:29:@4522.6]
  wire [57:0] _GEN_89; // @[CSR.scala 278:29:@4522.6]
  wire [31:0] _T_1421; // @[CSR.scala 277:72:@4531.8]
  wire [63:0] _T_1422; // @[Cat.scala 30:58:@4532.8]
  wire [57:0] _T_1423; // @[Util.scala 133:28:@4534.8]
  wire [63:0] _GEN_90; // @[CSR.scala 277:29:@4529.6]
  wire [57:0] _GEN_91; // @[CSR.scala 277:29:@4529.6]
  wire [31:0] _T_1424; // @[CSR.scala 278:45:@4538.8]
  wire [63:0] _T_1425; // @[Cat.scala 30:58:@4539.8]
  wire [57:0] _T_1426; // @[Util.scala 133:28:@4541.8]
  wire [63:0] _GEN_92; // @[CSR.scala 278:29:@4537.6]
  wire [57:0] _GEN_93; // @[CSR.scala 278:29:@4537.6]
  wire [31:0] _GEN_94; // @[CSR.scala 265:40:@4544.6]
  wire [31:0] _T_1429; // @[CSR.scala 267:78:@4549.8]
  wire [34:0] _GEN_225; // @[CSR.scala 267:86:@4550.8]
  wire [34:0] _T_1431; // @[CSR.scala 267:86:@4550.8]
  wire [34:0] _GEN_95; // @[CSR.scala 267:40:@4547.6]
  wire [31:0] _GEN_96; // @[CSR.scala 268:40:@4553.6]
  wire [31:0] _T_1433; // @[CSR.scala 269:62:@4557.8]
  wire [31:0] _GEN_97; // @[CSR.scala 269:40:@4556.6]
  wire [31:0] _GEN_98; // @[CSR.scala 270:40:@4560.6]
  wire [31:0] _GEN_99; // @[CSR.scala 271:42:@4564.6]
  wire  _GEN_100; // @[CSR.scala 242:14:@4093.4]
  wire  _GEN_101; // @[CSR.scala 242:14:@4093.4]
  wire  _GEN_102; // @[CSR.scala 242:14:@4093.4]
  wire  _GEN_103; // @[CSR.scala 242:14:@4093.4]
  wire  _GEN_104; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_105; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_106; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_107; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_108; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_109; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_110; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_111; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_112; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_113; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_114; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_115; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_116; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_117; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_118; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_119; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_120; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_121; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_122; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_123; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_124; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_125; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_126; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_127; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_128; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_129; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_130; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_131; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_132; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_133; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_134; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_135; // @[CSR.scala 242:14:@4093.4]
  wire [40:0] _GEN_136; // @[CSR.scala 242:14:@4093.4]
  wire [63:0] _GEN_137; // @[CSR.scala 242:14:@4093.4]
  wire [57:0] _GEN_138; // @[CSR.scala 242:14:@4093.4]
  wire [63:0] _GEN_139; // @[CSR.scala 242:14:@4093.4]
  wire [57:0] _GEN_140; // @[CSR.scala 242:14:@4093.4]
  wire [34:0] _GEN_142; // @[CSR.scala 242:14:@4093.4]
  assign _T_241 = _T_240 + 6'h1; // @[Util.scala 113:33:@3339.4]
  assign _T_245 = _T_241[6]; // @[Util.scala 118:20:@3342.4]
  assign _T_247 = _T_244 + 58'h1; // @[Util.scala 118:43:@3344.6]
  assign _T_248 = _T_244 + 58'h1; // @[Util.scala 118:43:@3345.6]
  assign _GEN_0 = _T_245 ? _T_248 : _T_244; // @[Util.scala 118:34:@3343.4]
  assign _T_249 = {_T_244,_T_240}; // @[Cat.scala 30:58:@3348.4]
  assign _GEN_147 = {{4'd0}, io_retire}; // @[Util.scala 113:33:@3350.4]
  assign _T_253 = _T_252 + _GEN_147; // @[Util.scala 113:33:@3350.4]
  assign _T_257 = _T_253[6]; // @[Util.scala 118:20:@3353.4]
  assign _T_259 = _T_256 + 58'h1; // @[Util.scala 118:43:@3355.6]
  assign _T_260 = _T_256 + 58'h1; // @[Util.scala 118:43:@3356.6]
  assign _GEN_1 = _T_257 ? _T_260 : _T_256; // @[Util.scala 118:34:@3354.4]
  assign _T_261 = {_T_256,_T_252}; // @[Cat.scala 30:58:@3359.4]
  assign _T_265 = {{1'd0}, _T_264}; // @[Util.scala 113:33:@3362.4]
  assign _T_268 = {{1'd0}, _T_267}; // @[Util.scala 113:33:@3365.4]
  assign _T_271 = {{1'd0}, _T_270}; // @[Util.scala 113:33:@3368.4]
  assign _T_274 = {{1'd0}, _T_273}; // @[Util.scala 113:33:@3371.4]
  assign _T_277 = {{1'd0}, _T_276}; // @[Util.scala 113:33:@3374.4]
  assign _T_280 = {{1'd0}, _T_279}; // @[Util.scala 113:33:@3377.4]
  assign _T_283 = {{1'd0}, _T_282}; // @[Util.scala 113:33:@3380.4]
  assign _T_286 = {{1'd0}, _T_285}; // @[Util.scala 113:33:@3383.4]
  assign _T_289 = {{1'd0}, _T_288}; // @[Util.scala 113:33:@3386.4]
  assign _T_292 = {{1'd0}, _T_291}; // @[Util.scala 113:33:@3389.4]
  assign _T_295 = {{1'd0}, _T_294}; // @[Util.scala 113:33:@3392.4]
  assign _T_298 = {{1'd0}, _T_297}; // @[Util.scala 113:33:@3395.4]
  assign _T_301 = {{1'd0}, _T_300}; // @[Util.scala 113:33:@3398.4]
  assign _T_304 = {{1'd0}, _T_303}; // @[Util.scala 113:33:@3401.4]
  assign _T_307 = {{1'd0}, _T_306}; // @[Util.scala 113:33:@3404.4]
  assign _T_310 = {{1'd0}, _T_309}; // @[Util.scala 113:33:@3407.4]
  assign _T_313 = {{1'd0}, _T_312}; // @[Util.scala 113:33:@3410.4]
  assign _T_316 = {{1'd0}, _T_315}; // @[Util.scala 113:33:@3413.4]
  assign _T_319 = {{1'd0}, _T_318}; // @[Util.scala 113:33:@3416.4]
  assign _T_322 = {{1'd0}, _T_321}; // @[Util.scala 113:33:@3419.4]
  assign _T_325 = {{1'd0}, _T_324}; // @[Util.scala 113:33:@3422.4]
  assign _T_328 = {{1'd0}, _T_327}; // @[Util.scala 113:33:@3425.4]
  assign _T_331 = {{1'd0}, _T_330}; // @[Util.scala 113:33:@3428.4]
  assign _T_334 = {{1'd0}, _T_333}; // @[Util.scala 113:33:@3431.4]
  assign _T_337 = {{1'd0}, _T_336}; // @[Util.scala 113:33:@3434.4]
  assign _T_340 = {{1'd0}, _T_339}; // @[Util.scala 113:33:@3437.4]
  assign _T_343 = {{1'd0}, _T_342}; // @[Util.scala 113:33:@3440.4]
  assign _T_346 = {{1'd0}, _T_345}; // @[Util.scala 113:33:@3443.4]
  assign _T_349 = {{1'd0}, _T_348}; // @[Util.scala 113:33:@3446.4]
  assign _T_352 = {{1'd0}, _T_351}; // @[Util.scala 113:33:@3449.4]
  assign _T_355 = {{1'd0}, _T_354}; // @[Util.scala 113:33:@3452.4]
  assign _T_358 = {{1'd0}, _T_357}; // @[Util.scala 113:33:@3455.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 137:31:@3546.4]
  assign _T_446 = io_rw_cmd != 3'h0; // @[CSR.scala 138:27:@3547.4]
  assign _T_448 = system_insn == 1'h0; // @[CSR.scala 138:40:@3548.4]
  assign cpu_ren = _T_446 & _T_448; // @[CSR.scala 138:37:@3549.4]
  assign read_mstatus = {io_status_prv,io_status_unimp5,io_status_mprv,io_status_unimp4,io_status_mpp,io_status_unimp3,io_status_mpie,io_status_unimp2,io_status_mie,io_status_unimp1}; // @[CSR.scala 140:32:@3558.4]
  assign _T_468 = {5'h0,3'h0,reg_mip_mtip,3'h0,reg_mip_msip,3'h0}; // @[CSR.scala 156:25:@3564.4]
  assign _T_474 = {5'h0,3'h0,reg_mie_mtip,3'h0,reg_mie_msip,3'h0}; // @[CSR.scala 157:25:@3570.4]
  assign _T_478 = io_rw_addr == 12'hb00; // @[CSR.scala 177:73:@3571.4]
  assign _T_480 = io_rw_addr == 12'hb02; // @[CSR.scala 177:73:@3572.4]
  assign _T_482 = io_rw_addr == 12'hf13; // @[CSR.scala 177:73:@3573.4]
  assign _T_488 = io_rw_addr == 12'h301; // @[CSR.scala 177:73:@3576.4]
  assign _T_490 = io_rw_addr == 12'h300; // @[CSR.scala 177:73:@3577.4]
  assign _T_492 = io_rw_addr == 12'h305; // @[CSR.scala 177:73:@3578.4]
  assign _T_494 = io_rw_addr == 12'h344; // @[CSR.scala 177:73:@3579.4]
  assign _T_496 = io_rw_addr == 12'h304; // @[CSR.scala 177:73:@3580.4]
  assign _T_498 = io_rw_addr == 12'h340; // @[CSR.scala 177:73:@3581.4]
  assign _T_500 = io_rw_addr == 12'h341; // @[CSR.scala 177:73:@3582.4]
  assign _T_502 = io_rw_addr == 12'h343; // @[CSR.scala 177:73:@3583.4]
  assign _T_504 = io_rw_addr == 12'h342; // @[CSR.scala 177:73:@3584.4]
  assign _T_508 = io_rw_addr == 12'h7b2; // @[CSR.scala 177:73:@3586.4]
  assign _T_510 = io_rw_addr == 12'h302; // @[CSR.scala 177:73:@3587.4]
  assign _T_512 = io_rw_addr == 12'hb03; // @[CSR.scala 177:73:@3588.4]
  assign _T_514 = io_rw_addr == 12'hb83; // @[CSR.scala 177:73:@3589.4]
  assign _T_516 = io_rw_addr == 12'hb04; // @[CSR.scala 177:73:@3590.4]
  assign _T_518 = io_rw_addr == 12'hb84; // @[CSR.scala 177:73:@3591.4]
  assign _T_520 = io_rw_addr == 12'hb05; // @[CSR.scala 177:73:@3592.4]
  assign _T_522 = io_rw_addr == 12'hb85; // @[CSR.scala 177:73:@3593.4]
  assign _T_524 = io_rw_addr == 12'hb06; // @[CSR.scala 177:73:@3594.4]
  assign _T_526 = io_rw_addr == 12'hb86; // @[CSR.scala 177:73:@3595.4]
  assign _T_528 = io_rw_addr == 12'hb07; // @[CSR.scala 177:73:@3596.4]
  assign _T_530 = io_rw_addr == 12'hb87; // @[CSR.scala 177:73:@3597.4]
  assign _T_532 = io_rw_addr == 12'hb08; // @[CSR.scala 177:73:@3598.4]
  assign _T_534 = io_rw_addr == 12'hb88; // @[CSR.scala 177:73:@3599.4]
  assign _T_536 = io_rw_addr == 12'hb09; // @[CSR.scala 177:73:@3600.4]
  assign _T_538 = io_rw_addr == 12'hb89; // @[CSR.scala 177:73:@3601.4]
  assign _T_540 = io_rw_addr == 12'hb0a; // @[CSR.scala 177:73:@3602.4]
  assign _T_542 = io_rw_addr == 12'hb8a; // @[CSR.scala 177:73:@3603.4]
  assign _T_544 = io_rw_addr == 12'hb0b; // @[CSR.scala 177:73:@3604.4]
  assign _T_546 = io_rw_addr == 12'hb8b; // @[CSR.scala 177:73:@3605.4]
  assign _T_548 = io_rw_addr == 12'hb0c; // @[CSR.scala 177:73:@3606.4]
  assign _T_550 = io_rw_addr == 12'hb8c; // @[CSR.scala 177:73:@3607.4]
  assign _T_552 = io_rw_addr == 12'hb0d; // @[CSR.scala 177:73:@3608.4]
  assign _T_554 = io_rw_addr == 12'hb8d; // @[CSR.scala 177:73:@3609.4]
  assign _T_556 = io_rw_addr == 12'hb0e; // @[CSR.scala 177:73:@3610.4]
  assign _T_558 = io_rw_addr == 12'hb8e; // @[CSR.scala 177:73:@3611.4]
  assign _T_560 = io_rw_addr == 12'hb0f; // @[CSR.scala 177:73:@3612.4]
  assign _T_562 = io_rw_addr == 12'hb8f; // @[CSR.scala 177:73:@3613.4]
  assign _T_564 = io_rw_addr == 12'hb10; // @[CSR.scala 177:73:@3614.4]
  assign _T_566 = io_rw_addr == 12'hb90; // @[CSR.scala 177:73:@3615.4]
  assign _T_568 = io_rw_addr == 12'hb11; // @[CSR.scala 177:73:@3616.4]
  assign _T_570 = io_rw_addr == 12'hb91; // @[CSR.scala 177:73:@3617.4]
  assign _T_572 = io_rw_addr == 12'hb12; // @[CSR.scala 177:73:@3618.4]
  assign _T_574 = io_rw_addr == 12'hb92; // @[CSR.scala 177:73:@3619.4]
  assign _T_576 = io_rw_addr == 12'hb13; // @[CSR.scala 177:73:@3620.4]
  assign _T_578 = io_rw_addr == 12'hb93; // @[CSR.scala 177:73:@3621.4]
  assign _T_580 = io_rw_addr == 12'hb14; // @[CSR.scala 177:73:@3622.4]
  assign _T_582 = io_rw_addr == 12'hb94; // @[CSR.scala 177:73:@3623.4]
  assign _T_584 = io_rw_addr == 12'hb15; // @[CSR.scala 177:73:@3624.4]
  assign _T_586 = io_rw_addr == 12'hb95; // @[CSR.scala 177:73:@3625.4]
  assign _T_588 = io_rw_addr == 12'hb16; // @[CSR.scala 177:73:@3626.4]
  assign _T_590 = io_rw_addr == 12'hb96; // @[CSR.scala 177:73:@3627.4]
  assign _T_592 = io_rw_addr == 12'hb17; // @[CSR.scala 177:73:@3628.4]
  assign _T_594 = io_rw_addr == 12'hb97; // @[CSR.scala 177:73:@3629.4]
  assign _T_596 = io_rw_addr == 12'hb18; // @[CSR.scala 177:73:@3630.4]
  assign _T_598 = io_rw_addr == 12'hb98; // @[CSR.scala 177:73:@3631.4]
  assign _T_600 = io_rw_addr == 12'hb19; // @[CSR.scala 177:73:@3632.4]
  assign _T_602 = io_rw_addr == 12'hb99; // @[CSR.scala 177:73:@3633.4]
  assign _T_604 = io_rw_addr == 12'hb1a; // @[CSR.scala 177:73:@3634.4]
  assign _T_606 = io_rw_addr == 12'hb9a; // @[CSR.scala 177:73:@3635.4]
  assign _T_608 = io_rw_addr == 12'hb1b; // @[CSR.scala 177:73:@3636.4]
  assign _T_610 = io_rw_addr == 12'hb9b; // @[CSR.scala 177:73:@3637.4]
  assign _T_612 = io_rw_addr == 12'hb1c; // @[CSR.scala 177:73:@3638.4]
  assign _T_614 = io_rw_addr == 12'hb9c; // @[CSR.scala 177:73:@3639.4]
  assign _T_616 = io_rw_addr == 12'hb1d; // @[CSR.scala 177:73:@3640.4]
  assign _T_618 = io_rw_addr == 12'hb9d; // @[CSR.scala 177:73:@3641.4]
  assign _T_620 = io_rw_addr == 12'hb1e; // @[CSR.scala 177:73:@3642.4]
  assign _T_622 = io_rw_addr == 12'hb9e; // @[CSR.scala 177:73:@3643.4]
  assign _T_624 = io_rw_addr == 12'hb1f; // @[CSR.scala 177:73:@3644.4]
  assign _T_626 = io_rw_addr == 12'hb9f; // @[CSR.scala 177:73:@3645.4]
  assign _T_628 = io_rw_addr == 12'hb20; // @[CSR.scala 177:73:@3646.4]
  assign _T_630 = io_rw_addr == 12'hba0; // @[CSR.scala 177:73:@3647.4]
  assign _T_632 = io_rw_addr == 12'hb21; // @[CSR.scala 177:73:@3648.4]
  assign _T_634 = io_rw_addr == 12'hba1; // @[CSR.scala 177:73:@3649.4]
  assign _T_636 = io_rw_addr == 12'hb22; // @[CSR.scala 177:73:@3650.4]
  assign _T_638 = io_rw_addr == 12'hba2; // @[CSR.scala 177:73:@3651.4]
  assign _T_640 = io_rw_addr == 12'hb80; // @[CSR.scala 177:73:@3652.4]
  assign _T_642 = io_rw_addr == 12'hb82; // @[CSR.scala 177:73:@3653.4]
  assign _T_643 = io_rw_addr[9:8]; // @[CSR.scala 179:54:@3654.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_643; // @[CSR.scala 179:41:@3655.4]
  assign _T_644 = io_rw_addr[11:10]; // @[CSR.scala 180:29:@3656.4]
  assign _T_645 = ~ _T_644; // @[CSR.scala 180:37:@3657.4]
  assign read_only = _T_645 == 2'h0; // @[CSR.scala 180:37:@3658.4]
  assign _T_647 = io_rw_cmd != 3'h5; // @[CSR.scala 181:38:@3659.4]
  assign _T_648 = cpu_ren & _T_647; // @[CSR.scala 181:25:@3660.4]
  assign cpu_wen = _T_648 & priv_sufficient; // @[CSR.scala 181:48:@3661.4]
  assign _T_650 = read_only == 1'h0; // @[CSR.scala 182:24:@3662.4]
  assign wen = cpu_wen & _T_650; // @[CSR.scala 182:21:@3663.4]
  assign _T_651 = io_rw_cmd == 3'h2; // @[Util.scala 23:47:@3664.4]
  assign _T_652 = io_rw_cmd == 3'h3; // @[Util.scala 23:47:@3665.4]
  assign _T_653 = _T_651 | _T_652; // @[Util.scala 23:62:@3666.4]
  assign _T_655 = _T_653 ? io_rw_rdata : 32'h0; // @[CSR.scala 281:9:@3667.4]
  assign _T_656 = _T_655 | io_rw_wdata; // @[CSR.scala 281:49:@3668.4]
  assign _T_659 = _T_652 ? io_rw_wdata : 32'h0; // @[CSR.scala 281:64:@3670.4]
  assign _T_660 = ~ _T_659; // @[CSR.scala 281:60:@3671.4]
  assign wdata = _T_656 & _T_660; // @[CSR.scala 281:58:@3672.4]
  assign _T_662 = io_rw_addr[2:0]; // @[CSR.scala 185:33:@3673.4]
  assign opcode = 8'h1 << _T_662; // @[CSR.scala 185:20:@3674.4]
  assign _T_663 = opcode[0]; // @[CSR.scala 186:40:@3675.4]
  assign insn_call = system_insn & _T_663; // @[CSR.scala 186:31:@3676.4]
  assign _T_664 = opcode[1]; // @[CSR.scala 187:41:@3677.4]
  assign insn_break = system_insn & _T_664; // @[CSR.scala 187:32:@3678.4]
  assign _T_665 = opcode[2]; // @[CSR.scala 188:39:@3679.4]
  assign _T_666 = system_insn & _T_665; // @[CSR.scala 188:30:@3680.4]
  assign insn_ret = _T_666 & priv_sufficient; // @[CSR.scala 188:43:@3681.4]
  assign _T_940 = insn_call | insn_break; // @[CSR.scala 199:24:@3880.4]
  assign _T_942 = {{1'd0}, insn_ret}; // @[Bitwise.scala 48:55:@3883.4]
  assign _T_944 = _T_942 <= 2'h1; // @[CSR.scala 201:50:@3884.4]
  assign _T_946 = _T_944 | reset; // @[CSR.scala 201:9:@3886.4]
  assign _T_948 = _T_946 == 1'h0; // @[CSR.scala 201:9:@3887.4]
  assign _T_951 = io_rw_addr[10]; // @[CSR.scala 208:32:@3896.4]
  assign _T_953 = _T_951 == 1'h0; // @[CSR.scala 208:21:@3897.4]
  assign _T_954 = insn_ret & _T_953; // @[CSR.scala 208:18:@3898.4]
  assign _GEN_3 = _T_954 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 208:38:@3899.4]
  assign _GEN_4 = _T_954 ? 1'h1 : reg_mstatus_mpie; // @[CSR.scala 208:38:@3899.4]
  assign new_prv = _T_954 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 208:38:@3899.4]
  assign _GEN_148 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 218:35:@3907.6]
  assign _T_958 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3907.6]
  assign _T_959 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3908.6]
  assign _GEN_7 = insn_call ? 32'h80000004 : reg_mepc; // @[CSR.scala 216:18:@3905.4]
  assign _GEN_8 = insn_call ? {{28'd0}, _T_959} : reg_mcause; // @[CSR.scala 216:18:@3905.4]
  assign _GEN_9 = insn_call ? io_pc : reg_mepc; // @[CSR.scala 216:18:@3905.4]
  assign _GEN_10 = insn_break ? 32'h80000004 : _GEN_7; // @[CSR.scala 223:19:@3912.4]
  assign _GEN_11 = insn_break ? 32'h3 : _GEN_8; // @[CSR.scala 223:19:@3912.4]
  assign _GEN_12 = insn_break ? io_pc : _GEN_9; // @[CSR.scala 223:19:@3912.4]
  assign _GEN_14 = io_xcpt ? io_cause : _GEN_11; // @[CSR.scala 229:17:@3917.4]
  assign _GEN_15 = io_xcpt ? io_pc : _GEN_12; // @[CSR.scala 229:17:@3917.4]
  assign _GEN_16 = io_xcpt ? io_tval : reg_mtval; // @[CSR.scala 229:17:@3917.4]
  assign _T_965 = _T_478 ? _T_249 : 64'h0; // @[Mux.scala 19:72:@3925.4]
  assign _T_967 = _T_480 ? _T_261 : 64'h0; // @[Mux.scala 19:72:@3926.4]
  assign _T_969 = _T_482 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:@3927.4]
  assign _T_975 = _T_488 ? 31'h40000100 : 31'h0; // @[Mux.scala 19:72:@3930.4]
  assign _T_977 = _T_490 ? read_mstatus : 32'h0; // @[Mux.scala 19:72:@3931.4]
  assign _T_979 = _T_492 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:@3932.4]
  assign _T_981 = _T_494 ? _T_468 : 16'h0; // @[Mux.scala 19:72:@3933.4]
  assign _T_983 = _T_496 ? _T_474 : 16'h0; // @[Mux.scala 19:72:@3934.4]
  assign _T_985 = _T_498 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:@3935.4]
  assign _T_987 = _T_500 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:@3936.4]
  assign _T_989 = _T_502 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:@3937.4]
  assign _T_991 = _T_504 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:@3938.4]
  assign _T_995 = _T_508 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:@3940.4]
  assign _T_997 = _T_510 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:@3941.4]
  assign _T_999 = _T_512 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3942.4]
  assign _T_1001 = _T_514 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3943.4]
  assign _T_1003 = _T_516 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3944.4]
  assign _T_1005 = _T_518 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3945.4]
  assign _T_1007 = _T_520 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3946.4]
  assign _T_1009 = _T_522 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3947.4]
  assign _T_1011 = _T_524 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3948.4]
  assign _T_1013 = _T_526 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3949.4]
  assign _T_1015 = _T_528 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3950.4]
  assign _T_1017 = _T_530 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3951.4]
  assign _T_1019 = _T_532 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3952.4]
  assign _T_1021 = _T_534 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3953.4]
  assign _T_1023 = _T_536 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3954.4]
  assign _T_1025 = _T_538 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3955.4]
  assign _T_1027 = _T_540 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3956.4]
  assign _T_1029 = _T_542 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3957.4]
  assign _T_1031 = _T_544 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3958.4]
  assign _T_1033 = _T_546 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3959.4]
  assign _T_1035 = _T_548 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3960.4]
  assign _T_1037 = _T_550 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3961.4]
  assign _T_1039 = _T_552 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3962.4]
  assign _T_1041 = _T_554 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3963.4]
  assign _T_1043 = _T_556 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3964.4]
  assign _T_1045 = _T_558 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3965.4]
  assign _T_1047 = _T_560 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3966.4]
  assign _T_1049 = _T_562 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3967.4]
  assign _T_1051 = _T_564 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3968.4]
  assign _T_1053 = _T_566 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3969.4]
  assign _T_1055 = _T_568 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3970.4]
  assign _T_1057 = _T_570 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3971.4]
  assign _T_1059 = _T_572 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3972.4]
  assign _T_1061 = _T_574 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3973.4]
  assign _T_1063 = _T_576 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3974.4]
  assign _T_1065 = _T_578 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3975.4]
  assign _T_1067 = _T_580 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3976.4]
  assign _T_1069 = _T_582 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3977.4]
  assign _T_1071 = _T_584 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3978.4]
  assign _T_1073 = _T_586 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3979.4]
  assign _T_1075 = _T_588 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3980.4]
  assign _T_1077 = _T_590 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3981.4]
  assign _T_1079 = _T_592 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3982.4]
  assign _T_1081 = _T_594 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3983.4]
  assign _T_1083 = _T_596 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3984.4]
  assign _T_1085 = _T_598 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3985.4]
  assign _T_1087 = _T_600 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3986.4]
  assign _T_1089 = _T_602 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3987.4]
  assign _T_1091 = _T_604 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3988.4]
  assign _T_1093 = _T_606 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3989.4]
  assign _T_1095 = _T_608 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3990.4]
  assign _T_1097 = _T_610 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3991.4]
  assign _T_1099 = _T_612 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3992.4]
  assign _T_1101 = _T_614 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3993.4]
  assign _T_1103 = _T_616 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3994.4]
  assign _T_1105 = _T_618 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3995.4]
  assign _T_1107 = _T_620 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3996.4]
  assign _T_1109 = _T_622 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3997.4]
  assign _T_1111 = _T_624 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3998.4]
  assign _T_1113 = _T_626 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3999.4]
  assign _T_1115 = _T_628 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@4000.4]
  assign _T_1117 = _T_630 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@4001.4]
  assign _T_1119 = _T_632 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@4002.4]
  assign _T_1121 = _T_634 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@4003.4]
  assign _T_1123 = _T_636 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@4004.4]
  assign _T_1125 = _T_638 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@4005.4]
  assign _T_1130 = _T_965 | _T_967; // @[Mux.scala 19:72:@4008.4]
  assign _GEN_149 = {{48'd0}, _T_969}; // @[Mux.scala 19:72:@4009.4]
  assign _T_1131 = _T_1130 | _GEN_149; // @[Mux.scala 19:72:@4009.4]
  assign _GEN_150 = {{33'd0}, _T_975}; // @[Mux.scala 19:72:@4012.4]
  assign _T_1134 = _T_1131 | _GEN_150; // @[Mux.scala 19:72:@4012.4]
  assign _GEN_151 = {{32'd0}, _T_977}; // @[Mux.scala 19:72:@4013.4]
  assign _T_1135 = _T_1134 | _GEN_151; // @[Mux.scala 19:72:@4013.4]
  assign _GEN_152 = {{55'd0}, _T_979}; // @[Mux.scala 19:72:@4014.4]
  assign _T_1136 = _T_1135 | _GEN_152; // @[Mux.scala 19:72:@4014.4]
  assign _GEN_153 = {{48'd0}, _T_981}; // @[Mux.scala 19:72:@4015.4]
  assign _T_1137 = _T_1136 | _GEN_153; // @[Mux.scala 19:72:@4015.4]
  assign _GEN_154 = {{48'd0}, _T_983}; // @[Mux.scala 19:72:@4016.4]
  assign _T_1138 = _T_1137 | _GEN_154; // @[Mux.scala 19:72:@4016.4]
  assign _GEN_155 = {{32'd0}, _T_985}; // @[Mux.scala 19:72:@4017.4]
  assign _T_1139 = _T_1138 | _GEN_155; // @[Mux.scala 19:72:@4017.4]
  assign _GEN_156 = {{32'd0}, _T_987}; // @[Mux.scala 19:72:@4018.4]
  assign _T_1140 = _T_1139 | _GEN_156; // @[Mux.scala 19:72:@4018.4]
  assign _GEN_157 = {{32'd0}, _T_989}; // @[Mux.scala 19:72:@4019.4]
  assign _T_1141 = _T_1140 | _GEN_157; // @[Mux.scala 19:72:@4019.4]
  assign _GEN_158 = {{32'd0}, _T_991}; // @[Mux.scala 19:72:@4020.4]
  assign _T_1142 = _T_1141 | _GEN_158; // @[Mux.scala 19:72:@4020.4]
  assign _GEN_159 = {{32'd0}, _T_995}; // @[Mux.scala 19:72:@4022.4]
  assign _T_1144 = _T_1142 | _GEN_159; // @[Mux.scala 19:72:@4022.4]
  assign _GEN_160 = {{32'd0}, _T_997}; // @[Mux.scala 19:72:@4023.4]
  assign _T_1145 = _T_1144 | _GEN_160; // @[Mux.scala 19:72:@4023.4]
  assign _GEN_161 = {{24'd0}, _T_999}; // @[Mux.scala 19:72:@4024.4]
  assign _T_1146 = _T_1145 | _GEN_161; // @[Mux.scala 19:72:@4024.4]
  assign _GEN_162 = {{24'd0}, _T_1001}; // @[Mux.scala 19:72:@4025.4]
  assign _T_1147 = _T_1146 | _GEN_162; // @[Mux.scala 19:72:@4025.4]
  assign _GEN_163 = {{24'd0}, _T_1003}; // @[Mux.scala 19:72:@4026.4]
  assign _T_1148 = _T_1147 | _GEN_163; // @[Mux.scala 19:72:@4026.4]
  assign _GEN_164 = {{24'd0}, _T_1005}; // @[Mux.scala 19:72:@4027.4]
  assign _T_1149 = _T_1148 | _GEN_164; // @[Mux.scala 19:72:@4027.4]
  assign _GEN_165 = {{24'd0}, _T_1007}; // @[Mux.scala 19:72:@4028.4]
  assign _T_1150 = _T_1149 | _GEN_165; // @[Mux.scala 19:72:@4028.4]
  assign _GEN_166 = {{24'd0}, _T_1009}; // @[Mux.scala 19:72:@4029.4]
  assign _T_1151 = _T_1150 | _GEN_166; // @[Mux.scala 19:72:@4029.4]
  assign _GEN_167 = {{24'd0}, _T_1011}; // @[Mux.scala 19:72:@4030.4]
  assign _T_1152 = _T_1151 | _GEN_167; // @[Mux.scala 19:72:@4030.4]
  assign _GEN_168 = {{24'd0}, _T_1013}; // @[Mux.scala 19:72:@4031.4]
  assign _T_1153 = _T_1152 | _GEN_168; // @[Mux.scala 19:72:@4031.4]
  assign _GEN_169 = {{24'd0}, _T_1015}; // @[Mux.scala 19:72:@4032.4]
  assign _T_1154 = _T_1153 | _GEN_169; // @[Mux.scala 19:72:@4032.4]
  assign _GEN_170 = {{24'd0}, _T_1017}; // @[Mux.scala 19:72:@4033.4]
  assign _T_1155 = _T_1154 | _GEN_170; // @[Mux.scala 19:72:@4033.4]
  assign _GEN_171 = {{24'd0}, _T_1019}; // @[Mux.scala 19:72:@4034.4]
  assign _T_1156 = _T_1155 | _GEN_171; // @[Mux.scala 19:72:@4034.4]
  assign _GEN_172 = {{24'd0}, _T_1021}; // @[Mux.scala 19:72:@4035.4]
  assign _T_1157 = _T_1156 | _GEN_172; // @[Mux.scala 19:72:@4035.4]
  assign _GEN_173 = {{24'd0}, _T_1023}; // @[Mux.scala 19:72:@4036.4]
  assign _T_1158 = _T_1157 | _GEN_173; // @[Mux.scala 19:72:@4036.4]
  assign _GEN_174 = {{24'd0}, _T_1025}; // @[Mux.scala 19:72:@4037.4]
  assign _T_1159 = _T_1158 | _GEN_174; // @[Mux.scala 19:72:@4037.4]
  assign _GEN_175 = {{24'd0}, _T_1027}; // @[Mux.scala 19:72:@4038.4]
  assign _T_1160 = _T_1159 | _GEN_175; // @[Mux.scala 19:72:@4038.4]
  assign _GEN_176 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:@4039.4]
  assign _T_1161 = _T_1160 | _GEN_176; // @[Mux.scala 19:72:@4039.4]
  assign _GEN_177 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:@4040.4]
  assign _T_1162 = _T_1161 | _GEN_177; // @[Mux.scala 19:72:@4040.4]
  assign _GEN_178 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:@4041.4]
  assign _T_1163 = _T_1162 | _GEN_178; // @[Mux.scala 19:72:@4041.4]
  assign _GEN_179 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:@4042.4]
  assign _T_1164 = _T_1163 | _GEN_179; // @[Mux.scala 19:72:@4042.4]
  assign _GEN_180 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:@4043.4]
  assign _T_1165 = _T_1164 | _GEN_180; // @[Mux.scala 19:72:@4043.4]
  assign _GEN_181 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:@4044.4]
  assign _T_1166 = _T_1165 | _GEN_181; // @[Mux.scala 19:72:@4044.4]
  assign _GEN_182 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:@4045.4]
  assign _T_1167 = _T_1166 | _GEN_182; // @[Mux.scala 19:72:@4045.4]
  assign _GEN_183 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:@4046.4]
  assign _T_1168 = _T_1167 | _GEN_183; // @[Mux.scala 19:72:@4046.4]
  assign _GEN_184 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:@4047.4]
  assign _T_1169 = _T_1168 | _GEN_184; // @[Mux.scala 19:72:@4047.4]
  assign _GEN_185 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:@4048.4]
  assign _T_1170 = _T_1169 | _GEN_185; // @[Mux.scala 19:72:@4048.4]
  assign _GEN_186 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:@4049.4]
  assign _T_1171 = _T_1170 | _GEN_186; // @[Mux.scala 19:72:@4049.4]
  assign _GEN_187 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:@4050.4]
  assign _T_1172 = _T_1171 | _GEN_187; // @[Mux.scala 19:72:@4050.4]
  assign _GEN_188 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:@4051.4]
  assign _T_1173 = _T_1172 | _GEN_188; // @[Mux.scala 19:72:@4051.4]
  assign _GEN_189 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:@4052.4]
  assign _T_1174 = _T_1173 | _GEN_189; // @[Mux.scala 19:72:@4052.4]
  assign _GEN_190 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:@4053.4]
  assign _T_1175 = _T_1174 | _GEN_190; // @[Mux.scala 19:72:@4053.4]
  assign _GEN_191 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:@4054.4]
  assign _T_1176 = _T_1175 | _GEN_191; // @[Mux.scala 19:72:@4054.4]
  assign _GEN_192 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:@4055.4]
  assign _T_1177 = _T_1176 | _GEN_192; // @[Mux.scala 19:72:@4055.4]
  assign _GEN_193 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:@4056.4]
  assign _T_1178 = _T_1177 | _GEN_193; // @[Mux.scala 19:72:@4056.4]
  assign _GEN_194 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:@4057.4]
  assign _T_1179 = _T_1178 | _GEN_194; // @[Mux.scala 19:72:@4057.4]
  assign _GEN_195 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:@4058.4]
  assign _T_1180 = _T_1179 | _GEN_195; // @[Mux.scala 19:72:@4058.4]
  assign _GEN_196 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:@4059.4]
  assign _T_1181 = _T_1180 | _GEN_196; // @[Mux.scala 19:72:@4059.4]
  assign _GEN_197 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:@4060.4]
  assign _T_1182 = _T_1181 | _GEN_197; // @[Mux.scala 19:72:@4060.4]
  assign _GEN_198 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:@4061.4]
  assign _T_1183 = _T_1182 | _GEN_198; // @[Mux.scala 19:72:@4061.4]
  assign _GEN_199 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:@4062.4]
  assign _T_1184 = _T_1183 | _GEN_199; // @[Mux.scala 19:72:@4062.4]
  assign _GEN_200 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:@4063.4]
  assign _T_1185 = _T_1184 | _GEN_200; // @[Mux.scala 19:72:@4063.4]
  assign _GEN_201 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:@4064.4]
  assign _T_1186 = _T_1185 | _GEN_201; // @[Mux.scala 19:72:@4064.4]
  assign _GEN_202 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:@4065.4]
  assign _T_1187 = _T_1186 | _GEN_202; // @[Mux.scala 19:72:@4065.4]
  assign _GEN_203 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:@4066.4]
  assign _T_1188 = _T_1187 | _GEN_203; // @[Mux.scala 19:72:@4066.4]
  assign _GEN_204 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:@4067.4]
  assign _T_1189 = _T_1188 | _GEN_204; // @[Mux.scala 19:72:@4067.4]
  assign _GEN_205 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:@4068.4]
  assign _T_1190 = _T_1189 | _GEN_205; // @[Mux.scala 19:72:@4068.4]
  assign _GEN_206 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:@4069.4]
  assign _T_1191 = _T_1190 | _GEN_206; // @[Mux.scala 19:72:@4069.4]
  assign _GEN_207 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:@4070.4]
  assign _T_1192 = _T_1191 | _GEN_207; // @[Mux.scala 19:72:@4070.4]
  assign _GEN_208 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:@4071.4]
  assign _T_1193 = _T_1192 | _GEN_208; // @[Mux.scala 19:72:@4071.4]
  assign _GEN_209 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:@4072.4]
  assign _T_1194 = _T_1193 | _GEN_209; // @[Mux.scala 19:72:@4072.4]
  assign _GEN_210 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:@4073.4]
  assign _T_1195 = _T_1194 | _GEN_210; // @[Mux.scala 19:72:@4073.4]
  assign _GEN_211 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:@4074.4]
  assign _T_1196 = _T_1195 | _GEN_211; // @[Mux.scala 19:72:@4074.4]
  assign _GEN_212 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:@4075.4]
  assign _T_1197 = _T_1196 | _GEN_212; // @[Mux.scala 19:72:@4075.4]
  assign _GEN_213 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:@4076.4]
  assign _T_1198 = _T_1197 | _GEN_213; // @[Mux.scala 19:72:@4076.4]
  assign _GEN_214 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:@4077.4]
  assign _T_1199 = _T_1198 | _GEN_214; // @[Mux.scala 19:72:@4077.4]
  assign _GEN_215 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:@4078.4]
  assign _T_1200 = _T_1199 | _GEN_215; // @[Mux.scala 19:72:@4078.4]
  assign _GEN_216 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:@4079.4]
  assign _T_1201 = _T_1200 | _GEN_216; // @[Mux.scala 19:72:@4079.4]
  assign _GEN_217 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:@4080.4]
  assign _T_1202 = _T_1201 | _GEN_217; // @[Mux.scala 19:72:@4080.4]
  assign _GEN_218 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:@4081.4]
  assign _T_1203 = _T_1202 | _GEN_218; // @[Mux.scala 19:72:@4081.4]
  assign _GEN_219 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:@4082.4]
  assign _T_1204 = _T_1203 | _GEN_219; // @[Mux.scala 19:72:@4082.4]
  assign _GEN_220 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:@4083.4]
  assign _T_1205 = _T_1204 | _GEN_220; // @[Mux.scala 19:72:@4083.4]
  assign _GEN_221 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:@4084.4]
  assign _T_1206 = _T_1205 | _GEN_221; // @[Mux.scala 19:72:@4084.4]
  assign _GEN_222 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:@4085.4]
  assign _T_1207 = _T_1206 | _GEN_222; // @[Mux.scala 19:72:@4085.4]
  assign _GEN_223 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:@4086.4]
  assign _T_1208 = _T_1207 | _GEN_223; // @[Mux.scala 19:72:@4086.4]
  assign _GEN_224 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:@4087.4]
  assign _T_1209 = _T_1208 | _GEN_224; // @[Mux.scala 19:72:@4087.4]
  assign _T_1220 = wdata[3]; // @[CSR.scala 245:39:@4100.8]
  assign _T_1222 = wdata[7]; // @[CSR.scala 245:39:@4104.8]
  assign _GEN_17 = _T_490 ? _T_1220 : _GEN_3; // @[CSR.scala 244:39:@4094.6]
  assign _GEN_18 = _T_490 ? _T_1222 : _GEN_4; // @[CSR.scala 244:39:@4094.6]
  assign _T_1233 = wdata[15:0]; // @[:@4123.8 :@4124.8]
  assign _T_1235 = _T_1233[3]; // @[CSR.scala 250:35:@4127.8]
  assign _T_1237 = _T_1233[7]; // @[CSR.scala 250:35:@4131.8]
  assign _GEN_19 = _T_494 ? _T_1235 : reg_mip_msip; // @[CSR.scala 249:35:@4121.6]
  assign _GEN_20 = _T_496 ? _T_1235 : reg_mie_msip; // @[CSR.scala 253:35:@4141.6]
  assign _GEN_21 = _T_496 ? _T_1237 : reg_mie_mtip; // @[CSR.scala 253:35:@4141.6]
  assign _T_1253 = wdata[7:0]; // @[CSR.scala 277:47:@4163.8]
  assign _T_1254 = _T_264[31:0]; // @[CSR.scala 277:72:@4164.8]
  assign _T_1255 = {_T_1253,_T_1254}; // @[Cat.scala 30:58:@4165.8]
  assign _GEN_22 = _T_514 ? {{1'd0}, _T_1255} : _T_265; // @[CSR.scala 277:29:@4162.6]
  assign _T_1256 = _T_264[39:32]; // @[CSR.scala 278:45:@4169.8]
  assign _T_1257 = {_T_1256,wdata}; // @[Cat.scala 30:58:@4170.8]
  assign _GEN_23 = _T_512 ? {{1'd0}, _T_1257} : _GEN_22; // @[CSR.scala 278:29:@4168.6]
  assign _T_1259 = _T_267[31:0]; // @[CSR.scala 277:72:@4175.8]
  assign _T_1260 = {_T_1253,_T_1259}; // @[Cat.scala 30:58:@4176.8]
  assign _GEN_24 = _T_518 ? {{1'd0}, _T_1260} : _T_268; // @[CSR.scala 277:29:@4173.6]
  assign _T_1261 = _T_267[39:32]; // @[CSR.scala 278:45:@4180.8]
  assign _T_1262 = {_T_1261,wdata}; // @[Cat.scala 30:58:@4181.8]
  assign _GEN_25 = _T_516 ? {{1'd0}, _T_1262} : _GEN_24; // @[CSR.scala 278:29:@4179.6]
  assign _T_1264 = _T_270[31:0]; // @[CSR.scala 277:72:@4186.8]
  assign _T_1265 = {_T_1253,_T_1264}; // @[Cat.scala 30:58:@4187.8]
  assign _GEN_26 = _T_522 ? {{1'd0}, _T_1265} : _T_271; // @[CSR.scala 277:29:@4184.6]
  assign _T_1266 = _T_270[39:32]; // @[CSR.scala 278:45:@4191.8]
  assign _T_1267 = {_T_1266,wdata}; // @[Cat.scala 30:58:@4192.8]
  assign _GEN_27 = _T_520 ? {{1'd0}, _T_1267} : _GEN_26; // @[CSR.scala 278:29:@4190.6]
  assign _T_1269 = _T_273[31:0]; // @[CSR.scala 277:72:@4197.8]
  assign _T_1270 = {_T_1253,_T_1269}; // @[Cat.scala 30:58:@4198.8]
  assign _GEN_28 = _T_526 ? {{1'd0}, _T_1270} : _T_274; // @[CSR.scala 277:29:@4195.6]
  assign _T_1271 = _T_273[39:32]; // @[CSR.scala 278:45:@4202.8]
  assign _T_1272 = {_T_1271,wdata}; // @[Cat.scala 30:58:@4203.8]
  assign _GEN_29 = _T_524 ? {{1'd0}, _T_1272} : _GEN_28; // @[CSR.scala 278:29:@4201.6]
  assign _T_1274 = _T_276[31:0]; // @[CSR.scala 277:72:@4208.8]
  assign _T_1275 = {_T_1253,_T_1274}; // @[Cat.scala 30:58:@4209.8]
  assign _GEN_30 = _T_530 ? {{1'd0}, _T_1275} : _T_277; // @[CSR.scala 277:29:@4206.6]
  assign _T_1276 = _T_276[39:32]; // @[CSR.scala 278:45:@4213.8]
  assign _T_1277 = {_T_1276,wdata}; // @[Cat.scala 30:58:@4214.8]
  assign _GEN_31 = _T_528 ? {{1'd0}, _T_1277} : _GEN_30; // @[CSR.scala 278:29:@4212.6]
  assign _T_1279 = _T_279[31:0]; // @[CSR.scala 277:72:@4219.8]
  assign _T_1280 = {_T_1253,_T_1279}; // @[Cat.scala 30:58:@4220.8]
  assign _GEN_32 = _T_534 ? {{1'd0}, _T_1280} : _T_280; // @[CSR.scala 277:29:@4217.6]
  assign _T_1281 = _T_279[39:32]; // @[CSR.scala 278:45:@4224.8]
  assign _T_1282 = {_T_1281,wdata}; // @[Cat.scala 30:58:@4225.8]
  assign _GEN_33 = _T_532 ? {{1'd0}, _T_1282} : _GEN_32; // @[CSR.scala 278:29:@4223.6]
  assign _T_1284 = _T_282[31:0]; // @[CSR.scala 277:72:@4230.8]
  assign _T_1285 = {_T_1253,_T_1284}; // @[Cat.scala 30:58:@4231.8]
  assign _GEN_34 = _T_538 ? {{1'd0}, _T_1285} : _T_283; // @[CSR.scala 277:29:@4228.6]
  assign _T_1286 = _T_282[39:32]; // @[CSR.scala 278:45:@4235.8]
  assign _T_1287 = {_T_1286,wdata}; // @[Cat.scala 30:58:@4236.8]
  assign _GEN_35 = _T_536 ? {{1'd0}, _T_1287} : _GEN_34; // @[CSR.scala 278:29:@4234.6]
  assign _T_1289 = _T_285[31:0]; // @[CSR.scala 277:72:@4241.8]
  assign _T_1290 = {_T_1253,_T_1289}; // @[Cat.scala 30:58:@4242.8]
  assign _GEN_36 = _T_542 ? {{1'd0}, _T_1290} : _T_286; // @[CSR.scala 277:29:@4239.6]
  assign _T_1291 = _T_285[39:32]; // @[CSR.scala 278:45:@4246.8]
  assign _T_1292 = {_T_1291,wdata}; // @[Cat.scala 30:58:@4247.8]
  assign _GEN_37 = _T_540 ? {{1'd0}, _T_1292} : _GEN_36; // @[CSR.scala 278:29:@4245.6]
  assign _T_1294 = _T_288[31:0]; // @[CSR.scala 277:72:@4252.8]
  assign _T_1295 = {_T_1253,_T_1294}; // @[Cat.scala 30:58:@4253.8]
  assign _GEN_38 = _T_546 ? {{1'd0}, _T_1295} : _T_289; // @[CSR.scala 277:29:@4250.6]
  assign _T_1296 = _T_288[39:32]; // @[CSR.scala 278:45:@4257.8]
  assign _T_1297 = {_T_1296,wdata}; // @[Cat.scala 30:58:@4258.8]
  assign _GEN_39 = _T_544 ? {{1'd0}, _T_1297} : _GEN_38; // @[CSR.scala 278:29:@4256.6]
  assign _T_1299 = _T_291[31:0]; // @[CSR.scala 277:72:@4263.8]
  assign _T_1300 = {_T_1253,_T_1299}; // @[Cat.scala 30:58:@4264.8]
  assign _GEN_40 = _T_550 ? {{1'd0}, _T_1300} : _T_292; // @[CSR.scala 277:29:@4261.6]
  assign _T_1301 = _T_291[39:32]; // @[CSR.scala 278:45:@4268.8]
  assign _T_1302 = {_T_1301,wdata}; // @[Cat.scala 30:58:@4269.8]
  assign _GEN_41 = _T_548 ? {{1'd0}, _T_1302} : _GEN_40; // @[CSR.scala 278:29:@4267.6]
  assign _T_1304 = _T_294[31:0]; // @[CSR.scala 277:72:@4274.8]
  assign _T_1305 = {_T_1253,_T_1304}; // @[Cat.scala 30:58:@4275.8]
  assign _GEN_42 = _T_554 ? {{1'd0}, _T_1305} : _T_295; // @[CSR.scala 277:29:@4272.6]
  assign _T_1306 = _T_294[39:32]; // @[CSR.scala 278:45:@4279.8]
  assign _T_1307 = {_T_1306,wdata}; // @[Cat.scala 30:58:@4280.8]
  assign _GEN_43 = _T_552 ? {{1'd0}, _T_1307} : _GEN_42; // @[CSR.scala 278:29:@4278.6]
  assign _T_1309 = _T_297[31:0]; // @[CSR.scala 277:72:@4285.8]
  assign _T_1310 = {_T_1253,_T_1309}; // @[Cat.scala 30:58:@4286.8]
  assign _GEN_44 = _T_558 ? {{1'd0}, _T_1310} : _T_298; // @[CSR.scala 277:29:@4283.6]
  assign _T_1311 = _T_297[39:32]; // @[CSR.scala 278:45:@4290.8]
  assign _T_1312 = {_T_1311,wdata}; // @[Cat.scala 30:58:@4291.8]
  assign _GEN_45 = _T_556 ? {{1'd0}, _T_1312} : _GEN_44; // @[CSR.scala 278:29:@4289.6]
  assign _T_1314 = _T_300[31:0]; // @[CSR.scala 277:72:@4296.8]
  assign _T_1315 = {_T_1253,_T_1314}; // @[Cat.scala 30:58:@4297.8]
  assign _GEN_46 = _T_562 ? {{1'd0}, _T_1315} : _T_301; // @[CSR.scala 277:29:@4294.6]
  assign _T_1316 = _T_300[39:32]; // @[CSR.scala 278:45:@4301.8]
  assign _T_1317 = {_T_1316,wdata}; // @[Cat.scala 30:58:@4302.8]
  assign _GEN_47 = _T_560 ? {{1'd0}, _T_1317} : _GEN_46; // @[CSR.scala 278:29:@4300.6]
  assign _T_1319 = _T_303[31:0]; // @[CSR.scala 277:72:@4307.8]
  assign _T_1320 = {_T_1253,_T_1319}; // @[Cat.scala 30:58:@4308.8]
  assign _GEN_48 = _T_566 ? {{1'd0}, _T_1320} : _T_304; // @[CSR.scala 277:29:@4305.6]
  assign _T_1321 = _T_303[39:32]; // @[CSR.scala 278:45:@4312.8]
  assign _T_1322 = {_T_1321,wdata}; // @[Cat.scala 30:58:@4313.8]
  assign _GEN_49 = _T_564 ? {{1'd0}, _T_1322} : _GEN_48; // @[CSR.scala 278:29:@4311.6]
  assign _T_1324 = _T_306[31:0]; // @[CSR.scala 277:72:@4318.8]
  assign _T_1325 = {_T_1253,_T_1324}; // @[Cat.scala 30:58:@4319.8]
  assign _GEN_50 = _T_570 ? {{1'd0}, _T_1325} : _T_307; // @[CSR.scala 277:29:@4316.6]
  assign _T_1326 = _T_306[39:32]; // @[CSR.scala 278:45:@4323.8]
  assign _T_1327 = {_T_1326,wdata}; // @[Cat.scala 30:58:@4324.8]
  assign _GEN_51 = _T_568 ? {{1'd0}, _T_1327} : _GEN_50; // @[CSR.scala 278:29:@4322.6]
  assign _T_1329 = _T_309[31:0]; // @[CSR.scala 277:72:@4329.8]
  assign _T_1330 = {_T_1253,_T_1329}; // @[Cat.scala 30:58:@4330.8]
  assign _GEN_52 = _T_574 ? {{1'd0}, _T_1330} : _T_310; // @[CSR.scala 277:29:@4327.6]
  assign _T_1331 = _T_309[39:32]; // @[CSR.scala 278:45:@4334.8]
  assign _T_1332 = {_T_1331,wdata}; // @[Cat.scala 30:58:@4335.8]
  assign _GEN_53 = _T_572 ? {{1'd0}, _T_1332} : _GEN_52; // @[CSR.scala 278:29:@4333.6]
  assign _T_1334 = _T_312[31:0]; // @[CSR.scala 277:72:@4340.8]
  assign _T_1335 = {_T_1253,_T_1334}; // @[Cat.scala 30:58:@4341.8]
  assign _GEN_54 = _T_578 ? {{1'd0}, _T_1335} : _T_313; // @[CSR.scala 277:29:@4338.6]
  assign _T_1336 = _T_312[39:32]; // @[CSR.scala 278:45:@4345.8]
  assign _T_1337 = {_T_1336,wdata}; // @[Cat.scala 30:58:@4346.8]
  assign _GEN_55 = _T_576 ? {{1'd0}, _T_1337} : _GEN_54; // @[CSR.scala 278:29:@4344.6]
  assign _T_1339 = _T_315[31:0]; // @[CSR.scala 277:72:@4351.8]
  assign _T_1340 = {_T_1253,_T_1339}; // @[Cat.scala 30:58:@4352.8]
  assign _GEN_56 = _T_582 ? {{1'd0}, _T_1340} : _T_316; // @[CSR.scala 277:29:@4349.6]
  assign _T_1341 = _T_315[39:32]; // @[CSR.scala 278:45:@4356.8]
  assign _T_1342 = {_T_1341,wdata}; // @[Cat.scala 30:58:@4357.8]
  assign _GEN_57 = _T_580 ? {{1'd0}, _T_1342} : _GEN_56; // @[CSR.scala 278:29:@4355.6]
  assign _T_1344 = _T_318[31:0]; // @[CSR.scala 277:72:@4362.8]
  assign _T_1345 = {_T_1253,_T_1344}; // @[Cat.scala 30:58:@4363.8]
  assign _GEN_58 = _T_586 ? {{1'd0}, _T_1345} : _T_319; // @[CSR.scala 277:29:@4360.6]
  assign _T_1346 = _T_318[39:32]; // @[CSR.scala 278:45:@4367.8]
  assign _T_1347 = {_T_1346,wdata}; // @[Cat.scala 30:58:@4368.8]
  assign _GEN_59 = _T_584 ? {{1'd0}, _T_1347} : _GEN_58; // @[CSR.scala 278:29:@4366.6]
  assign _T_1349 = _T_321[31:0]; // @[CSR.scala 277:72:@4373.8]
  assign _T_1350 = {_T_1253,_T_1349}; // @[Cat.scala 30:58:@4374.8]
  assign _GEN_60 = _T_590 ? {{1'd0}, _T_1350} : _T_322; // @[CSR.scala 277:29:@4371.6]
  assign _T_1351 = _T_321[39:32]; // @[CSR.scala 278:45:@4378.8]
  assign _T_1352 = {_T_1351,wdata}; // @[Cat.scala 30:58:@4379.8]
  assign _GEN_61 = _T_588 ? {{1'd0}, _T_1352} : _GEN_60; // @[CSR.scala 278:29:@4377.6]
  assign _T_1354 = _T_324[31:0]; // @[CSR.scala 277:72:@4384.8]
  assign _T_1355 = {_T_1253,_T_1354}; // @[Cat.scala 30:58:@4385.8]
  assign _GEN_62 = _T_594 ? {{1'd0}, _T_1355} : _T_325; // @[CSR.scala 277:29:@4382.6]
  assign _T_1356 = _T_324[39:32]; // @[CSR.scala 278:45:@4389.8]
  assign _T_1357 = {_T_1356,wdata}; // @[Cat.scala 30:58:@4390.8]
  assign _GEN_63 = _T_592 ? {{1'd0}, _T_1357} : _GEN_62; // @[CSR.scala 278:29:@4388.6]
  assign _T_1359 = _T_327[31:0]; // @[CSR.scala 277:72:@4395.8]
  assign _T_1360 = {_T_1253,_T_1359}; // @[Cat.scala 30:58:@4396.8]
  assign _GEN_64 = _T_598 ? {{1'd0}, _T_1360} : _T_328; // @[CSR.scala 277:29:@4393.6]
  assign _T_1361 = _T_327[39:32]; // @[CSR.scala 278:45:@4400.8]
  assign _T_1362 = {_T_1361,wdata}; // @[Cat.scala 30:58:@4401.8]
  assign _GEN_65 = _T_596 ? {{1'd0}, _T_1362} : _GEN_64; // @[CSR.scala 278:29:@4399.6]
  assign _T_1364 = _T_330[31:0]; // @[CSR.scala 277:72:@4406.8]
  assign _T_1365 = {_T_1253,_T_1364}; // @[Cat.scala 30:58:@4407.8]
  assign _GEN_66 = _T_602 ? {{1'd0}, _T_1365} : _T_331; // @[CSR.scala 277:29:@4404.6]
  assign _T_1366 = _T_330[39:32]; // @[CSR.scala 278:45:@4411.8]
  assign _T_1367 = {_T_1366,wdata}; // @[Cat.scala 30:58:@4412.8]
  assign _GEN_67 = _T_600 ? {{1'd0}, _T_1367} : _GEN_66; // @[CSR.scala 278:29:@4410.6]
  assign _T_1369 = _T_333[31:0]; // @[CSR.scala 277:72:@4417.8]
  assign _T_1370 = {_T_1253,_T_1369}; // @[Cat.scala 30:58:@4418.8]
  assign _GEN_68 = _T_606 ? {{1'd0}, _T_1370} : _T_334; // @[CSR.scala 277:29:@4415.6]
  assign _T_1371 = _T_333[39:32]; // @[CSR.scala 278:45:@4422.8]
  assign _T_1372 = {_T_1371,wdata}; // @[Cat.scala 30:58:@4423.8]
  assign _GEN_69 = _T_604 ? {{1'd0}, _T_1372} : _GEN_68; // @[CSR.scala 278:29:@4421.6]
  assign _T_1374 = _T_336[31:0]; // @[CSR.scala 277:72:@4428.8]
  assign _T_1375 = {_T_1253,_T_1374}; // @[Cat.scala 30:58:@4429.8]
  assign _GEN_70 = _T_610 ? {{1'd0}, _T_1375} : _T_337; // @[CSR.scala 277:29:@4426.6]
  assign _T_1376 = _T_336[39:32]; // @[CSR.scala 278:45:@4433.8]
  assign _T_1377 = {_T_1376,wdata}; // @[Cat.scala 30:58:@4434.8]
  assign _GEN_71 = _T_608 ? {{1'd0}, _T_1377} : _GEN_70; // @[CSR.scala 278:29:@4432.6]
  assign _T_1379 = _T_339[31:0]; // @[CSR.scala 277:72:@4439.8]
  assign _T_1380 = {_T_1253,_T_1379}; // @[Cat.scala 30:58:@4440.8]
  assign _GEN_72 = _T_614 ? {{1'd0}, _T_1380} : _T_340; // @[CSR.scala 277:29:@4437.6]
  assign _T_1381 = _T_339[39:32]; // @[CSR.scala 278:45:@4444.8]
  assign _T_1382 = {_T_1381,wdata}; // @[Cat.scala 30:58:@4445.8]
  assign _GEN_73 = _T_612 ? {{1'd0}, _T_1382} : _GEN_72; // @[CSR.scala 278:29:@4443.6]
  assign _T_1384 = _T_342[31:0]; // @[CSR.scala 277:72:@4450.8]
  assign _T_1385 = {_T_1253,_T_1384}; // @[Cat.scala 30:58:@4451.8]
  assign _GEN_74 = _T_618 ? {{1'd0}, _T_1385} : _T_343; // @[CSR.scala 277:29:@4448.6]
  assign _T_1386 = _T_342[39:32]; // @[CSR.scala 278:45:@4455.8]
  assign _T_1387 = {_T_1386,wdata}; // @[Cat.scala 30:58:@4456.8]
  assign _GEN_75 = _T_616 ? {{1'd0}, _T_1387} : _GEN_74; // @[CSR.scala 278:29:@4454.6]
  assign _T_1389 = _T_345[31:0]; // @[CSR.scala 277:72:@4461.8]
  assign _T_1390 = {_T_1253,_T_1389}; // @[Cat.scala 30:58:@4462.8]
  assign _GEN_76 = _T_622 ? {{1'd0}, _T_1390} : _T_346; // @[CSR.scala 277:29:@4459.6]
  assign _T_1391 = _T_345[39:32]; // @[CSR.scala 278:45:@4466.8]
  assign _T_1392 = {_T_1391,wdata}; // @[Cat.scala 30:58:@4467.8]
  assign _GEN_77 = _T_620 ? {{1'd0}, _T_1392} : _GEN_76; // @[CSR.scala 278:29:@4465.6]
  assign _T_1394 = _T_348[31:0]; // @[CSR.scala 277:72:@4472.8]
  assign _T_1395 = {_T_1253,_T_1394}; // @[Cat.scala 30:58:@4473.8]
  assign _GEN_78 = _T_626 ? {{1'd0}, _T_1395} : _T_349; // @[CSR.scala 277:29:@4470.6]
  assign _T_1396 = _T_348[39:32]; // @[CSR.scala 278:45:@4477.8]
  assign _T_1397 = {_T_1396,wdata}; // @[Cat.scala 30:58:@4478.8]
  assign _GEN_79 = _T_624 ? {{1'd0}, _T_1397} : _GEN_78; // @[CSR.scala 278:29:@4476.6]
  assign _T_1399 = _T_351[31:0]; // @[CSR.scala 277:72:@4483.8]
  assign _T_1400 = {_T_1253,_T_1399}; // @[Cat.scala 30:58:@4484.8]
  assign _GEN_80 = _T_630 ? {{1'd0}, _T_1400} : _T_352; // @[CSR.scala 277:29:@4481.6]
  assign _T_1401 = _T_351[39:32]; // @[CSR.scala 278:45:@4488.8]
  assign _T_1402 = {_T_1401,wdata}; // @[Cat.scala 30:58:@4489.8]
  assign _GEN_81 = _T_628 ? {{1'd0}, _T_1402} : _GEN_80; // @[CSR.scala 278:29:@4487.6]
  assign _T_1404 = _T_354[31:0]; // @[CSR.scala 277:72:@4494.8]
  assign _T_1405 = {_T_1253,_T_1404}; // @[Cat.scala 30:58:@4495.8]
  assign _GEN_82 = _T_634 ? {{1'd0}, _T_1405} : _T_355; // @[CSR.scala 277:29:@4492.6]
  assign _T_1406 = _T_354[39:32]; // @[CSR.scala 278:45:@4499.8]
  assign _T_1407 = {_T_1406,wdata}; // @[Cat.scala 30:58:@4500.8]
  assign _GEN_83 = _T_632 ? {{1'd0}, _T_1407} : _GEN_82; // @[CSR.scala 278:29:@4498.6]
  assign _T_1409 = _T_357[31:0]; // @[CSR.scala 277:72:@4505.8]
  assign _T_1410 = {_T_1253,_T_1409}; // @[Cat.scala 30:58:@4506.8]
  assign _GEN_84 = _T_638 ? {{1'd0}, _T_1410} : _T_358; // @[CSR.scala 277:29:@4503.6]
  assign _T_1411 = _T_357[39:32]; // @[CSR.scala 278:45:@4510.8]
  assign _T_1412 = {_T_1411,wdata}; // @[Cat.scala 30:58:@4511.8]
  assign _GEN_85 = _T_636 ? {{1'd0}, _T_1412} : _GEN_84; // @[CSR.scala 278:29:@4509.6]
  assign _T_1414 = _T_249[31:0]; // @[CSR.scala 277:72:@4516.8]
  assign _T_1415 = {wdata,_T_1414}; // @[Cat.scala 30:58:@4517.8]
  assign _T_1416 = _T_1415[63:6]; // @[Util.scala 133:28:@4519.8]
  assign _GEN_86 = _T_640 ? _T_1415 : {{57'd0}, _T_241}; // @[CSR.scala 277:29:@4514.6]
  assign _GEN_87 = _T_640 ? _T_1416 : _GEN_0; // @[CSR.scala 277:29:@4514.6]
  assign _T_1417 = _T_249[63:32]; // @[CSR.scala 278:45:@4523.8]
  assign _T_1418 = {_T_1417,wdata}; // @[Cat.scala 30:58:@4524.8]
  assign _T_1419 = _T_1418[63:6]; // @[Util.scala 133:28:@4526.8]
  assign _GEN_88 = _T_478 ? _T_1418 : _GEN_86; // @[CSR.scala 278:29:@4522.6]
  assign _GEN_89 = _T_478 ? _T_1419 : _GEN_87; // @[CSR.scala 278:29:@4522.6]
  assign _T_1421 = _T_261[31:0]; // @[CSR.scala 277:72:@4531.8]
  assign _T_1422 = {wdata,_T_1421}; // @[Cat.scala 30:58:@4532.8]
  assign _T_1423 = _T_1422[63:6]; // @[Util.scala 133:28:@4534.8]
  assign _GEN_90 = _T_642 ? _T_1422 : {{57'd0}, _T_253}; // @[CSR.scala 277:29:@4529.6]
  assign _GEN_91 = _T_642 ? _T_1423 : _GEN_1; // @[CSR.scala 277:29:@4529.6]
  assign _T_1424 = _T_261[63:32]; // @[CSR.scala 278:45:@4538.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:@4539.8]
  assign _T_1426 = _T_1425[63:6]; // @[Util.scala 133:28:@4541.8]
  assign _GEN_92 = _T_480 ? _T_1425 : _GEN_90; // @[CSR.scala 278:29:@4537.6]
  assign _GEN_93 = _T_480 ? _T_1426 : _GEN_91; // @[CSR.scala 278:29:@4537.6]
  assign _GEN_94 = _T_508 ? wdata : reg_dscratch; // @[CSR.scala 265:40:@4544.6]
  assign _T_1429 = wdata >> 2'h2; // @[CSR.scala 267:78:@4549.8]
  assign _GEN_225 = {{3'd0}, _T_1429}; // @[CSR.scala 267:86:@4550.8]
  assign _T_1431 = _GEN_225 << 2'h2; // @[CSR.scala 267:86:@4550.8]
  assign _GEN_95 = _T_500 ? _T_1431 : {{3'd0}, _GEN_15}; // @[CSR.scala 267:40:@4547.6]
  assign _GEN_96 = _T_498 ? wdata : reg_mscratch; // @[CSR.scala 268:40:@4553.6]
  assign _T_1433 = wdata & 32'h8000001f; // @[CSR.scala 269:62:@4557.8]
  assign _GEN_97 = _T_504 ? _T_1433 : _GEN_14; // @[CSR.scala 269:40:@4556.6]
  assign _GEN_98 = _T_502 ? wdata : _GEN_16; // @[CSR.scala 270:40:@4560.6]
  assign _GEN_99 = _T_510 ? wdata : reg_medeleg; // @[CSR.scala 271:42:@4564.6]
  assign _GEN_100 = wen ? _GEN_17 : _GEN_3; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_101 = wen ? _GEN_18 : _GEN_4; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_102 = wen ? _GEN_19 : reg_mip_msip; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_103 = wen ? _GEN_20 : reg_mie_msip; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_104 = wen ? _GEN_21 : reg_mie_mtip; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_105 = wen ? _GEN_23 : _T_265; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_106 = wen ? _GEN_25 : _T_268; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_107 = wen ? _GEN_27 : _T_271; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_108 = wen ? _GEN_29 : _T_274; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_109 = wen ? _GEN_31 : _T_277; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_110 = wen ? _GEN_33 : _T_280; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_111 = wen ? _GEN_35 : _T_283; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_112 = wen ? _GEN_37 : _T_286; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_113 = wen ? _GEN_39 : _T_289; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_114 = wen ? _GEN_41 : _T_292; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_115 = wen ? _GEN_43 : _T_295; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_116 = wen ? _GEN_45 : _T_298; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_117 = wen ? _GEN_47 : _T_301; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_118 = wen ? _GEN_49 : _T_304; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_119 = wen ? _GEN_51 : _T_307; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_120 = wen ? _GEN_53 : _T_310; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_121 = wen ? _GEN_55 : _T_313; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_122 = wen ? _GEN_57 : _T_316; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_123 = wen ? _GEN_59 : _T_319; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_124 = wen ? _GEN_61 : _T_322; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_125 = wen ? _GEN_63 : _T_325; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_126 = wen ? _GEN_65 : _T_328; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_127 = wen ? _GEN_67 : _T_331; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_128 = wen ? _GEN_69 : _T_334; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_129 = wen ? _GEN_71 : _T_337; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_130 = wen ? _GEN_73 : _T_340; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_131 = wen ? _GEN_75 : _T_343; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_132 = wen ? _GEN_77 : _T_346; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_133 = wen ? _GEN_79 : _T_349; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_134 = wen ? _GEN_81 : _T_352; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_135 = wen ? _GEN_83 : _T_355; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_136 = wen ? _GEN_85 : _T_358; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_137 = wen ? _GEN_88 : {{57'd0}, _T_241}; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_138 = wen ? _GEN_89 : _GEN_0; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_139 = wen ? _GEN_92 : {{57'd0}, _T_253}; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_140 = wen ? _GEN_93 : _GEN_1; // @[CSR.scala 242:14:@4093.4]
  assign _GEN_142 = wen ? _GEN_95 : {{3'd0}, _GEN_15}; // @[CSR.scala 242:14:@4093.4]
  assign io_rw_rdata = _T_1209[31:0]; // @[CSR.scala 240:15:@4092.4]
  assign io_eret = _T_940 | insn_ret; // @[CSR.scala 199:11:@3882.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 197:13:@3879.4]
  assign io_status_unimp5 = 14'h0; // @[CSR.scala 197:13:@3878.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 197:13:@3877.4]
  assign io_status_unimp4 = 2'h0; // @[CSR.scala 197:13:@3876.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 197:13:@3875.4]
  assign io_status_unimp3 = 3'h0; // @[CSR.scala 197:13:@3874.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 197:13:@3873.4]
  assign io_status_unimp2 = 3'h0; // @[CSR.scala 197:13:@3872.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 197:13:@3871.4]
  assign io_status_unimp1 = 3'h0; // @[CSR.scala 197:13:@3870.4]
  assign io_evec = io_xcpt ? 32'h80000004 : _GEN_10; // @[CSR.scala 212:13:@3903.6 CSR.scala 217:13:@3906.6 CSR.scala 224:13:@3913.6 CSR.scala 230:13:@3918.6]
  assign io_time = _T_249[31:0]; // @[CSR.scala 236:11:@3923.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_240 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_244 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_252 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_256 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_264 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_267 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_270 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_273 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_276 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_279 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_282 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_285 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_288 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_291 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_294 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_297 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_300 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_303 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_306 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_309 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_312 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_315 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_318 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_321 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_324 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_327 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_330 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_333 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_336 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_339 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_342 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_345 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_348 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_351 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_354 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_357 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_954) begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mpie <= _T_1222;
        end else begin
          if (_T_954) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mpie <= 1'h1;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mie <= _T_1220;
        end else begin
          if (_T_954) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end
    end
    reg_mepc <= _GEN_142[31:0];
    if (wen) begin
      if (_T_504) begin
        reg_mcause <= _T_1433;
      end else begin
        if (io_xcpt) begin
          reg_mcause <= io_cause;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_959};
            end
          end
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mcause <= io_cause;
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_959};
          end
        end
      end
    end
    if (wen) begin
      if (_T_502) begin
        reg_mtval <= wdata;
      end else begin
        if (io_xcpt) begin
          reg_mtval <= io_tval;
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mtval <= io_tval;
      end
    end
    if (wen) begin
      if (_T_498) begin
        reg_mscratch <= wdata;
      end
    end
    if (wen) begin
      if (_T_510) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (reset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_494) begin
          reg_mip_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_mtip <= _T_1237;
        end
      end
    end
    if (reset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      _T_240 <= 6'h0;
    end else begin
      _T_240 <= _GEN_137[5:0];
    end
    if (reset) begin
      _T_244 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_478) begin
          _T_244 <= _T_1419;
        end else begin
          if (_T_640) begin
            _T_244 <= _T_1416;
          end else begin
            if (_T_245) begin
              _T_244 <= _T_248;
            end
          end
        end
      end else begin
        if (_T_245) begin
          _T_244 <= _T_248;
        end
      end
    end
    if (reset) begin
      _T_252 <= 6'h0;
    end else begin
      _T_252 <= _GEN_139[5:0];
    end
    if (reset) begin
      _T_256 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_480) begin
          _T_256 <= _T_1426;
        end else begin
          if (_T_642) begin
            _T_256 <= _T_1423;
          end else begin
            if (_T_257) begin
              _T_256 <= _T_260;
            end
          end
        end
      end else begin
        if (_T_257) begin
          _T_256 <= _T_260;
        end
      end
    end
    _T_264 <= _GEN_105[39:0];
    _T_267 <= _GEN_106[39:0];
    _T_270 <= _GEN_107[39:0];
    _T_273 <= _GEN_108[39:0];
    _T_276 <= _GEN_109[39:0];
    _T_279 <= _GEN_110[39:0];
    _T_282 <= _GEN_111[39:0];
    _T_285 <= _GEN_112[39:0];
    _T_288 <= _GEN_113[39:0];
    _T_291 <= _GEN_114[39:0];
    _T_294 <= _GEN_115[39:0];
    _T_297 <= _GEN_116[39:0];
    _T_300 <= _GEN_117[39:0];
    _T_303 <= _GEN_118[39:0];
    _T_306 <= _GEN_119[39:0];
    _T_309 <= _GEN_120[39:0];
    _T_312 <= _GEN_121[39:0];
    _T_315 <= _GEN_122[39:0];
    _T_318 <= _GEN_123[39:0];
    _T_321 <= _GEN_124[39:0];
    _T_324 <= _GEN_125[39:0];
    _T_327 <= _GEN_126[39:0];
    _T_330 <= _GEN_127[39:0];
    _T_333 <= _GEN_128[39:0];
    _T_336 <= _GEN_129[39:0];
    _T_339 <= _GEN_130[39:0];
    _T_342 <= _GEN_131[39:0];
    _T_345 <= _GEN_132[39:0];
    _T_348 <= _GEN_133[39:0];
    _T_351 <= _GEN_134[39:0];
    _T_354 <= _GEN_135[39:0];
    _T_357 <= _GEN_136[39:0];
    if (wen) begin
      if (_T_508) begin
        reg_dscratch <= wdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:201 assert(PopCount(insn_ret :: io.illegal :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 201:9:@3889.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[CSR.scala 201:9:@3890.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module InstDecoder( // @[:@4570.2]
  input  [31:0] io_inst, // @[:@4573.4]
  output [3:0]  io_cinfo_br_type, // @[:@4573.4]
  output [1:0]  io_cinfo_op1_sel, // @[:@4573.4]
  output [2:0]  io_cinfo_op2_sel, // @[:@4573.4]
  output        io_cinfo_rs1_oen, // @[:@4573.4]
  output        io_cinfo_rs2_oen, // @[:@4573.4]
  output [3:0]  io_cinfo_alu_fun, // @[:@4573.4]
  output [1:0]  io_cinfo_wb_sel, // @[:@4573.4]
  output        io_cinfo_rf_wen, // @[:@4573.4]
  output        io_cinfo_mem_en, // @[:@4573.4]
  output        io_cinfo_mem_fcn, // @[:@4573.4]
  output [2:0]  io_cinfo_mem_typ, // @[:@4573.4]
  output [2:0]  io_cinfo_csr_cmd, // @[:@4573.4]
  output        io_cinfo_illegal, // @[:@4573.4]
  output        io_cinfo_is_branch, // @[:@4573.4]
  output        io_cinfo_jal, // @[:@4573.4]
  output        io_cinfo_ret, // @[:@4573.4]
  output [4:0]  io_cinfo_rs1_addr, // @[:@4573.4]
  output [4:0]  io_cinfo_rs2_addr, // @[:@4573.4]
  output [4:0]  io_cinfo_wbaddr, // @[:@4573.4]
  output [31:0] io_dinfo_imm_i, // @[:@4573.4]
  output [31:0] io_dinfo_imm_s, // @[:@4573.4]
  output [31:0] io_dinfo_imm_sb, // @[:@4573.4]
  output [31:0] io_dinfo_imm_u, // @[:@4573.4]
  output [31:0] io_dinfo_imm_uj, // @[:@4573.4]
  output [31:0] io_dinfo_imm_z // @[:@4573.4]
);
  wire [31:0] _T_13; // @[Lookup.scala 9:38:@4575.4]
  wire  _T_14; // @[Lookup.scala 9:38:@4576.4]
  wire  _T_18; // @[Lookup.scala 9:38:@4578.4]
  wire  _T_22; // @[Lookup.scala 9:38:@4580.4]
  wire  _T_26; // @[Lookup.scala 9:38:@4582.4]
  wire  _T_30; // @[Lookup.scala 9:38:@4584.4]
  wire  _T_34; // @[Lookup.scala 9:38:@4586.4]
  wire  _T_38; // @[Lookup.scala 9:38:@4588.4]
  wire  _T_42; // @[Lookup.scala 9:38:@4590.4]
  wire [31:0] _T_45; // @[Lookup.scala 9:38:@4591.4]
  wire  _T_46; // @[Lookup.scala 9:38:@4592.4]
  wire  _T_50; // @[Lookup.scala 9:38:@4594.4]
  wire  _T_54; // @[Lookup.scala 9:38:@4596.4]
  wire  _T_58; // @[Lookup.scala 9:38:@4598.4]
  wire  _T_62; // @[Lookup.scala 9:38:@4600.4]
  wire  _T_66; // @[Lookup.scala 9:38:@4602.4]
  wire  _T_70; // @[Lookup.scala 9:38:@4604.4]
  wire  _T_74; // @[Lookup.scala 9:38:@4606.4]
  wire [31:0] _T_77; // @[Lookup.scala 9:38:@4607.4]
  wire  _T_78; // @[Lookup.scala 9:38:@4608.4]
  wire  _T_82; // @[Lookup.scala 9:38:@4610.4]
  wire  _T_86; // @[Lookup.scala 9:38:@4612.4]
  wire [31:0] _T_89; // @[Lookup.scala 9:38:@4613.4]
  wire  _T_90; // @[Lookup.scala 9:38:@4614.4]
  wire  _T_94; // @[Lookup.scala 9:38:@4616.4]
  wire  _T_98; // @[Lookup.scala 9:38:@4618.4]
  wire  _T_102; // @[Lookup.scala 9:38:@4620.4]
  wire  _T_106; // @[Lookup.scala 9:38:@4622.4]
  wire  _T_110; // @[Lookup.scala 9:38:@4624.4]
  wire  _T_114; // @[Lookup.scala 9:38:@4626.4]
  wire  _T_118; // @[Lookup.scala 9:38:@4628.4]
  wire  _T_122; // @[Lookup.scala 9:38:@4630.4]
  wire  _T_126; // @[Lookup.scala 9:38:@4632.4]
  wire  _T_130; // @[Lookup.scala 9:38:@4634.4]
  wire  _T_134; // @[Lookup.scala 9:38:@4636.4]
  wire  _T_138; // @[Lookup.scala 9:38:@4638.4]
  wire  _T_142; // @[Lookup.scala 9:38:@4640.4]
  wire  _T_146; // @[Lookup.scala 9:38:@4642.4]
  wire  _T_150; // @[Lookup.scala 9:38:@4644.4]
  wire  _T_154; // @[Lookup.scala 9:38:@4646.4]
  wire  _T_158; // @[Lookup.scala 9:38:@4648.4]
  wire  _T_162; // @[Lookup.scala 9:38:@4650.4]
  wire  _T_166; // @[Lookup.scala 9:38:@4652.4]
  wire  _T_170; // @[Lookup.scala 9:38:@4654.4]
  wire  _T_174; // @[Lookup.scala 9:38:@4656.4]
  wire  _T_178; // @[Lookup.scala 9:38:@4658.4]
  wire  _T_182; // @[Lookup.scala 9:38:@4660.4]
  wire  _T_186; // @[Lookup.scala 9:38:@4662.4]
  wire  _T_190; // @[Lookup.scala 9:38:@4664.4]
  wire  _T_194; // @[Lookup.scala 9:38:@4666.4]
  wire  _T_198; // @[Lookup.scala 9:38:@4668.4]
  wire  _T_202; // @[Lookup.scala 9:38:@4670.4]
  wire  _T_206; // @[Lookup.scala 9:38:@4672.4]
  wire  _T_210; // @[Lookup.scala 9:38:@4674.4]
  wire  _T_212; // @[Lookup.scala 11:37:@4676.4]
  wire  _T_213; // @[Lookup.scala 11:37:@4677.4]
  wire  _T_214; // @[Lookup.scala 11:37:@4678.4]
  wire  _T_215; // @[Lookup.scala 11:37:@4679.4]
  wire  _T_216; // @[Lookup.scala 11:37:@4680.4]
  wire  _T_217; // @[Lookup.scala 11:37:@4681.4]
  wire  _T_218; // @[Lookup.scala 11:37:@4682.4]
  wire  _T_219; // @[Lookup.scala 11:37:@4683.4]
  wire  _T_220; // @[Lookup.scala 11:37:@4684.4]
  wire  _T_221; // @[Lookup.scala 11:37:@4685.4]
  wire  _T_222; // @[Lookup.scala 11:37:@4686.4]
  wire  _T_223; // @[Lookup.scala 11:37:@4687.4]
  wire  _T_224; // @[Lookup.scala 11:37:@4688.4]
  wire  _T_225; // @[Lookup.scala 11:37:@4689.4]
  wire  _T_226; // @[Lookup.scala 11:37:@4690.4]
  wire  _T_227; // @[Lookup.scala 11:37:@4691.4]
  wire  _T_228; // @[Lookup.scala 11:37:@4692.4]
  wire  _T_229; // @[Lookup.scala 11:37:@4693.4]
  wire  _T_230; // @[Lookup.scala 11:37:@4694.4]
  wire  _T_231; // @[Lookup.scala 11:37:@4695.4]
  wire  _T_232; // @[Lookup.scala 11:37:@4696.4]
  wire  _T_233; // @[Lookup.scala 11:37:@4697.4]
  wire  _T_234; // @[Lookup.scala 11:37:@4698.4]
  wire  _T_235; // @[Lookup.scala 11:37:@4699.4]
  wire  _T_236; // @[Lookup.scala 11:37:@4700.4]
  wire  _T_237; // @[Lookup.scala 11:37:@4701.4]
  wire  _T_238; // @[Lookup.scala 11:37:@4702.4]
  wire  _T_239; // @[Lookup.scala 11:37:@4703.4]
  wire  _T_240; // @[Lookup.scala 11:37:@4704.4]
  wire  _T_241; // @[Lookup.scala 11:37:@4705.4]
  wire  _T_242; // @[Lookup.scala 11:37:@4706.4]
  wire  _T_243; // @[Lookup.scala 11:37:@4707.4]
  wire  _T_244; // @[Lookup.scala 11:37:@4708.4]
  wire  _T_245; // @[Lookup.scala 11:37:@4709.4]
  wire  _T_246; // @[Lookup.scala 11:37:@4710.4]
  wire  _T_247; // @[Lookup.scala 11:37:@4711.4]
  wire  _T_248; // @[Lookup.scala 11:37:@4712.4]
  wire  _T_249; // @[Lookup.scala 11:37:@4713.4]
  wire  _T_250; // @[Lookup.scala 11:37:@4714.4]
  wire  _T_251; // @[Lookup.scala 11:37:@4715.4]
  wire  _T_252; // @[Lookup.scala 11:37:@4716.4]
  wire  _T_253; // @[Lookup.scala 11:37:@4717.4]
  wire  _T_254; // @[Lookup.scala 11:37:@4718.4]
  wire  _T_255; // @[Lookup.scala 11:37:@4719.4]
  wire  _T_256; // @[Lookup.scala 11:37:@4720.4]
  wire  _T_257; // @[Lookup.scala 11:37:@4721.4]
  wire  _T_258; // @[Lookup.scala 11:37:@4722.4]
  wire  _T_259; // @[Lookup.scala 11:37:@4723.4]
  wire  signals_0; // @[Lookup.scala 11:37:@4724.4]
  wire [3:0] _T_273; // @[Lookup.scala 11:37:@4738.4]
  wire [3:0] _T_274; // @[Lookup.scala 11:37:@4739.4]
  wire [3:0] _T_275; // @[Lookup.scala 11:37:@4740.4]
  wire [3:0] _T_276; // @[Lookup.scala 11:37:@4741.4]
  wire [3:0] _T_277; // @[Lookup.scala 11:37:@4742.4]
  wire [3:0] _T_278; // @[Lookup.scala 11:37:@4743.4]
  wire [3:0] _T_279; // @[Lookup.scala 11:37:@4744.4]
  wire [3:0] _T_280; // @[Lookup.scala 11:37:@4745.4]
  wire [3:0] _T_281; // @[Lookup.scala 11:37:@4746.4]
  wire [3:0] _T_282; // @[Lookup.scala 11:37:@4747.4]
  wire [3:0] _T_283; // @[Lookup.scala 11:37:@4748.4]
  wire [3:0] _T_284; // @[Lookup.scala 11:37:@4749.4]
  wire [3:0] _T_285; // @[Lookup.scala 11:37:@4750.4]
  wire [3:0] _T_286; // @[Lookup.scala 11:37:@4751.4]
  wire [3:0] _T_287; // @[Lookup.scala 11:37:@4752.4]
  wire [3:0] _T_288; // @[Lookup.scala 11:37:@4753.4]
  wire [3:0] _T_289; // @[Lookup.scala 11:37:@4754.4]
  wire [3:0] _T_290; // @[Lookup.scala 11:37:@4755.4]
  wire [3:0] _T_291; // @[Lookup.scala 11:37:@4756.4]
  wire [3:0] _T_292; // @[Lookup.scala 11:37:@4757.4]
  wire [3:0] _T_293; // @[Lookup.scala 11:37:@4758.4]
  wire [3:0] _T_294; // @[Lookup.scala 11:37:@4759.4]
  wire [3:0] _T_295; // @[Lookup.scala 11:37:@4760.4]
  wire [3:0] _T_296; // @[Lookup.scala 11:37:@4761.4]
  wire [3:0] _T_297; // @[Lookup.scala 11:37:@4762.4]
  wire [3:0] _T_298; // @[Lookup.scala 11:37:@4763.4]
  wire [3:0] _T_299; // @[Lookup.scala 11:37:@4764.4]
  wire [3:0] _T_300; // @[Lookup.scala 11:37:@4765.4]
  wire [3:0] _T_301; // @[Lookup.scala 11:37:@4766.4]
  wire [3:0] _T_302; // @[Lookup.scala 11:37:@4767.4]
  wire [3:0] _T_303; // @[Lookup.scala 11:37:@4768.4]
  wire [3:0] _T_304; // @[Lookup.scala 11:37:@4769.4]
  wire [3:0] _T_305; // @[Lookup.scala 11:37:@4770.4]
  wire [3:0] _T_306; // @[Lookup.scala 11:37:@4771.4]
  wire [3:0] _T_307; // @[Lookup.scala 11:37:@4772.4]
  wire [3:0] _T_308; // @[Lookup.scala 11:37:@4773.4]
  wire [1:0] _T_316; // @[Lookup.scala 11:37:@4782.4]
  wire [1:0] _T_317; // @[Lookup.scala 11:37:@4783.4]
  wire [1:0] _T_318; // @[Lookup.scala 11:37:@4784.4]
  wire [1:0] _T_319; // @[Lookup.scala 11:37:@4785.4]
  wire [1:0] _T_320; // @[Lookup.scala 11:37:@4786.4]
  wire [1:0] _T_321; // @[Lookup.scala 11:37:@4787.4]
  wire [1:0] _T_322; // @[Lookup.scala 11:37:@4788.4]
  wire [1:0] _T_323; // @[Lookup.scala 11:37:@4789.4]
  wire [1:0] _T_324; // @[Lookup.scala 11:37:@4790.4]
  wire [1:0] _T_325; // @[Lookup.scala 11:37:@4791.4]
  wire [1:0] _T_326; // @[Lookup.scala 11:37:@4792.4]
  wire [1:0] _T_327; // @[Lookup.scala 11:37:@4793.4]
  wire [1:0] _T_328; // @[Lookup.scala 11:37:@4794.4]
  wire [1:0] _T_329; // @[Lookup.scala 11:37:@4795.4]
  wire [1:0] _T_330; // @[Lookup.scala 11:37:@4796.4]
  wire [1:0] _T_331; // @[Lookup.scala 11:37:@4797.4]
  wire [1:0] _T_332; // @[Lookup.scala 11:37:@4798.4]
  wire [1:0] _T_333; // @[Lookup.scala 11:37:@4799.4]
  wire [1:0] _T_334; // @[Lookup.scala 11:37:@4800.4]
  wire [1:0] _T_335; // @[Lookup.scala 11:37:@4801.4]
  wire [1:0] _T_336; // @[Lookup.scala 11:37:@4802.4]
  wire [1:0] _T_337; // @[Lookup.scala 11:37:@4803.4]
  wire [1:0] _T_338; // @[Lookup.scala 11:37:@4804.4]
  wire [1:0] _T_339; // @[Lookup.scala 11:37:@4805.4]
  wire [1:0] _T_340; // @[Lookup.scala 11:37:@4806.4]
  wire [1:0] _T_341; // @[Lookup.scala 11:37:@4807.4]
  wire [1:0] _T_342; // @[Lookup.scala 11:37:@4808.4]
  wire [1:0] _T_343; // @[Lookup.scala 11:37:@4809.4]
  wire [1:0] _T_344; // @[Lookup.scala 11:37:@4810.4]
  wire [1:0] _T_345; // @[Lookup.scala 11:37:@4811.4]
  wire [1:0] _T_346; // @[Lookup.scala 11:37:@4812.4]
  wire [1:0] _T_347; // @[Lookup.scala 11:37:@4813.4]
  wire [1:0] _T_348; // @[Lookup.scala 11:37:@4814.4]
  wire [1:0] _T_349; // @[Lookup.scala 11:37:@4815.4]
  wire [1:0] _T_350; // @[Lookup.scala 11:37:@4816.4]
  wire [1:0] _T_351; // @[Lookup.scala 11:37:@4817.4]
  wire [1:0] _T_352; // @[Lookup.scala 11:37:@4818.4]
  wire [1:0] _T_353; // @[Lookup.scala 11:37:@4819.4]
  wire [1:0] _T_354; // @[Lookup.scala 11:37:@4820.4]
  wire [1:0] _T_355; // @[Lookup.scala 11:37:@4821.4]
  wire [1:0] _T_356; // @[Lookup.scala 11:37:@4822.4]
  wire [1:0] _T_357; // @[Lookup.scala 11:37:@4823.4]
  wire [2:0] _T_371; // @[Lookup.scala 11:37:@4838.4]
  wire [2:0] _T_372; // @[Lookup.scala 11:37:@4839.4]
  wire [2:0] _T_373; // @[Lookup.scala 11:37:@4840.4]
  wire [2:0] _T_374; // @[Lookup.scala 11:37:@4841.4]
  wire [2:0] _T_375; // @[Lookup.scala 11:37:@4842.4]
  wire [2:0] _T_376; // @[Lookup.scala 11:37:@4843.4]
  wire [2:0] _T_377; // @[Lookup.scala 11:37:@4844.4]
  wire [2:0] _T_378; // @[Lookup.scala 11:37:@4845.4]
  wire [2:0] _T_379; // @[Lookup.scala 11:37:@4846.4]
  wire [2:0] _T_380; // @[Lookup.scala 11:37:@4847.4]
  wire [2:0] _T_381; // @[Lookup.scala 11:37:@4848.4]
  wire [2:0] _T_382; // @[Lookup.scala 11:37:@4849.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@4850.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@4851.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@4852.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@4853.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@4854.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@4855.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@4856.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@4857.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@4858.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@4859.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@4860.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@4861.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@4862.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@4863.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@4864.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@4865.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@4866.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@4867.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@4868.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@4869.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@4870.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@4871.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@4872.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@4873.4]
  wire  _T_415; // @[Lookup.scala 11:37:@4883.4]
  wire  _T_416; // @[Lookup.scala 11:37:@4884.4]
  wire  _T_417; // @[Lookup.scala 11:37:@4885.4]
  wire  _T_418; // @[Lookup.scala 11:37:@4886.4]
  wire  _T_419; // @[Lookup.scala 11:37:@4887.4]
  wire  _T_420; // @[Lookup.scala 11:37:@4888.4]
  wire  _T_421; // @[Lookup.scala 11:37:@4889.4]
  wire  _T_422; // @[Lookup.scala 11:37:@4890.4]
  wire  _T_423; // @[Lookup.scala 11:37:@4891.4]
  wire  _T_424; // @[Lookup.scala 11:37:@4892.4]
  wire  _T_425; // @[Lookup.scala 11:37:@4893.4]
  wire  _T_426; // @[Lookup.scala 11:37:@4894.4]
  wire  _T_427; // @[Lookup.scala 11:37:@4895.4]
  wire  _T_428; // @[Lookup.scala 11:37:@4896.4]
  wire  _T_429; // @[Lookup.scala 11:37:@4897.4]
  wire  _T_430; // @[Lookup.scala 11:37:@4898.4]
  wire  _T_431; // @[Lookup.scala 11:37:@4899.4]
  wire  _T_432; // @[Lookup.scala 11:37:@4900.4]
  wire  _T_433; // @[Lookup.scala 11:37:@4901.4]
  wire  _T_434; // @[Lookup.scala 11:37:@4902.4]
  wire  _T_435; // @[Lookup.scala 11:37:@4903.4]
  wire  _T_436; // @[Lookup.scala 11:37:@4904.4]
  wire  _T_437; // @[Lookup.scala 11:37:@4905.4]
  wire  _T_438; // @[Lookup.scala 11:37:@4906.4]
  wire  _T_439; // @[Lookup.scala 11:37:@4907.4]
  wire  _T_440; // @[Lookup.scala 11:37:@4908.4]
  wire  _T_441; // @[Lookup.scala 11:37:@4909.4]
  wire  _T_442; // @[Lookup.scala 11:37:@4910.4]
  wire  _T_443; // @[Lookup.scala 11:37:@4911.4]
  wire  _T_444; // @[Lookup.scala 11:37:@4912.4]
  wire  _T_445; // @[Lookup.scala 11:37:@4913.4]
  wire  _T_446; // @[Lookup.scala 11:37:@4914.4]
  wire  _T_447; // @[Lookup.scala 11:37:@4915.4]
  wire  _T_448; // @[Lookup.scala 11:37:@4916.4]
  wire  _T_449; // @[Lookup.scala 11:37:@4917.4]
  wire  _T_450; // @[Lookup.scala 11:37:@4918.4]
  wire  _T_451; // @[Lookup.scala 11:37:@4919.4]
  wire  _T_452; // @[Lookup.scala 11:37:@4920.4]
  wire  _T_453; // @[Lookup.scala 11:37:@4921.4]
  wire  _T_454; // @[Lookup.scala 11:37:@4922.4]
  wire  _T_455; // @[Lookup.scala 11:37:@4923.4]
  wire  _T_475; // @[Lookup.scala 11:37:@4944.4]
  wire  _T_476; // @[Lookup.scala 11:37:@4945.4]
  wire  _T_477; // @[Lookup.scala 11:37:@4946.4]
  wire  _T_478; // @[Lookup.scala 11:37:@4947.4]
  wire  _T_479; // @[Lookup.scala 11:37:@4948.4]
  wire  _T_480; // @[Lookup.scala 11:37:@4949.4]
  wire  _T_481; // @[Lookup.scala 11:37:@4950.4]
  wire  _T_482; // @[Lookup.scala 11:37:@4951.4]
  wire  _T_483; // @[Lookup.scala 11:37:@4952.4]
  wire  _T_484; // @[Lookup.scala 11:37:@4953.4]
  wire  _T_485; // @[Lookup.scala 11:37:@4954.4]
  wire  _T_486; // @[Lookup.scala 11:37:@4955.4]
  wire  _T_487; // @[Lookup.scala 11:37:@4956.4]
  wire  _T_488; // @[Lookup.scala 11:37:@4957.4]
  wire  _T_489; // @[Lookup.scala 11:37:@4958.4]
  wire  _T_490; // @[Lookup.scala 11:37:@4959.4]
  wire  _T_491; // @[Lookup.scala 11:37:@4960.4]
  wire  _T_492; // @[Lookup.scala 11:37:@4961.4]
  wire  _T_493; // @[Lookup.scala 11:37:@4962.4]
  wire  _T_494; // @[Lookup.scala 11:37:@4963.4]
  wire  _T_495; // @[Lookup.scala 11:37:@4964.4]
  wire  _T_496; // @[Lookup.scala 11:37:@4965.4]
  wire  _T_497; // @[Lookup.scala 11:37:@4966.4]
  wire  _T_498; // @[Lookup.scala 11:37:@4967.4]
  wire  _T_499; // @[Lookup.scala 11:37:@4968.4]
  wire  _T_500; // @[Lookup.scala 11:37:@4969.4]
  wire  _T_501; // @[Lookup.scala 11:37:@4970.4]
  wire  _T_502; // @[Lookup.scala 11:37:@4971.4]
  wire  _T_503; // @[Lookup.scala 11:37:@4972.4]
  wire  _T_504; // @[Lookup.scala 11:37:@4973.4]
  wire [3:0] _T_512; // @[Lookup.scala 11:37:@4982.4]
  wire [3:0] _T_513; // @[Lookup.scala 11:37:@4983.4]
  wire [3:0] _T_514; // @[Lookup.scala 11:37:@4984.4]
  wire [3:0] _T_515; // @[Lookup.scala 11:37:@4985.4]
  wire [3:0] _T_516; // @[Lookup.scala 11:37:@4986.4]
  wire [3:0] _T_517; // @[Lookup.scala 11:37:@4987.4]
  wire [3:0] _T_518; // @[Lookup.scala 11:37:@4988.4]
  wire [3:0] _T_519; // @[Lookup.scala 11:37:@4989.4]
  wire [3:0] _T_520; // @[Lookup.scala 11:37:@4990.4]
  wire [3:0] _T_521; // @[Lookup.scala 11:37:@4991.4]
  wire [3:0] _T_522; // @[Lookup.scala 11:37:@4992.4]
  wire [3:0] _T_523; // @[Lookup.scala 11:37:@4993.4]
  wire [3:0] _T_524; // @[Lookup.scala 11:37:@4994.4]
  wire [3:0] _T_525; // @[Lookup.scala 11:37:@4995.4]
  wire [3:0] _T_526; // @[Lookup.scala 11:37:@4996.4]
  wire [3:0] _T_527; // @[Lookup.scala 11:37:@4997.4]
  wire [3:0] _T_528; // @[Lookup.scala 11:37:@4998.4]
  wire [3:0] _T_529; // @[Lookup.scala 11:37:@4999.4]
  wire [3:0] _T_530; // @[Lookup.scala 11:37:@5000.4]
  wire [3:0] _T_531; // @[Lookup.scala 11:37:@5001.4]
  wire [3:0] _T_532; // @[Lookup.scala 11:37:@5002.4]
  wire [3:0] _T_533; // @[Lookup.scala 11:37:@5003.4]
  wire [3:0] _T_534; // @[Lookup.scala 11:37:@5004.4]
  wire [3:0] _T_535; // @[Lookup.scala 11:37:@5005.4]
  wire [3:0] _T_536; // @[Lookup.scala 11:37:@5006.4]
  wire [3:0] _T_537; // @[Lookup.scala 11:37:@5007.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:@5008.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:@5009.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:@5010.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:@5011.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:@5012.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:@5013.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:@5014.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:@5015.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:@5016.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:@5017.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:@5018.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:@5019.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:@5020.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:@5021.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:@5022.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:@5023.4]
  wire [1:0] _T_561; // @[Lookup.scala 11:37:@5032.4]
  wire [1:0] _T_562; // @[Lookup.scala 11:37:@5033.4]
  wire [1:0] _T_563; // @[Lookup.scala 11:37:@5034.4]
  wire [1:0] _T_564; // @[Lookup.scala 11:37:@5035.4]
  wire [1:0] _T_565; // @[Lookup.scala 11:37:@5036.4]
  wire [1:0] _T_566; // @[Lookup.scala 11:37:@5037.4]
  wire [1:0] _T_567; // @[Lookup.scala 11:37:@5038.4]
  wire [1:0] _T_568; // @[Lookup.scala 11:37:@5039.4]
  wire [1:0] _T_569; // @[Lookup.scala 11:37:@5040.4]
  wire [1:0] _T_570; // @[Lookup.scala 11:37:@5041.4]
  wire [1:0] _T_571; // @[Lookup.scala 11:37:@5042.4]
  wire [1:0] _T_572; // @[Lookup.scala 11:37:@5043.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@5044.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@5045.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@5046.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@5047.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@5048.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@5049.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@5050.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@5051.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@5052.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@5053.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@5054.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@5055.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@5056.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@5057.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@5058.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@5059.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@5060.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@5061.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@5062.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@5063.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@5064.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@5065.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@5066.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@5067.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@5068.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@5069.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@5070.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@5071.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@5072.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@5073.4]
  wire  _T_616; // @[Lookup.scala 11:37:@5088.4]
  wire  _T_617; // @[Lookup.scala 11:37:@5089.4]
  wire  _T_618; // @[Lookup.scala 11:37:@5090.4]
  wire  _T_619; // @[Lookup.scala 11:37:@5091.4]
  wire  _T_620; // @[Lookup.scala 11:37:@5092.4]
  wire  _T_621; // @[Lookup.scala 11:37:@5093.4]
  wire  _T_622; // @[Lookup.scala 11:37:@5094.4]
  wire  _T_623; // @[Lookup.scala 11:37:@5095.4]
  wire  _T_624; // @[Lookup.scala 11:37:@5096.4]
  wire  _T_625; // @[Lookup.scala 11:37:@5097.4]
  wire  _T_626; // @[Lookup.scala 11:37:@5098.4]
  wire  _T_627; // @[Lookup.scala 11:37:@5099.4]
  wire  _T_628; // @[Lookup.scala 11:37:@5100.4]
  wire  _T_629; // @[Lookup.scala 11:37:@5101.4]
  wire  _T_630; // @[Lookup.scala 11:37:@5102.4]
  wire  _T_631; // @[Lookup.scala 11:37:@5103.4]
  wire  _T_632; // @[Lookup.scala 11:37:@5104.4]
  wire  _T_633; // @[Lookup.scala 11:37:@5105.4]
  wire  _T_634; // @[Lookup.scala 11:37:@5106.4]
  wire  _T_635; // @[Lookup.scala 11:37:@5107.4]
  wire  _T_636; // @[Lookup.scala 11:37:@5108.4]
  wire  _T_637; // @[Lookup.scala 11:37:@5109.4]
  wire  _T_638; // @[Lookup.scala 11:37:@5110.4]
  wire  _T_639; // @[Lookup.scala 11:37:@5111.4]
  wire  _T_640; // @[Lookup.scala 11:37:@5112.4]
  wire  _T_641; // @[Lookup.scala 11:37:@5113.4]
  wire  _T_642; // @[Lookup.scala 11:37:@5114.4]
  wire  _T_643; // @[Lookup.scala 11:37:@5115.4]
  wire  _T_644; // @[Lookup.scala 11:37:@5116.4]
  wire  _T_645; // @[Lookup.scala 11:37:@5117.4]
  wire  _T_646; // @[Lookup.scala 11:37:@5118.4]
  wire  _T_647; // @[Lookup.scala 11:37:@5119.4]
  wire  _T_648; // @[Lookup.scala 11:37:@5120.4]
  wire  _T_649; // @[Lookup.scala 11:37:@5121.4]
  wire  _T_650; // @[Lookup.scala 11:37:@5122.4]
  wire  _T_651; // @[Lookup.scala 11:37:@5123.4]
  wire  _T_653; // @[Lookup.scala 11:37:@5126.4]
  wire  _T_654; // @[Lookup.scala 11:37:@5127.4]
  wire  _T_655; // @[Lookup.scala 11:37:@5128.4]
  wire  _T_656; // @[Lookup.scala 11:37:@5129.4]
  wire  _T_657; // @[Lookup.scala 11:37:@5130.4]
  wire  _T_658; // @[Lookup.scala 11:37:@5131.4]
  wire  _T_659; // @[Lookup.scala 11:37:@5132.4]
  wire  _T_660; // @[Lookup.scala 11:37:@5133.4]
  wire  _T_661; // @[Lookup.scala 11:37:@5134.4]
  wire  _T_662; // @[Lookup.scala 11:37:@5135.4]
  wire  _T_663; // @[Lookup.scala 11:37:@5136.4]
  wire  _T_664; // @[Lookup.scala 11:37:@5137.4]
  wire  _T_665; // @[Lookup.scala 11:37:@5138.4]
  wire  _T_666; // @[Lookup.scala 11:37:@5139.4]
  wire  _T_667; // @[Lookup.scala 11:37:@5140.4]
  wire  _T_668; // @[Lookup.scala 11:37:@5141.4]
  wire  _T_669; // @[Lookup.scala 11:37:@5142.4]
  wire  _T_670; // @[Lookup.scala 11:37:@5143.4]
  wire  _T_671; // @[Lookup.scala 11:37:@5144.4]
  wire  _T_672; // @[Lookup.scala 11:37:@5145.4]
  wire  _T_673; // @[Lookup.scala 11:37:@5146.4]
  wire  _T_674; // @[Lookup.scala 11:37:@5147.4]
  wire  _T_675; // @[Lookup.scala 11:37:@5148.4]
  wire  _T_676; // @[Lookup.scala 11:37:@5149.4]
  wire  _T_677; // @[Lookup.scala 11:37:@5150.4]
  wire  _T_678; // @[Lookup.scala 11:37:@5151.4]
  wire  _T_679; // @[Lookup.scala 11:37:@5152.4]
  wire  _T_680; // @[Lookup.scala 11:37:@5153.4]
  wire  _T_681; // @[Lookup.scala 11:37:@5154.4]
  wire  _T_682; // @[Lookup.scala 11:37:@5155.4]
  wire  _T_683; // @[Lookup.scala 11:37:@5156.4]
  wire  _T_684; // @[Lookup.scala 11:37:@5157.4]
  wire  _T_685; // @[Lookup.scala 11:37:@5158.4]
  wire  _T_686; // @[Lookup.scala 11:37:@5159.4]
  wire  _T_687; // @[Lookup.scala 11:37:@5160.4]
  wire  _T_688; // @[Lookup.scala 11:37:@5161.4]
  wire  _T_689; // @[Lookup.scala 11:37:@5162.4]
  wire  _T_690; // @[Lookup.scala 11:37:@5163.4]
  wire  _T_691; // @[Lookup.scala 11:37:@5164.4]
  wire  _T_692; // @[Lookup.scala 11:37:@5165.4]
  wire  _T_693; // @[Lookup.scala 11:37:@5166.4]
  wire  _T_694; // @[Lookup.scala 11:37:@5167.4]
  wire  _T_695; // @[Lookup.scala 11:37:@5168.4]
  wire  _T_696; // @[Lookup.scala 11:37:@5169.4]
  wire  _T_697; // @[Lookup.scala 11:37:@5170.4]
  wire  _T_698; // @[Lookup.scala 11:37:@5171.4]
  wire  _T_699; // @[Lookup.scala 11:37:@5172.4]
  wire  _T_700; // @[Lookup.scala 11:37:@5173.4]
  wire  _T_744; // @[Lookup.scala 11:37:@5218.4]
  wire  _T_745; // @[Lookup.scala 11:37:@5219.4]
  wire  _T_746; // @[Lookup.scala 11:37:@5220.4]
  wire  _T_747; // @[Lookup.scala 11:37:@5221.4]
  wire  _T_748; // @[Lookup.scala 11:37:@5222.4]
  wire  _T_749; // @[Lookup.scala 11:37:@5223.4]
  wire [2:0] _T_792; // @[Lookup.scala 11:37:@5267.4]
  wire [2:0] _T_793; // @[Lookup.scala 11:37:@5268.4]
  wire [2:0] _T_794; // @[Lookup.scala 11:37:@5269.4]
  wire [2:0] _T_795; // @[Lookup.scala 11:37:@5270.4]
  wire [2:0] _T_796; // @[Lookup.scala 11:37:@5271.4]
  wire [2:0] _T_797; // @[Lookup.scala 11:37:@5272.4]
  wire [2:0] _T_798; // @[Lookup.scala 11:37:@5273.4]
  wire [2:0] _T_802; // @[Lookup.scala 11:37:@5278.4]
  wire [2:0] _T_803; // @[Lookup.scala 11:37:@5279.4]
  wire [2:0] _T_804; // @[Lookup.scala 11:37:@5280.4]
  wire [2:0] _T_805; // @[Lookup.scala 11:37:@5281.4]
  wire [2:0] _T_806; // @[Lookup.scala 11:37:@5282.4]
  wire [2:0] _T_807; // @[Lookup.scala 11:37:@5283.4]
  wire [2:0] _T_808; // @[Lookup.scala 11:37:@5284.4]
  wire [2:0] _T_809; // @[Lookup.scala 11:37:@5285.4]
  wire [2:0] _T_810; // @[Lookup.scala 11:37:@5286.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@5287.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@5288.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@5289.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@5290.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@5291.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@5292.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@5293.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@5294.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@5295.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@5296.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@5297.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@5298.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@5299.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@5300.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@5301.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@5302.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@5303.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@5304.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@5305.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@5306.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@5307.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@5308.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@5309.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@5310.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@5311.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@5312.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@5313.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@5314.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@5315.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@5316.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@5317.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@5318.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@5319.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@5320.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@5321.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@5322.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@5323.4]
  wire [4:0] _T_899; // @[InstDecoder.scala 130:31:@5390.4]
  wire [4:0] _T_901; // @[InstDecoder.scala 132:31:@5394.4]
  wire [4:0] func; // @[InstDecoder.scala 134:21:@5396.4]
  wire  _T_905; // @[InstDecoder.scala 137:24:@5399.4]
  wire  _T_907; // @[InstDecoder.scala 135:37:@5400.4]
  wire  _T_909; // @[InstDecoder.scala 135:53:@5401.4]
  wire  _T_910; // @[InstDecoder.scala 135:45:@5402.4]
  wire  _T_913; // @[InstDecoder.scala 138:24:@5405.4]
  wire  _T_915; // @[InstDecoder.scala 135:37:@5406.4]
  wire  _T_917; // @[InstDecoder.scala 135:53:@5407.4]
  wire  _T_918; // @[InstDecoder.scala 135:45:@5408.4]
  wire  _T_919; // @[InstDecoder.scala 138:39:@5409.4]
  wire  _T_926; // @[InstDecoder.scala 138:69:@5413.4]
  wire [11:0] imm_itype; // @[InstDecoder.scala 141:27:@5416.4]
  wire [6:0] _T_928; // @[InstDecoder.scala 142:31:@5417.4]
  wire [11:0] imm_stype; // @[Cat.scala 30:58:@5419.4]
  wire  _T_930; // @[InstDecoder.scala 143:31:@5420.4]
  wire  _T_931; // @[InstDecoder.scala 143:44:@5421.4]
  wire [5:0] _T_932; // @[InstDecoder.scala 143:56:@5422.4]
  wire [3:0] _T_933; // @[InstDecoder.scala 143:73:@5423.4]
  wire [11:0] imm_sbtype; // @[Cat.scala 30:58:@5426.4]
  wire [19:0] imm_utype; // @[InstDecoder.scala 144:27:@5427.4]
  wire [7:0] _T_937; // @[InstDecoder.scala 145:44:@5429.4]
  wire  _T_938; // @[InstDecoder.scala 145:60:@5430.4]
  wire [9:0] _T_939; // @[InstDecoder.scala 145:73:@5431.4]
  wire [19:0] imm_ujtype; // @[Cat.scala 30:58:@5434.4]
  wire  _T_942; // @[InstDecoder.scala 148:43:@5435.4]
  wire [19:0] _T_946; // @[Bitwise.scala 72:12:@5437.4]
  wire  _T_948; // @[InstDecoder.scala 149:43:@5440.4]
  wire [19:0] _T_952; // @[Bitwise.scala 72:12:@5442.4]
  wire  _T_954; // @[InstDecoder.scala 150:44:@5445.4]
  wire [18:0] _T_958; // @[Bitwise.scala 72:12:@5447.4]
  wire [30:0] _T_960; // @[Cat.scala 30:58:@5448.4]
  wire  _T_968; // @[InstDecoder.scala 152:44:@5454.4]
  wire [10:0] _T_972; // @[Bitwise.scala 72:12:@5456.4]
  wire [30:0] _T_974; // @[Cat.scala 30:58:@5457.4]
  assign _T_13 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@4575.4]
  assign _T_14 = 32'h2003 == _T_13; // @[Lookup.scala 9:38:@4576.4]
  assign _T_18 = 32'h3 == _T_13; // @[Lookup.scala 9:38:@4578.4]
  assign _T_22 = 32'h4003 == _T_13; // @[Lookup.scala 9:38:@4580.4]
  assign _T_26 = 32'h1003 == _T_13; // @[Lookup.scala 9:38:@4582.4]
  assign _T_30 = 32'h5003 == _T_13; // @[Lookup.scala 9:38:@4584.4]
  assign _T_34 = 32'h2023 == _T_13; // @[Lookup.scala 9:38:@4586.4]
  assign _T_38 = 32'h23 == _T_13; // @[Lookup.scala 9:38:@4588.4]
  assign _T_42 = 32'h1023 == _T_13; // @[Lookup.scala 9:38:@4590.4]
  assign _T_45 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@4591.4]
  assign _T_46 = 32'h17 == _T_45; // @[Lookup.scala 9:38:@4592.4]
  assign _T_50 = 32'h37 == _T_45; // @[Lookup.scala 9:38:@4594.4]
  assign _T_54 = 32'h13 == _T_13; // @[Lookup.scala 9:38:@4596.4]
  assign _T_58 = 32'h7013 == _T_13; // @[Lookup.scala 9:38:@4598.4]
  assign _T_62 = 32'h6013 == _T_13; // @[Lookup.scala 9:38:@4600.4]
  assign _T_66 = 32'h4013 == _T_13; // @[Lookup.scala 9:38:@4602.4]
  assign _T_70 = 32'h2013 == _T_13; // @[Lookup.scala 9:38:@4604.4]
  assign _T_74 = 32'h3013 == _T_13; // @[Lookup.scala 9:38:@4606.4]
  assign _T_77 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@4607.4]
  assign _T_78 = 32'h1013 == _T_77; // @[Lookup.scala 9:38:@4608.4]
  assign _T_82 = 32'h40005013 == _T_77; // @[Lookup.scala 9:38:@4610.4]
  assign _T_86 = 32'h5013 == _T_77; // @[Lookup.scala 9:38:@4612.4]
  assign _T_89 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@4613.4]
  assign _T_90 = 32'h1033 == _T_89; // @[Lookup.scala 9:38:@4614.4]
  assign _T_94 = 32'h33 == _T_89; // @[Lookup.scala 9:38:@4616.4]
  assign _T_98 = 32'h40000033 == _T_89; // @[Lookup.scala 9:38:@4618.4]
  assign _T_102 = 32'h2033 == _T_89; // @[Lookup.scala 9:38:@4620.4]
  assign _T_106 = 32'h3033 == _T_89; // @[Lookup.scala 9:38:@4622.4]
  assign _T_110 = 32'h7033 == _T_89; // @[Lookup.scala 9:38:@4624.4]
  assign _T_114 = 32'h6033 == _T_89; // @[Lookup.scala 9:38:@4626.4]
  assign _T_118 = 32'h4033 == _T_89; // @[Lookup.scala 9:38:@4628.4]
  assign _T_122 = 32'h40005033 == _T_89; // @[Lookup.scala 9:38:@4630.4]
  assign _T_126 = 32'h5033 == _T_89; // @[Lookup.scala 9:38:@4632.4]
  assign _T_130 = 32'h6f == _T_45; // @[Lookup.scala 9:38:@4634.4]
  assign _T_134 = 32'h67 == _T_13; // @[Lookup.scala 9:38:@4636.4]
  assign _T_138 = 32'h63 == _T_13; // @[Lookup.scala 9:38:@4638.4]
  assign _T_142 = 32'h1063 == _T_13; // @[Lookup.scala 9:38:@4640.4]
  assign _T_146 = 32'h5063 == _T_13; // @[Lookup.scala 9:38:@4642.4]
  assign _T_150 = 32'h7063 == _T_13; // @[Lookup.scala 9:38:@4644.4]
  assign _T_154 = 32'h4063 == _T_13; // @[Lookup.scala 9:38:@4646.4]
  assign _T_158 = 32'h6063 == _T_13; // @[Lookup.scala 9:38:@4648.4]
  assign _T_162 = 32'h5073 == _T_13; // @[Lookup.scala 9:38:@4650.4]
  assign _T_166 = 32'h6073 == _T_13; // @[Lookup.scala 9:38:@4652.4]
  assign _T_170 = 32'h1073 == _T_13; // @[Lookup.scala 9:38:@4654.4]
  assign _T_174 = 32'h2073 == _T_13; // @[Lookup.scala 9:38:@4656.4]
  assign _T_178 = 32'h3073 == _T_13; // @[Lookup.scala 9:38:@4658.4]
  assign _T_182 = 32'h7073 == _T_13; // @[Lookup.scala 9:38:@4660.4]
  assign _T_186 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@4662.4]
  assign _T_190 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@4664.4]
  assign _T_194 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@4666.4]
  assign _T_198 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@4668.4]
  assign _T_202 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@4670.4]
  assign _T_206 = 32'h100f == _T_13; // @[Lookup.scala 9:38:@4672.4]
  assign _T_210 = 32'hf == _T_13; // @[Lookup.scala 9:38:@4674.4]
  assign _T_212 = _T_206 ? 1'h1 : _T_210; // @[Lookup.scala 11:37:@4676.4]
  assign _T_213 = _T_202 ? 1'h1 : _T_212; // @[Lookup.scala 11:37:@4677.4]
  assign _T_214 = _T_198 ? 1'h1 : _T_213; // @[Lookup.scala 11:37:@4678.4]
  assign _T_215 = _T_194 ? 1'h1 : _T_214; // @[Lookup.scala 11:37:@4679.4]
  assign _T_216 = _T_190 ? 1'h1 : _T_215; // @[Lookup.scala 11:37:@4680.4]
  assign _T_217 = _T_186 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@4681.4]
  assign _T_218 = _T_182 ? 1'h1 : _T_217; // @[Lookup.scala 11:37:@4682.4]
  assign _T_219 = _T_178 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@4683.4]
  assign _T_220 = _T_174 ? 1'h1 : _T_219; // @[Lookup.scala 11:37:@4684.4]
  assign _T_221 = _T_170 ? 1'h1 : _T_220; // @[Lookup.scala 11:37:@4685.4]
  assign _T_222 = _T_166 ? 1'h1 : _T_221; // @[Lookup.scala 11:37:@4686.4]
  assign _T_223 = _T_162 ? 1'h1 : _T_222; // @[Lookup.scala 11:37:@4687.4]
  assign _T_224 = _T_158 ? 1'h1 : _T_223; // @[Lookup.scala 11:37:@4688.4]
  assign _T_225 = _T_154 ? 1'h1 : _T_224; // @[Lookup.scala 11:37:@4689.4]
  assign _T_226 = _T_150 ? 1'h1 : _T_225; // @[Lookup.scala 11:37:@4690.4]
  assign _T_227 = _T_146 ? 1'h1 : _T_226; // @[Lookup.scala 11:37:@4691.4]
  assign _T_228 = _T_142 ? 1'h1 : _T_227; // @[Lookup.scala 11:37:@4692.4]
  assign _T_229 = _T_138 ? 1'h1 : _T_228; // @[Lookup.scala 11:37:@4693.4]
  assign _T_230 = _T_134 ? 1'h1 : _T_229; // @[Lookup.scala 11:37:@4694.4]
  assign _T_231 = _T_130 ? 1'h1 : _T_230; // @[Lookup.scala 11:37:@4695.4]
  assign _T_232 = _T_126 ? 1'h1 : _T_231; // @[Lookup.scala 11:37:@4696.4]
  assign _T_233 = _T_122 ? 1'h1 : _T_232; // @[Lookup.scala 11:37:@4697.4]
  assign _T_234 = _T_118 ? 1'h1 : _T_233; // @[Lookup.scala 11:37:@4698.4]
  assign _T_235 = _T_114 ? 1'h1 : _T_234; // @[Lookup.scala 11:37:@4699.4]
  assign _T_236 = _T_110 ? 1'h1 : _T_235; // @[Lookup.scala 11:37:@4700.4]
  assign _T_237 = _T_106 ? 1'h1 : _T_236; // @[Lookup.scala 11:37:@4701.4]
  assign _T_238 = _T_102 ? 1'h1 : _T_237; // @[Lookup.scala 11:37:@4702.4]
  assign _T_239 = _T_98 ? 1'h1 : _T_238; // @[Lookup.scala 11:37:@4703.4]
  assign _T_240 = _T_94 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@4704.4]
  assign _T_241 = _T_90 ? 1'h1 : _T_240; // @[Lookup.scala 11:37:@4705.4]
  assign _T_242 = _T_86 ? 1'h1 : _T_241; // @[Lookup.scala 11:37:@4706.4]
  assign _T_243 = _T_82 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@4707.4]
  assign _T_244 = _T_78 ? 1'h1 : _T_243; // @[Lookup.scala 11:37:@4708.4]
  assign _T_245 = _T_74 ? 1'h1 : _T_244; // @[Lookup.scala 11:37:@4709.4]
  assign _T_246 = _T_70 ? 1'h1 : _T_245; // @[Lookup.scala 11:37:@4710.4]
  assign _T_247 = _T_66 ? 1'h1 : _T_246; // @[Lookup.scala 11:37:@4711.4]
  assign _T_248 = _T_62 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@4712.4]
  assign _T_249 = _T_58 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@4713.4]
  assign _T_250 = _T_54 ? 1'h1 : _T_249; // @[Lookup.scala 11:37:@4714.4]
  assign _T_251 = _T_50 ? 1'h1 : _T_250; // @[Lookup.scala 11:37:@4715.4]
  assign _T_252 = _T_46 ? 1'h1 : _T_251; // @[Lookup.scala 11:37:@4716.4]
  assign _T_253 = _T_42 ? 1'h1 : _T_252; // @[Lookup.scala 11:37:@4717.4]
  assign _T_254 = _T_38 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@4718.4]
  assign _T_255 = _T_34 ? 1'h1 : _T_254; // @[Lookup.scala 11:37:@4719.4]
  assign _T_256 = _T_30 ? 1'h1 : _T_255; // @[Lookup.scala 11:37:@4720.4]
  assign _T_257 = _T_26 ? 1'h1 : _T_256; // @[Lookup.scala 11:37:@4721.4]
  assign _T_258 = _T_22 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:@4722.4]
  assign _T_259 = _T_18 ? 1'h1 : _T_258; // @[Lookup.scala 11:37:@4723.4]
  assign signals_0 = _T_14 ? 1'h1 : _T_259; // @[Lookup.scala 11:37:@4724.4]
  assign _T_273 = _T_158 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@4738.4]
  assign _T_274 = _T_154 ? 4'h5 : _T_273; // @[Lookup.scala 11:37:@4739.4]
  assign _T_275 = _T_150 ? 4'h4 : _T_274; // @[Lookup.scala 11:37:@4740.4]
  assign _T_276 = _T_146 ? 4'h3 : _T_275; // @[Lookup.scala 11:37:@4741.4]
  assign _T_277 = _T_142 ? 4'h1 : _T_276; // @[Lookup.scala 11:37:@4742.4]
  assign _T_278 = _T_138 ? 4'h2 : _T_277; // @[Lookup.scala 11:37:@4743.4]
  assign _T_279 = _T_134 ? 4'h8 : _T_278; // @[Lookup.scala 11:37:@4744.4]
  assign _T_280 = _T_130 ? 4'h7 : _T_279; // @[Lookup.scala 11:37:@4745.4]
  assign _T_281 = _T_126 ? 4'h0 : _T_280; // @[Lookup.scala 11:37:@4746.4]
  assign _T_282 = _T_122 ? 4'h0 : _T_281; // @[Lookup.scala 11:37:@4747.4]
  assign _T_283 = _T_118 ? 4'h0 : _T_282; // @[Lookup.scala 11:37:@4748.4]
  assign _T_284 = _T_114 ? 4'h0 : _T_283; // @[Lookup.scala 11:37:@4749.4]
  assign _T_285 = _T_110 ? 4'h0 : _T_284; // @[Lookup.scala 11:37:@4750.4]
  assign _T_286 = _T_106 ? 4'h0 : _T_285; // @[Lookup.scala 11:37:@4751.4]
  assign _T_287 = _T_102 ? 4'h0 : _T_286; // @[Lookup.scala 11:37:@4752.4]
  assign _T_288 = _T_98 ? 4'h0 : _T_287; // @[Lookup.scala 11:37:@4753.4]
  assign _T_289 = _T_94 ? 4'h0 : _T_288; // @[Lookup.scala 11:37:@4754.4]
  assign _T_290 = _T_90 ? 4'h0 : _T_289; // @[Lookup.scala 11:37:@4755.4]
  assign _T_291 = _T_86 ? 4'h0 : _T_290; // @[Lookup.scala 11:37:@4756.4]
  assign _T_292 = _T_82 ? 4'h0 : _T_291; // @[Lookup.scala 11:37:@4757.4]
  assign _T_293 = _T_78 ? 4'h0 : _T_292; // @[Lookup.scala 11:37:@4758.4]
  assign _T_294 = _T_74 ? 4'h0 : _T_293; // @[Lookup.scala 11:37:@4759.4]
  assign _T_295 = _T_70 ? 4'h0 : _T_294; // @[Lookup.scala 11:37:@4760.4]
  assign _T_296 = _T_66 ? 4'h0 : _T_295; // @[Lookup.scala 11:37:@4761.4]
  assign _T_297 = _T_62 ? 4'h0 : _T_296; // @[Lookup.scala 11:37:@4762.4]
  assign _T_298 = _T_58 ? 4'h0 : _T_297; // @[Lookup.scala 11:37:@4763.4]
  assign _T_299 = _T_54 ? 4'h0 : _T_298; // @[Lookup.scala 11:37:@4764.4]
  assign _T_300 = _T_50 ? 4'h0 : _T_299; // @[Lookup.scala 11:37:@4765.4]
  assign _T_301 = _T_46 ? 4'h0 : _T_300; // @[Lookup.scala 11:37:@4766.4]
  assign _T_302 = _T_42 ? 4'h0 : _T_301; // @[Lookup.scala 11:37:@4767.4]
  assign _T_303 = _T_38 ? 4'h0 : _T_302; // @[Lookup.scala 11:37:@4768.4]
  assign _T_304 = _T_34 ? 4'h0 : _T_303; // @[Lookup.scala 11:37:@4769.4]
  assign _T_305 = _T_30 ? 4'h0 : _T_304; // @[Lookup.scala 11:37:@4770.4]
  assign _T_306 = _T_26 ? 4'h0 : _T_305; // @[Lookup.scala 11:37:@4771.4]
  assign _T_307 = _T_22 ? 4'h0 : _T_306; // @[Lookup.scala 11:37:@4772.4]
  assign _T_308 = _T_18 ? 4'h0 : _T_307; // @[Lookup.scala 11:37:@4773.4]
  assign _T_316 = _T_182 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@4782.4]
  assign _T_317 = _T_178 ? 2'h0 : _T_316; // @[Lookup.scala 11:37:@4783.4]
  assign _T_318 = _T_174 ? 2'h0 : _T_317; // @[Lookup.scala 11:37:@4784.4]
  assign _T_319 = _T_170 ? 2'h0 : _T_318; // @[Lookup.scala 11:37:@4785.4]
  assign _T_320 = _T_166 ? 2'h2 : _T_319; // @[Lookup.scala 11:37:@4786.4]
  assign _T_321 = _T_162 ? 2'h2 : _T_320; // @[Lookup.scala 11:37:@4787.4]
  assign _T_322 = _T_158 ? 2'h0 : _T_321; // @[Lookup.scala 11:37:@4788.4]
  assign _T_323 = _T_154 ? 2'h0 : _T_322; // @[Lookup.scala 11:37:@4789.4]
  assign _T_324 = _T_150 ? 2'h0 : _T_323; // @[Lookup.scala 11:37:@4790.4]
  assign _T_325 = _T_146 ? 2'h0 : _T_324; // @[Lookup.scala 11:37:@4791.4]
  assign _T_326 = _T_142 ? 2'h0 : _T_325; // @[Lookup.scala 11:37:@4792.4]
  assign _T_327 = _T_138 ? 2'h0 : _T_326; // @[Lookup.scala 11:37:@4793.4]
  assign _T_328 = _T_134 ? 2'h0 : _T_327; // @[Lookup.scala 11:37:@4794.4]
  assign _T_329 = _T_130 ? 2'h0 : _T_328; // @[Lookup.scala 11:37:@4795.4]
  assign _T_330 = _T_126 ? 2'h0 : _T_329; // @[Lookup.scala 11:37:@4796.4]
  assign _T_331 = _T_122 ? 2'h0 : _T_330; // @[Lookup.scala 11:37:@4797.4]
  assign _T_332 = _T_118 ? 2'h0 : _T_331; // @[Lookup.scala 11:37:@4798.4]
  assign _T_333 = _T_114 ? 2'h0 : _T_332; // @[Lookup.scala 11:37:@4799.4]
  assign _T_334 = _T_110 ? 2'h0 : _T_333; // @[Lookup.scala 11:37:@4800.4]
  assign _T_335 = _T_106 ? 2'h0 : _T_334; // @[Lookup.scala 11:37:@4801.4]
  assign _T_336 = _T_102 ? 2'h0 : _T_335; // @[Lookup.scala 11:37:@4802.4]
  assign _T_337 = _T_98 ? 2'h0 : _T_336; // @[Lookup.scala 11:37:@4803.4]
  assign _T_338 = _T_94 ? 2'h0 : _T_337; // @[Lookup.scala 11:37:@4804.4]
  assign _T_339 = _T_90 ? 2'h0 : _T_338; // @[Lookup.scala 11:37:@4805.4]
  assign _T_340 = _T_86 ? 2'h0 : _T_339; // @[Lookup.scala 11:37:@4806.4]
  assign _T_341 = _T_82 ? 2'h0 : _T_340; // @[Lookup.scala 11:37:@4807.4]
  assign _T_342 = _T_78 ? 2'h0 : _T_341; // @[Lookup.scala 11:37:@4808.4]
  assign _T_343 = _T_74 ? 2'h0 : _T_342; // @[Lookup.scala 11:37:@4809.4]
  assign _T_344 = _T_70 ? 2'h0 : _T_343; // @[Lookup.scala 11:37:@4810.4]
  assign _T_345 = _T_66 ? 2'h0 : _T_344; // @[Lookup.scala 11:37:@4811.4]
  assign _T_346 = _T_62 ? 2'h0 : _T_345; // @[Lookup.scala 11:37:@4812.4]
  assign _T_347 = _T_58 ? 2'h0 : _T_346; // @[Lookup.scala 11:37:@4813.4]
  assign _T_348 = _T_54 ? 2'h0 : _T_347; // @[Lookup.scala 11:37:@4814.4]
  assign _T_349 = _T_50 ? 2'h0 : _T_348; // @[Lookup.scala 11:37:@4815.4]
  assign _T_350 = _T_46 ? 2'h1 : _T_349; // @[Lookup.scala 11:37:@4816.4]
  assign _T_351 = _T_42 ? 2'h0 : _T_350; // @[Lookup.scala 11:37:@4817.4]
  assign _T_352 = _T_38 ? 2'h0 : _T_351; // @[Lookup.scala 11:37:@4818.4]
  assign _T_353 = _T_34 ? 2'h0 : _T_352; // @[Lookup.scala 11:37:@4819.4]
  assign _T_354 = _T_30 ? 2'h0 : _T_353; // @[Lookup.scala 11:37:@4820.4]
  assign _T_355 = _T_26 ? 2'h0 : _T_354; // @[Lookup.scala 11:37:@4821.4]
  assign _T_356 = _T_22 ? 2'h0 : _T_355; // @[Lookup.scala 11:37:@4822.4]
  assign _T_357 = _T_18 ? 2'h0 : _T_356; // @[Lookup.scala 11:37:@4823.4]
  assign _T_371 = _T_158 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37:@4838.4]
  assign _T_372 = _T_154 ? 3'h3 : _T_371; // @[Lookup.scala 11:37:@4839.4]
  assign _T_373 = _T_150 ? 3'h3 : _T_372; // @[Lookup.scala 11:37:@4840.4]
  assign _T_374 = _T_146 ? 3'h3 : _T_373; // @[Lookup.scala 11:37:@4841.4]
  assign _T_375 = _T_142 ? 3'h3 : _T_374; // @[Lookup.scala 11:37:@4842.4]
  assign _T_376 = _T_138 ? 3'h3 : _T_375; // @[Lookup.scala 11:37:@4843.4]
  assign _T_377 = _T_134 ? 3'h1 : _T_376; // @[Lookup.scala 11:37:@4844.4]
  assign _T_378 = _T_130 ? 3'h5 : _T_377; // @[Lookup.scala 11:37:@4845.4]
  assign _T_379 = _T_126 ? 3'h0 : _T_378; // @[Lookup.scala 11:37:@4846.4]
  assign _T_380 = _T_122 ? 3'h0 : _T_379; // @[Lookup.scala 11:37:@4847.4]
  assign _T_381 = _T_118 ? 3'h0 : _T_380; // @[Lookup.scala 11:37:@4848.4]
  assign _T_382 = _T_114 ? 3'h0 : _T_381; // @[Lookup.scala 11:37:@4849.4]
  assign _T_383 = _T_110 ? 3'h0 : _T_382; // @[Lookup.scala 11:37:@4850.4]
  assign _T_384 = _T_106 ? 3'h0 : _T_383; // @[Lookup.scala 11:37:@4851.4]
  assign _T_385 = _T_102 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@4852.4]
  assign _T_386 = _T_98 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@4853.4]
  assign _T_387 = _T_94 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@4854.4]
  assign _T_388 = _T_90 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@4855.4]
  assign _T_389 = _T_86 ? 3'h1 : _T_388; // @[Lookup.scala 11:37:@4856.4]
  assign _T_390 = _T_82 ? 3'h1 : _T_389; // @[Lookup.scala 11:37:@4857.4]
  assign _T_391 = _T_78 ? 3'h1 : _T_390; // @[Lookup.scala 11:37:@4858.4]
  assign _T_392 = _T_74 ? 3'h1 : _T_391; // @[Lookup.scala 11:37:@4859.4]
  assign _T_393 = _T_70 ? 3'h1 : _T_392; // @[Lookup.scala 11:37:@4860.4]
  assign _T_394 = _T_66 ? 3'h1 : _T_393; // @[Lookup.scala 11:37:@4861.4]
  assign _T_395 = _T_62 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@4862.4]
  assign _T_396 = _T_58 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@4863.4]
  assign _T_397 = _T_54 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@4864.4]
  assign _T_398 = _T_50 ? 3'h4 : _T_397; // @[Lookup.scala 11:37:@4865.4]
  assign _T_399 = _T_46 ? 3'h4 : _T_398; // @[Lookup.scala 11:37:@4866.4]
  assign _T_400 = _T_42 ? 3'h2 : _T_399; // @[Lookup.scala 11:37:@4867.4]
  assign _T_401 = _T_38 ? 3'h2 : _T_400; // @[Lookup.scala 11:37:@4868.4]
  assign _T_402 = _T_34 ? 3'h2 : _T_401; // @[Lookup.scala 11:37:@4869.4]
  assign _T_403 = _T_30 ? 3'h1 : _T_402; // @[Lookup.scala 11:37:@4870.4]
  assign _T_404 = _T_26 ? 3'h1 : _T_403; // @[Lookup.scala 11:37:@4871.4]
  assign _T_405 = _T_22 ? 3'h1 : _T_404; // @[Lookup.scala 11:37:@4872.4]
  assign _T_406 = _T_18 ? 3'h1 : _T_405; // @[Lookup.scala 11:37:@4873.4]
  assign _T_415 = _T_178 ? 1'h1 : _T_182; // @[Lookup.scala 11:37:@4883.4]
  assign _T_416 = _T_174 ? 1'h1 : _T_415; // @[Lookup.scala 11:37:@4884.4]
  assign _T_417 = _T_170 ? 1'h1 : _T_416; // @[Lookup.scala 11:37:@4885.4]
  assign _T_418 = _T_166 ? 1'h1 : _T_417; // @[Lookup.scala 11:37:@4886.4]
  assign _T_419 = _T_162 ? 1'h1 : _T_418; // @[Lookup.scala 11:37:@4887.4]
  assign _T_420 = _T_158 ? 1'h1 : _T_419; // @[Lookup.scala 11:37:@4888.4]
  assign _T_421 = _T_154 ? 1'h1 : _T_420; // @[Lookup.scala 11:37:@4889.4]
  assign _T_422 = _T_150 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@4890.4]
  assign _T_423 = _T_146 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@4891.4]
  assign _T_424 = _T_142 ? 1'h1 : _T_423; // @[Lookup.scala 11:37:@4892.4]
  assign _T_425 = _T_138 ? 1'h1 : _T_424; // @[Lookup.scala 11:37:@4893.4]
  assign _T_426 = _T_134 ? 1'h1 : _T_425; // @[Lookup.scala 11:37:@4894.4]
  assign _T_427 = _T_130 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:@4895.4]
  assign _T_428 = _T_126 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@4896.4]
  assign _T_429 = _T_122 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@4897.4]
  assign _T_430 = _T_118 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@4898.4]
  assign _T_431 = _T_114 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@4899.4]
  assign _T_432 = _T_110 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@4900.4]
  assign _T_433 = _T_106 ? 1'h1 : _T_432; // @[Lookup.scala 11:37:@4901.4]
  assign _T_434 = _T_102 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@4902.4]
  assign _T_435 = _T_98 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@4903.4]
  assign _T_436 = _T_94 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@4904.4]
  assign _T_437 = _T_90 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@4905.4]
  assign _T_438 = _T_86 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@4906.4]
  assign _T_439 = _T_82 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@4907.4]
  assign _T_440 = _T_78 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@4908.4]
  assign _T_441 = _T_74 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@4909.4]
  assign _T_442 = _T_70 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@4910.4]
  assign _T_443 = _T_66 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@4911.4]
  assign _T_444 = _T_62 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@4912.4]
  assign _T_445 = _T_58 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@4913.4]
  assign _T_446 = _T_54 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@4914.4]
  assign _T_447 = _T_50 ? 1'h0 : _T_446; // @[Lookup.scala 11:37:@4915.4]
  assign _T_448 = _T_46 ? 1'h0 : _T_447; // @[Lookup.scala 11:37:@4916.4]
  assign _T_449 = _T_42 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@4917.4]
  assign _T_450 = _T_38 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@4918.4]
  assign _T_451 = _T_34 ? 1'h1 : _T_450; // @[Lookup.scala 11:37:@4919.4]
  assign _T_452 = _T_30 ? 1'h1 : _T_451; // @[Lookup.scala 11:37:@4920.4]
  assign _T_453 = _T_26 ? 1'h1 : _T_452; // @[Lookup.scala 11:37:@4921.4]
  assign _T_454 = _T_22 ? 1'h1 : _T_453; // @[Lookup.scala 11:37:@4922.4]
  assign _T_455 = _T_18 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@4923.4]
  assign _T_475 = _T_134 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@4944.4]
  assign _T_476 = _T_130 ? 1'h0 : _T_475; // @[Lookup.scala 11:37:@4945.4]
  assign _T_477 = _T_126 ? 1'h1 : _T_476; // @[Lookup.scala 11:37:@4946.4]
  assign _T_478 = _T_122 ? 1'h1 : _T_477; // @[Lookup.scala 11:37:@4947.4]
  assign _T_479 = _T_118 ? 1'h1 : _T_478; // @[Lookup.scala 11:37:@4948.4]
  assign _T_480 = _T_114 ? 1'h1 : _T_479; // @[Lookup.scala 11:37:@4949.4]
  assign _T_481 = _T_110 ? 1'h1 : _T_480; // @[Lookup.scala 11:37:@4950.4]
  assign _T_482 = _T_106 ? 1'h1 : _T_481; // @[Lookup.scala 11:37:@4951.4]
  assign _T_483 = _T_102 ? 1'h1 : _T_482; // @[Lookup.scala 11:37:@4952.4]
  assign _T_484 = _T_98 ? 1'h1 : _T_483; // @[Lookup.scala 11:37:@4953.4]
  assign _T_485 = _T_94 ? 1'h1 : _T_484; // @[Lookup.scala 11:37:@4954.4]
  assign _T_486 = _T_90 ? 1'h1 : _T_485; // @[Lookup.scala 11:37:@4955.4]
  assign _T_487 = _T_86 ? 1'h0 : _T_486; // @[Lookup.scala 11:37:@4956.4]
  assign _T_488 = _T_82 ? 1'h0 : _T_487; // @[Lookup.scala 11:37:@4957.4]
  assign _T_489 = _T_78 ? 1'h0 : _T_488; // @[Lookup.scala 11:37:@4958.4]
  assign _T_490 = _T_74 ? 1'h0 : _T_489; // @[Lookup.scala 11:37:@4959.4]
  assign _T_491 = _T_70 ? 1'h0 : _T_490; // @[Lookup.scala 11:37:@4960.4]
  assign _T_492 = _T_66 ? 1'h0 : _T_491; // @[Lookup.scala 11:37:@4961.4]
  assign _T_493 = _T_62 ? 1'h0 : _T_492; // @[Lookup.scala 11:37:@4962.4]
  assign _T_494 = _T_58 ? 1'h0 : _T_493; // @[Lookup.scala 11:37:@4963.4]
  assign _T_495 = _T_54 ? 1'h0 : _T_494; // @[Lookup.scala 11:37:@4964.4]
  assign _T_496 = _T_50 ? 1'h0 : _T_495; // @[Lookup.scala 11:37:@4965.4]
  assign _T_497 = _T_46 ? 1'h0 : _T_496; // @[Lookup.scala 11:37:@4966.4]
  assign _T_498 = _T_42 ? 1'h1 : _T_497; // @[Lookup.scala 11:37:@4967.4]
  assign _T_499 = _T_38 ? 1'h1 : _T_498; // @[Lookup.scala 11:37:@4968.4]
  assign _T_500 = _T_34 ? 1'h1 : _T_499; // @[Lookup.scala 11:37:@4969.4]
  assign _T_501 = _T_30 ? 1'h0 : _T_500; // @[Lookup.scala 11:37:@4970.4]
  assign _T_502 = _T_26 ? 1'h0 : _T_501; // @[Lookup.scala 11:37:@4971.4]
  assign _T_503 = _T_22 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@4972.4]
  assign _T_504 = _T_18 ? 1'h0 : _T_503; // @[Lookup.scala 11:37:@4973.4]
  assign _T_512 = _T_182 ? 4'ha : 4'h0; // @[Lookup.scala 11:37:@4982.4]
  assign _T_513 = _T_178 ? 4'ha : _T_512; // @[Lookup.scala 11:37:@4983.4]
  assign _T_514 = _T_174 ? 4'ha : _T_513; // @[Lookup.scala 11:37:@4984.4]
  assign _T_515 = _T_170 ? 4'ha : _T_514; // @[Lookup.scala 11:37:@4985.4]
  assign _T_516 = _T_166 ? 4'ha : _T_515; // @[Lookup.scala 11:37:@4986.4]
  assign _T_517 = _T_162 ? 4'ha : _T_516; // @[Lookup.scala 11:37:@4987.4]
  assign _T_518 = _T_158 ? 4'h0 : _T_517; // @[Lookup.scala 11:37:@4988.4]
  assign _T_519 = _T_154 ? 4'h0 : _T_518; // @[Lookup.scala 11:37:@4989.4]
  assign _T_520 = _T_150 ? 4'h0 : _T_519; // @[Lookup.scala 11:37:@4990.4]
  assign _T_521 = _T_146 ? 4'h0 : _T_520; // @[Lookup.scala 11:37:@4991.4]
  assign _T_522 = _T_142 ? 4'h0 : _T_521; // @[Lookup.scala 11:37:@4992.4]
  assign _T_523 = _T_138 ? 4'h0 : _T_522; // @[Lookup.scala 11:37:@4993.4]
  assign _T_524 = _T_134 ? 4'h0 : _T_523; // @[Lookup.scala 11:37:@4994.4]
  assign _T_525 = _T_130 ? 4'h0 : _T_524; // @[Lookup.scala 11:37:@4995.4]
  assign _T_526 = _T_126 ? 4'h3 : _T_525; // @[Lookup.scala 11:37:@4996.4]
  assign _T_527 = _T_122 ? 4'h4 : _T_526; // @[Lookup.scala 11:37:@4997.4]
  assign _T_528 = _T_118 ? 4'h7 : _T_527; // @[Lookup.scala 11:37:@4998.4]
  assign _T_529 = _T_114 ? 4'h6 : _T_528; // @[Lookup.scala 11:37:@4999.4]
  assign _T_530 = _T_110 ? 4'h5 : _T_529; // @[Lookup.scala 11:37:@5000.4]
  assign _T_531 = _T_106 ? 4'h9 : _T_530; // @[Lookup.scala 11:37:@5001.4]
  assign _T_532 = _T_102 ? 4'h8 : _T_531; // @[Lookup.scala 11:37:@5002.4]
  assign _T_533 = _T_98 ? 4'h1 : _T_532; // @[Lookup.scala 11:37:@5003.4]
  assign _T_534 = _T_94 ? 4'h0 : _T_533; // @[Lookup.scala 11:37:@5004.4]
  assign _T_535 = _T_90 ? 4'h2 : _T_534; // @[Lookup.scala 11:37:@5005.4]
  assign _T_536 = _T_86 ? 4'h3 : _T_535; // @[Lookup.scala 11:37:@5006.4]
  assign _T_537 = _T_82 ? 4'h4 : _T_536; // @[Lookup.scala 11:37:@5007.4]
  assign _T_538 = _T_78 ? 4'h2 : _T_537; // @[Lookup.scala 11:37:@5008.4]
  assign _T_539 = _T_74 ? 4'h9 : _T_538; // @[Lookup.scala 11:37:@5009.4]
  assign _T_540 = _T_70 ? 4'h8 : _T_539; // @[Lookup.scala 11:37:@5010.4]
  assign _T_541 = _T_66 ? 4'h7 : _T_540; // @[Lookup.scala 11:37:@5011.4]
  assign _T_542 = _T_62 ? 4'h6 : _T_541; // @[Lookup.scala 11:37:@5012.4]
  assign _T_543 = _T_58 ? 4'h5 : _T_542; // @[Lookup.scala 11:37:@5013.4]
  assign _T_544 = _T_54 ? 4'h0 : _T_543; // @[Lookup.scala 11:37:@5014.4]
  assign _T_545 = _T_50 ? 4'hb : _T_544; // @[Lookup.scala 11:37:@5015.4]
  assign _T_546 = _T_46 ? 4'h0 : _T_545; // @[Lookup.scala 11:37:@5016.4]
  assign _T_547 = _T_42 ? 4'h0 : _T_546; // @[Lookup.scala 11:37:@5017.4]
  assign _T_548 = _T_38 ? 4'h0 : _T_547; // @[Lookup.scala 11:37:@5018.4]
  assign _T_549 = _T_34 ? 4'h0 : _T_548; // @[Lookup.scala 11:37:@5019.4]
  assign _T_550 = _T_30 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:@5020.4]
  assign _T_551 = _T_26 ? 4'h0 : _T_550; // @[Lookup.scala 11:37:@5021.4]
  assign _T_552 = _T_22 ? 4'h0 : _T_551; // @[Lookup.scala 11:37:@5022.4]
  assign _T_553 = _T_18 ? 4'h0 : _T_552; // @[Lookup.scala 11:37:@5023.4]
  assign _T_561 = _T_182 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@5032.4]
  assign _T_562 = _T_178 ? 2'h3 : _T_561; // @[Lookup.scala 11:37:@5033.4]
  assign _T_563 = _T_174 ? 2'h3 : _T_562; // @[Lookup.scala 11:37:@5034.4]
  assign _T_564 = _T_170 ? 2'h3 : _T_563; // @[Lookup.scala 11:37:@5035.4]
  assign _T_565 = _T_166 ? 2'h3 : _T_564; // @[Lookup.scala 11:37:@5036.4]
  assign _T_566 = _T_162 ? 2'h3 : _T_565; // @[Lookup.scala 11:37:@5037.4]
  assign _T_567 = _T_158 ? 2'h0 : _T_566; // @[Lookup.scala 11:37:@5038.4]
  assign _T_568 = _T_154 ? 2'h0 : _T_567; // @[Lookup.scala 11:37:@5039.4]
  assign _T_569 = _T_150 ? 2'h0 : _T_568; // @[Lookup.scala 11:37:@5040.4]
  assign _T_570 = _T_146 ? 2'h0 : _T_569; // @[Lookup.scala 11:37:@5041.4]
  assign _T_571 = _T_142 ? 2'h0 : _T_570; // @[Lookup.scala 11:37:@5042.4]
  assign _T_572 = _T_138 ? 2'h0 : _T_571; // @[Lookup.scala 11:37:@5043.4]
  assign _T_573 = _T_134 ? 2'h2 : _T_572; // @[Lookup.scala 11:37:@5044.4]
  assign _T_574 = _T_130 ? 2'h2 : _T_573; // @[Lookup.scala 11:37:@5045.4]
  assign _T_575 = _T_126 ? 2'h0 : _T_574; // @[Lookup.scala 11:37:@5046.4]
  assign _T_576 = _T_122 ? 2'h0 : _T_575; // @[Lookup.scala 11:37:@5047.4]
  assign _T_577 = _T_118 ? 2'h0 : _T_576; // @[Lookup.scala 11:37:@5048.4]
  assign _T_578 = _T_114 ? 2'h0 : _T_577; // @[Lookup.scala 11:37:@5049.4]
  assign _T_579 = _T_110 ? 2'h0 : _T_578; // @[Lookup.scala 11:37:@5050.4]
  assign _T_580 = _T_106 ? 2'h0 : _T_579; // @[Lookup.scala 11:37:@5051.4]
  assign _T_581 = _T_102 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@5052.4]
  assign _T_582 = _T_98 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@5053.4]
  assign _T_583 = _T_94 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@5054.4]
  assign _T_584 = _T_90 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@5055.4]
  assign _T_585 = _T_86 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@5056.4]
  assign _T_586 = _T_82 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@5057.4]
  assign _T_587 = _T_78 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@5058.4]
  assign _T_588 = _T_74 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@5059.4]
  assign _T_589 = _T_70 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@5060.4]
  assign _T_590 = _T_66 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@5061.4]
  assign _T_591 = _T_62 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@5062.4]
  assign _T_592 = _T_58 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@5063.4]
  assign _T_593 = _T_54 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@5064.4]
  assign _T_594 = _T_50 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@5065.4]
  assign _T_595 = _T_46 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@5066.4]
  assign _T_596 = _T_42 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@5067.4]
  assign _T_597 = _T_38 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@5068.4]
  assign _T_598 = _T_34 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@5069.4]
  assign _T_599 = _T_30 ? 2'h1 : _T_598; // @[Lookup.scala 11:37:@5070.4]
  assign _T_600 = _T_26 ? 2'h1 : _T_599; // @[Lookup.scala 11:37:@5071.4]
  assign _T_601 = _T_22 ? 2'h1 : _T_600; // @[Lookup.scala 11:37:@5072.4]
  assign _T_602 = _T_18 ? 2'h1 : _T_601; // @[Lookup.scala 11:37:@5073.4]
  assign _T_616 = _T_158 ? 1'h0 : _T_419; // @[Lookup.scala 11:37:@5088.4]
  assign _T_617 = _T_154 ? 1'h0 : _T_616; // @[Lookup.scala 11:37:@5089.4]
  assign _T_618 = _T_150 ? 1'h0 : _T_617; // @[Lookup.scala 11:37:@5090.4]
  assign _T_619 = _T_146 ? 1'h0 : _T_618; // @[Lookup.scala 11:37:@5091.4]
  assign _T_620 = _T_142 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@5092.4]
  assign _T_621 = _T_138 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@5093.4]
  assign _T_622 = _T_134 ? 1'h1 : _T_621; // @[Lookup.scala 11:37:@5094.4]
  assign _T_623 = _T_130 ? 1'h1 : _T_622; // @[Lookup.scala 11:37:@5095.4]
  assign _T_624 = _T_126 ? 1'h1 : _T_623; // @[Lookup.scala 11:37:@5096.4]
  assign _T_625 = _T_122 ? 1'h1 : _T_624; // @[Lookup.scala 11:37:@5097.4]
  assign _T_626 = _T_118 ? 1'h1 : _T_625; // @[Lookup.scala 11:37:@5098.4]
  assign _T_627 = _T_114 ? 1'h1 : _T_626; // @[Lookup.scala 11:37:@5099.4]
  assign _T_628 = _T_110 ? 1'h1 : _T_627; // @[Lookup.scala 11:37:@5100.4]
  assign _T_629 = _T_106 ? 1'h1 : _T_628; // @[Lookup.scala 11:37:@5101.4]
  assign _T_630 = _T_102 ? 1'h1 : _T_629; // @[Lookup.scala 11:37:@5102.4]
  assign _T_631 = _T_98 ? 1'h1 : _T_630; // @[Lookup.scala 11:37:@5103.4]
  assign _T_632 = _T_94 ? 1'h1 : _T_631; // @[Lookup.scala 11:37:@5104.4]
  assign _T_633 = _T_90 ? 1'h1 : _T_632; // @[Lookup.scala 11:37:@5105.4]
  assign _T_634 = _T_86 ? 1'h1 : _T_633; // @[Lookup.scala 11:37:@5106.4]
  assign _T_635 = _T_82 ? 1'h1 : _T_634; // @[Lookup.scala 11:37:@5107.4]
  assign _T_636 = _T_78 ? 1'h1 : _T_635; // @[Lookup.scala 11:37:@5108.4]
  assign _T_637 = _T_74 ? 1'h1 : _T_636; // @[Lookup.scala 11:37:@5109.4]
  assign _T_638 = _T_70 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:@5110.4]
  assign _T_639 = _T_66 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:@5111.4]
  assign _T_640 = _T_62 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:@5112.4]
  assign _T_641 = _T_58 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:@5113.4]
  assign _T_642 = _T_54 ? 1'h1 : _T_641; // @[Lookup.scala 11:37:@5114.4]
  assign _T_643 = _T_50 ? 1'h1 : _T_642; // @[Lookup.scala 11:37:@5115.4]
  assign _T_644 = _T_46 ? 1'h1 : _T_643; // @[Lookup.scala 11:37:@5116.4]
  assign _T_645 = _T_42 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:@5117.4]
  assign _T_646 = _T_38 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:@5118.4]
  assign _T_647 = _T_34 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:@5119.4]
  assign _T_648 = _T_30 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:@5120.4]
  assign _T_649 = _T_26 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:@5121.4]
  assign _T_650 = _T_22 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:@5122.4]
  assign _T_651 = _T_18 ? 1'h1 : _T_650; // @[Lookup.scala 11:37:@5123.4]
  assign _T_653 = _T_206 ? 1'h0 : _T_210; // @[Lookup.scala 11:37:@5126.4]
  assign _T_654 = _T_202 ? 1'h0 : _T_653; // @[Lookup.scala 11:37:@5127.4]
  assign _T_655 = _T_198 ? 1'h0 : _T_654; // @[Lookup.scala 11:37:@5128.4]
  assign _T_656 = _T_194 ? 1'h0 : _T_655; // @[Lookup.scala 11:37:@5129.4]
  assign _T_657 = _T_190 ? 1'h0 : _T_656; // @[Lookup.scala 11:37:@5130.4]
  assign _T_658 = _T_186 ? 1'h0 : _T_657; // @[Lookup.scala 11:37:@5131.4]
  assign _T_659 = _T_182 ? 1'h0 : _T_658; // @[Lookup.scala 11:37:@5132.4]
  assign _T_660 = _T_178 ? 1'h0 : _T_659; // @[Lookup.scala 11:37:@5133.4]
  assign _T_661 = _T_174 ? 1'h0 : _T_660; // @[Lookup.scala 11:37:@5134.4]
  assign _T_662 = _T_170 ? 1'h0 : _T_661; // @[Lookup.scala 11:37:@5135.4]
  assign _T_663 = _T_166 ? 1'h0 : _T_662; // @[Lookup.scala 11:37:@5136.4]
  assign _T_664 = _T_162 ? 1'h0 : _T_663; // @[Lookup.scala 11:37:@5137.4]
  assign _T_665 = _T_158 ? 1'h0 : _T_664; // @[Lookup.scala 11:37:@5138.4]
  assign _T_666 = _T_154 ? 1'h0 : _T_665; // @[Lookup.scala 11:37:@5139.4]
  assign _T_667 = _T_150 ? 1'h0 : _T_666; // @[Lookup.scala 11:37:@5140.4]
  assign _T_668 = _T_146 ? 1'h0 : _T_667; // @[Lookup.scala 11:37:@5141.4]
  assign _T_669 = _T_142 ? 1'h0 : _T_668; // @[Lookup.scala 11:37:@5142.4]
  assign _T_670 = _T_138 ? 1'h0 : _T_669; // @[Lookup.scala 11:37:@5143.4]
  assign _T_671 = _T_134 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:@5144.4]
  assign _T_672 = _T_130 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:@5145.4]
  assign _T_673 = _T_126 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:@5146.4]
  assign _T_674 = _T_122 ? 1'h0 : _T_673; // @[Lookup.scala 11:37:@5147.4]
  assign _T_675 = _T_118 ? 1'h0 : _T_674; // @[Lookup.scala 11:37:@5148.4]
  assign _T_676 = _T_114 ? 1'h0 : _T_675; // @[Lookup.scala 11:37:@5149.4]
  assign _T_677 = _T_110 ? 1'h0 : _T_676; // @[Lookup.scala 11:37:@5150.4]
  assign _T_678 = _T_106 ? 1'h0 : _T_677; // @[Lookup.scala 11:37:@5151.4]
  assign _T_679 = _T_102 ? 1'h0 : _T_678; // @[Lookup.scala 11:37:@5152.4]
  assign _T_680 = _T_98 ? 1'h0 : _T_679; // @[Lookup.scala 11:37:@5153.4]
  assign _T_681 = _T_94 ? 1'h0 : _T_680; // @[Lookup.scala 11:37:@5154.4]
  assign _T_682 = _T_90 ? 1'h0 : _T_681; // @[Lookup.scala 11:37:@5155.4]
  assign _T_683 = _T_86 ? 1'h0 : _T_682; // @[Lookup.scala 11:37:@5156.4]
  assign _T_684 = _T_82 ? 1'h0 : _T_683; // @[Lookup.scala 11:37:@5157.4]
  assign _T_685 = _T_78 ? 1'h0 : _T_684; // @[Lookup.scala 11:37:@5158.4]
  assign _T_686 = _T_74 ? 1'h0 : _T_685; // @[Lookup.scala 11:37:@5159.4]
  assign _T_687 = _T_70 ? 1'h0 : _T_686; // @[Lookup.scala 11:37:@5160.4]
  assign _T_688 = _T_66 ? 1'h0 : _T_687; // @[Lookup.scala 11:37:@5161.4]
  assign _T_689 = _T_62 ? 1'h0 : _T_688; // @[Lookup.scala 11:37:@5162.4]
  assign _T_690 = _T_58 ? 1'h0 : _T_689; // @[Lookup.scala 11:37:@5163.4]
  assign _T_691 = _T_54 ? 1'h0 : _T_690; // @[Lookup.scala 11:37:@5164.4]
  assign _T_692 = _T_50 ? 1'h0 : _T_691; // @[Lookup.scala 11:37:@5165.4]
  assign _T_693 = _T_46 ? 1'h0 : _T_692; // @[Lookup.scala 11:37:@5166.4]
  assign _T_694 = _T_42 ? 1'h1 : _T_693; // @[Lookup.scala 11:37:@5167.4]
  assign _T_695 = _T_38 ? 1'h1 : _T_694; // @[Lookup.scala 11:37:@5168.4]
  assign _T_696 = _T_34 ? 1'h1 : _T_695; // @[Lookup.scala 11:37:@5169.4]
  assign _T_697 = _T_30 ? 1'h1 : _T_696; // @[Lookup.scala 11:37:@5170.4]
  assign _T_698 = _T_26 ? 1'h1 : _T_697; // @[Lookup.scala 11:37:@5171.4]
  assign _T_699 = _T_22 ? 1'h1 : _T_698; // @[Lookup.scala 11:37:@5172.4]
  assign _T_700 = _T_18 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:@5173.4]
  assign _T_744 = _T_38 ? 1'h1 : _T_42; // @[Lookup.scala 11:37:@5218.4]
  assign _T_745 = _T_34 ? 1'h1 : _T_744; // @[Lookup.scala 11:37:@5219.4]
  assign _T_746 = _T_30 ? 1'h0 : _T_745; // @[Lookup.scala 11:37:@5220.4]
  assign _T_747 = _T_26 ? 1'h0 : _T_746; // @[Lookup.scala 11:37:@5221.4]
  assign _T_748 = _T_22 ? 1'h0 : _T_747; // @[Lookup.scala 11:37:@5222.4]
  assign _T_749 = _T_18 ? 1'h0 : _T_748; // @[Lookup.scala 11:37:@5223.4]
  assign _T_792 = _T_42 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@5267.4]
  assign _T_793 = _T_38 ? 3'h1 : _T_792; // @[Lookup.scala 11:37:@5268.4]
  assign _T_794 = _T_34 ? 3'h3 : _T_793; // @[Lookup.scala 11:37:@5269.4]
  assign _T_795 = _T_30 ? 3'h6 : _T_794; // @[Lookup.scala 11:37:@5270.4]
  assign _T_796 = _T_26 ? 3'h2 : _T_795; // @[Lookup.scala 11:37:@5271.4]
  assign _T_797 = _T_22 ? 3'h5 : _T_796; // @[Lookup.scala 11:37:@5272.4]
  assign _T_798 = _T_18 ? 3'h1 : _T_797; // @[Lookup.scala 11:37:@5273.4]
  assign _T_802 = _T_198 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@5278.4]
  assign _T_803 = _T_194 ? 3'h4 : _T_802; // @[Lookup.scala 11:37:@5279.4]
  assign _T_804 = _T_190 ? 3'h4 : _T_803; // @[Lookup.scala 11:37:@5280.4]
  assign _T_805 = _T_186 ? 3'h4 : _T_804; // @[Lookup.scala 11:37:@5281.4]
  assign _T_806 = _T_182 ? 3'h3 : _T_805; // @[Lookup.scala 11:37:@5282.4]
  assign _T_807 = _T_178 ? 3'h3 : _T_806; // @[Lookup.scala 11:37:@5283.4]
  assign _T_808 = _T_174 ? 3'h2 : _T_807; // @[Lookup.scala 11:37:@5284.4]
  assign _T_809 = _T_170 ? 3'h1 : _T_808; // @[Lookup.scala 11:37:@5285.4]
  assign _T_810 = _T_166 ? 3'h2 : _T_809; // @[Lookup.scala 11:37:@5286.4]
  assign _T_811 = _T_162 ? 3'h1 : _T_810; // @[Lookup.scala 11:37:@5287.4]
  assign _T_812 = _T_158 ? 3'h0 : _T_811; // @[Lookup.scala 11:37:@5288.4]
  assign _T_813 = _T_154 ? 3'h0 : _T_812; // @[Lookup.scala 11:37:@5289.4]
  assign _T_814 = _T_150 ? 3'h0 : _T_813; // @[Lookup.scala 11:37:@5290.4]
  assign _T_815 = _T_146 ? 3'h0 : _T_814; // @[Lookup.scala 11:37:@5291.4]
  assign _T_816 = _T_142 ? 3'h0 : _T_815; // @[Lookup.scala 11:37:@5292.4]
  assign _T_817 = _T_138 ? 3'h0 : _T_816; // @[Lookup.scala 11:37:@5293.4]
  assign _T_818 = _T_134 ? 3'h0 : _T_817; // @[Lookup.scala 11:37:@5294.4]
  assign _T_819 = _T_130 ? 3'h0 : _T_818; // @[Lookup.scala 11:37:@5295.4]
  assign _T_820 = _T_126 ? 3'h0 : _T_819; // @[Lookup.scala 11:37:@5296.4]
  assign _T_821 = _T_122 ? 3'h0 : _T_820; // @[Lookup.scala 11:37:@5297.4]
  assign _T_822 = _T_118 ? 3'h0 : _T_821; // @[Lookup.scala 11:37:@5298.4]
  assign _T_823 = _T_114 ? 3'h0 : _T_822; // @[Lookup.scala 11:37:@5299.4]
  assign _T_824 = _T_110 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@5300.4]
  assign _T_825 = _T_106 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@5301.4]
  assign _T_826 = _T_102 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@5302.4]
  assign _T_827 = _T_98 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@5303.4]
  assign _T_828 = _T_94 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@5304.4]
  assign _T_829 = _T_90 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@5305.4]
  assign _T_830 = _T_86 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@5306.4]
  assign _T_831 = _T_82 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@5307.4]
  assign _T_832 = _T_78 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@5308.4]
  assign _T_833 = _T_74 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@5309.4]
  assign _T_834 = _T_70 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@5310.4]
  assign _T_835 = _T_66 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@5311.4]
  assign _T_836 = _T_62 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@5312.4]
  assign _T_837 = _T_58 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@5313.4]
  assign _T_838 = _T_54 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@5314.4]
  assign _T_839 = _T_50 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@5315.4]
  assign _T_840 = _T_46 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@5316.4]
  assign _T_841 = _T_42 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@5317.4]
  assign _T_842 = _T_38 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@5318.4]
  assign _T_843 = _T_34 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@5319.4]
  assign _T_844 = _T_30 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@5320.4]
  assign _T_845 = _T_26 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@5321.4]
  assign _T_846 = _T_22 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@5322.4]
  assign _T_847 = _T_18 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@5323.4]
  assign _T_899 = io_inst[19:15]; // @[InstDecoder.scala 130:31:@5390.4]
  assign _T_901 = io_inst[11:7]; // @[InstDecoder.scala 132:31:@5394.4]
  assign func = io_inst[6:2]; // @[InstDecoder.scala 134:21:@5396.4]
  assign _T_905 = func == 5'h1b; // @[InstDecoder.scala 137:24:@5399.4]
  assign _T_907 = io_cinfo_wbaddr == 5'h1; // @[InstDecoder.scala 135:37:@5400.4]
  assign _T_909 = io_cinfo_wbaddr == 5'h5; // @[InstDecoder.scala 135:53:@5401.4]
  assign _T_910 = _T_907 | _T_909; // @[InstDecoder.scala 135:45:@5402.4]
  assign _T_913 = func == 5'h19; // @[InstDecoder.scala 138:24:@5405.4]
  assign _T_915 = io_cinfo_rs1_addr == 5'h1; // @[InstDecoder.scala 135:37:@5406.4]
  assign _T_917 = io_cinfo_rs1_addr == 5'h5; // @[InstDecoder.scala 135:53:@5407.4]
  assign _T_918 = _T_915 | _T_917; // @[InstDecoder.scala 135:45:@5408.4]
  assign _T_919 = _T_913 & _T_918; // @[InstDecoder.scala 138:39:@5409.4]
  assign _T_926 = _T_910 == 1'h0; // @[InstDecoder.scala 138:69:@5413.4]
  assign imm_itype = io_inst[31:20]; // @[InstDecoder.scala 141:27:@5416.4]
  assign _T_928 = io_inst[31:25]; // @[InstDecoder.scala 142:31:@5417.4]
  assign imm_stype = {_T_928,_T_901}; // @[Cat.scala 30:58:@5419.4]
  assign _T_930 = io_inst[31]; // @[InstDecoder.scala 143:31:@5420.4]
  assign _T_931 = io_inst[7]; // @[InstDecoder.scala 143:44:@5421.4]
  assign _T_932 = io_inst[30:25]; // @[InstDecoder.scala 143:56:@5422.4]
  assign _T_933 = io_inst[11:8]; // @[InstDecoder.scala 143:73:@5423.4]
  assign imm_sbtype = {_T_930,_T_931,_T_932,_T_933}; // @[Cat.scala 30:58:@5426.4]
  assign imm_utype = io_inst[31:12]; // @[InstDecoder.scala 144:27:@5427.4]
  assign _T_937 = io_inst[19:12]; // @[InstDecoder.scala 145:44:@5429.4]
  assign _T_938 = io_inst[20]; // @[InstDecoder.scala 145:60:@5430.4]
  assign _T_939 = io_inst[30:21]; // @[InstDecoder.scala 145:73:@5431.4]
  assign imm_ujtype = {_T_930,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@5434.4]
  assign _T_942 = imm_itype[11]; // @[InstDecoder.scala 148:43:@5435.4]
  assign _T_946 = _T_942 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@5437.4]
  assign _T_948 = imm_stype[11]; // @[InstDecoder.scala 149:43:@5440.4]
  assign _T_952 = _T_948 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@5442.4]
  assign _T_954 = imm_sbtype[11]; // @[InstDecoder.scala 150:44:@5445.4]
  assign _T_958 = _T_954 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@5447.4]
  assign _T_960 = {_T_958,_T_930,_T_931,_T_932,_T_933}; // @[Cat.scala 30:58:@5448.4]
  assign _T_968 = imm_ujtype[19]; // @[InstDecoder.scala 152:44:@5454.4]
  assign _T_972 = _T_968 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@5456.4]
  assign _T_974 = {_T_972,_T_930,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@5457.4]
  assign io_cinfo_br_type = _T_14 ? 4'h0 : _T_308; // @[InstDecoder.scala 115:20:@5375.4]
  assign io_cinfo_op1_sel = _T_14 ? 2'h0 : _T_357; // @[InstDecoder.scala 116:20:@5376.4]
  assign io_cinfo_op2_sel = _T_14 ? 3'h1 : _T_406; // @[InstDecoder.scala 117:20:@5377.4]
  assign io_cinfo_rs1_oen = _T_14 ? 1'h1 : _T_455; // @[InstDecoder.scala 118:20:@5378.4]
  assign io_cinfo_rs2_oen = _T_14 ? 1'h0 : _T_504; // @[InstDecoder.scala 119:20:@5379.4]
  assign io_cinfo_alu_fun = _T_14 ? 4'h0 : _T_553; // @[InstDecoder.scala 120:20:@5380.4]
  assign io_cinfo_wb_sel = _T_14 ? 2'h1 : _T_602; // @[InstDecoder.scala 121:20:@5381.4]
  assign io_cinfo_rf_wen = _T_14 ? 1'h1 : _T_651; // @[InstDecoder.scala 122:20:@5382.4]
  assign io_cinfo_mem_en = _T_14 ? 1'h1 : _T_700; // @[InstDecoder.scala 123:20:@5383.4]
  assign io_cinfo_mem_fcn = _T_14 ? 1'h0 : _T_749; // @[InstDecoder.scala 124:20:@5384.4]
  assign io_cinfo_mem_typ = _T_14 ? 3'h3 : _T_798; // @[InstDecoder.scala 125:20:@5385.4]
  assign io_cinfo_csr_cmd = _T_14 ? 3'h0 : _T_847; // @[InstDecoder.scala 126:20:@5386.4]
  assign io_cinfo_illegal = signals_0 == 1'h0; // @[InstDecoder.scala 127:20:@5388.4]
  assign io_cinfo_is_branch = func == 5'h18; // @[InstDecoder.scala 136:22:@5398.4]
  assign io_cinfo_jal = _T_905 & _T_910; // @[InstDecoder.scala 137:16:@5404.4]
  assign io_cinfo_ret = _T_919 & _T_926; // @[InstDecoder.scala 138:16:@5415.4]
  assign io_cinfo_rs1_addr = io_inst[19:15]; // @[InstDecoder.scala 130:21:@5391.4]
  assign io_cinfo_rs2_addr = io_inst[24:20]; // @[InstDecoder.scala 131:21:@5393.4]
  assign io_cinfo_wbaddr = io_inst[11:7]; // @[InstDecoder.scala 132:21:@5395.4]
  assign io_dinfo_imm_i = {_T_946,imm_itype}; // @[InstDecoder.scala 148:19:@5439.4]
  assign io_dinfo_imm_s = {_T_952,imm_stype}; // @[InstDecoder.scala 149:19:@5444.4]
  assign io_dinfo_imm_sb = {_T_960,1'h0}; // @[InstDecoder.scala 150:19:@5450.4]
  assign io_dinfo_imm_u = {imm_utype,12'h0}; // @[InstDecoder.scala 151:19:@5453.4]
  assign io_dinfo_imm_uj = {_T_974,1'h0}; // @[InstDecoder.scala 152:19:@5459.4]
  assign io_dinfo_imm_z = {27'h0,_T_899}; // @[InstDecoder.scala 153:19:@5463.4]
endmodule
module Regfile( // @[:@5465.2]
  input         clock, // @[:@5466.4]
  input  [4:0]  io_rs1_addr, // @[:@5468.4]
  output [31:0] io_rs1_data, // @[:@5468.4]
  input  [4:0]  io_rs2_addr, // @[:@5468.4]
  output [31:0] io_rs2_data, // @[:@5468.4]
  input  [4:0]  io_waddr, // @[:@5468.4]
  input  [31:0] io_wdata, // @[:@5468.4]
  input         io_wen // @[:@5468.4]
);
  reg [31:0] regfile [0:31]; // @[Regfile.scala 27:21:@5470.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_27_data; // @[Regfile.scala 27:21:@5470.4]
  wire [4:0] regfile__T_27_addr; // @[Regfile.scala 27:21:@5470.4]
  wire [31:0] regfile__T_32_data; // @[Regfile.scala 27:21:@5470.4]
  wire [4:0] regfile__T_32_addr; // @[Regfile.scala 27:21:@5470.4]
  wire [31:0] regfile__T_24_data; // @[Regfile.scala 27:21:@5470.4]
  wire [4:0] regfile__T_24_addr; // @[Regfile.scala 27:21:@5470.4]
  wire  regfile__T_24_mask; // @[Regfile.scala 27:21:@5470.4]
  wire  regfile__T_24_en; // @[Regfile.scala 27:21:@5470.4]
  wire  _T_22; // @[Regfile.scala 29:30:@5471.4]
  wire  _T_26; // @[Regfile.scala 34:35:@5477.4]
  wire  _T_31; // @[Regfile.scala 35:35:@5481.4]
  assign regfile__T_27_addr = io_rs1_addr;
  assign regfile__T_27_data = regfile[regfile__T_27_addr]; // @[Regfile.scala 27:21:@5470.4]
  assign regfile__T_32_addr = io_rs2_addr;
  assign regfile__T_32_data = regfile[regfile__T_32_addr]; // @[Regfile.scala 27:21:@5470.4]
  assign regfile__T_24_data = io_wdata;
  assign regfile__T_24_addr = io_waddr;
  assign regfile__T_24_mask = 1'h1;
  assign regfile__T_24_en = io_wen & _T_22;
  assign _T_22 = io_waddr != 5'h0; // @[Regfile.scala 29:30:@5471.4]
  assign _T_26 = io_rs1_addr != 5'h0; // @[Regfile.scala 34:35:@5477.4]
  assign _T_31 = io_rs2_addr != 5'h0; // @[Regfile.scala 35:35:@5481.4]
  assign io_rs1_data = _T_26 ? regfile__T_27_data : 32'h0; // @[Regfile.scala 34:16:@5480.4]
  assign io_rs2_data = _T_31 ? regfile__T_32_data : 32'h0; // @[Regfile.scala 35:16:@5484.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(regfile__T_24_en & regfile__T_24_mask) begin
      regfile[regfile__T_24_addr] <= regfile__T_24_data; // @[Regfile.scala 27:21:@5470.4]
    end
  end
endmodule
module ALU( // @[:@5486.2]
  input  [31:0] io_op1, // @[:@5489.4]
  input  [31:0] io_op2, // @[:@5489.4]
  input  [31:0] io_pc, // @[:@5489.4]
  input  [3:0]  io_ctrl_fun, // @[:@5489.4]
  input  [3:0]  io_ctrl_br_type, // @[:@5489.4]
  input  [1:0]  io_ctrl_wb_sel, // @[:@5489.4]
  output [1:0]  io_ctrl_pc_sel, // @[:@5489.4]
  input  [31:0] io_rs2_data, // @[:@5489.4]
  output [31:0] io_result, // @[:@5489.4]
  output [31:0] io_target_brjmp, // @[:@5489.4]
  output [31:0] io_target_jpreg, // @[:@5489.4]
  output [31:0] io_target_conti // @[:@5489.4]
);
  wire [4:0] alu_shamt; // @[ALU.scala 32:32:@5491.4]
  wire [32:0] _T_25; // @[ALU.scala 33:34:@5492.4]
  wire [31:0] add_result; // @[ALU.scala 33:34:@5493.4]
  wire  _T_29; // @[ALU.scala 38:18:@5496.4]
  wire  _T_30; // @[ALU.scala 39:18:@5497.4]
  wire [32:0] _T_31; // @[ALU.scala 39:44:@5498.4]
  wire [32:0] _T_32; // @[ALU.scala 39:44:@5499.4]
  wire [31:0] _T_33; // @[ALU.scala 39:44:@5500.4]
  wire  _T_34; // @[ALU.scala 40:18:@5501.4]
  wire [31:0] _T_35; // @[ALU.scala 40:44:@5502.4]
  wire  _T_36; // @[ALU.scala 41:18:@5503.4]
  wire [31:0] _T_37; // @[ALU.scala 41:44:@5504.4]
  wire  _T_38; // @[ALU.scala 42:18:@5505.4]
  wire [31:0] _T_39; // @[ALU.scala 42:44:@5506.4]
  wire  _T_40; // @[ALU.scala 43:18:@5507.4]
  wire [31:0] _T_41; // @[ALU.scala 43:44:@5508.4]
  wire [31:0] _T_42; // @[ALU.scala 43:60:@5509.4]
  wire  _T_43; // @[ALU.scala 43:51:@5510.4]
  wire  _T_44; // @[ALU.scala 44:18:@5511.4]
  wire  _T_45; // @[ALU.scala 44:44:@5512.4]
  wire  _T_46; // @[ALU.scala 45:18:@5513.4]
  wire [62:0] _GEN_0; // @[ALU.scala 45:44:@5514.4]
  wire [62:0] _T_47; // @[ALU.scala 45:44:@5514.4]
  wire [31:0] _T_48; // @[ALU.scala 45:57:@5515.4]
  wire  _T_49; // @[ALU.scala 46:18:@5516.4]
  wire [31:0] _T_51; // @[ALU.scala 46:51:@5518.4]
  wire [31:0] _T_52; // @[ALU.scala 46:65:@5519.4]
  wire  _T_53; // @[ALU.scala 47:18:@5520.4]
  wire [31:0] _T_54; // @[ALU.scala 47:44:@5521.4]
  wire  _T_55; // @[ALU.scala 48:18:@5522.4]
  wire  _T_56; // @[ALU.scala 49:18:@5523.4]
  wire [31:0] _T_57; // @[Mux.scala 61:16:@5524.4]
  wire [31:0] _T_58; // @[Mux.scala 61:16:@5525.4]
  wire [31:0] _T_59; // @[Mux.scala 61:16:@5526.4]
  wire [31:0] _T_60; // @[Mux.scala 61:16:@5527.4]
  wire [31:0] _T_61; // @[Mux.scala 61:16:@5528.4]
  wire [31:0] _T_62; // @[Mux.scala 61:16:@5529.4]
  wire [31:0] _T_63; // @[Mux.scala 61:16:@5530.4]
  wire [31:0] _T_64; // @[Mux.scala 61:16:@5531.4]
  wire [31:0] _T_65; // @[Mux.scala 61:16:@5532.4]
  wire [31:0] _T_66; // @[Mux.scala 61:16:@5533.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@5534.4]
  wire [31:0] result; // @[Mux.scala 61:16:@5535.4]
  wire [32:0] _T_69; // @[ALU.scala 52:31:@5537.4]
  wire [30:0] _T_71; // @[ALU.scala 53:39:@5540.4]
  wire [32:0] _T_75; // @[ALU.scala 54:31:@5543.4]
  wire  _T_77; // @[ALU.scala 55:40:@5546.4]
  wire  br_eq; // @[ALU.scala 57:29:@5549.4]
  wire [31:0] _T_80; // @[ALU.scala 58:50:@5551.4]
  wire  br_lt; // @[ALU.scala 58:36:@5552.4]
  wire  br_ltu; // @[ALU.scala 59:36:@5553.4]
  wire  _T_81; // @[ALU.scala 63:25:@5554.4]
  wire  _T_82; // @[ALU.scala 64:25:@5555.4]
  wire  _T_84; // @[ALU.scala 64:41:@5556.4]
  wire [1:0] _T_85; // @[ALU.scala 64:40:@5557.4]
  wire  _T_86; // @[ALU.scala 65:25:@5558.4]
  wire [1:0] _T_87; // @[ALU.scala 65:40:@5559.4]
  wire  _T_88; // @[ALU.scala 66:25:@5560.4]
  wire  _T_90; // @[ALU.scala 66:41:@5561.4]
  wire [1:0] _T_91; // @[ALU.scala 66:40:@5562.4]
  wire  _T_92; // @[ALU.scala 67:25:@5563.4]
  wire  _T_94; // @[ALU.scala 67:41:@5564.4]
  wire [1:0] _T_95; // @[ALU.scala 67:40:@5565.4]
  wire  _T_96; // @[ALU.scala 68:25:@5566.4]
  wire [1:0] _T_97; // @[ALU.scala 68:40:@5567.4]
  wire  _T_98; // @[ALU.scala 69:25:@5568.4]
  wire [1:0] _T_99; // @[ALU.scala 69:40:@5569.4]
  wire  _T_100; // @[ALU.scala 70:25:@5570.4]
  wire  _T_101; // @[ALU.scala 71:25:@5571.4]
  wire [1:0] _T_102; // @[ALU.scala 71:8:@5572.4]
  wire [1:0] _T_103; // @[ALU.scala 70:8:@5573.4]
  wire [1:0] _T_104; // @[ALU.scala 69:8:@5574.4]
  wire [1:0] _T_105; // @[ALU.scala 68:8:@5575.4]
  wire [1:0] _T_106; // @[ALU.scala 67:8:@5576.4]
  wire [1:0] _T_107; // @[ALU.scala 66:8:@5577.4]
  wire [1:0] _T_108; // @[ALU.scala 65:8:@5578.4]
  wire [1:0] _T_109; // @[ALU.scala 64:8:@5579.4]
  assign alu_shamt = io_op2[4:0]; // @[ALU.scala 32:32:@5491.4]
  assign _T_25 = io_op1 + io_op2; // @[ALU.scala 33:34:@5492.4]
  assign add_result = io_op1 + io_op2; // @[ALU.scala 33:34:@5493.4]
  assign _T_29 = io_ctrl_fun == 4'h0; // @[ALU.scala 38:18:@5496.4]
  assign _T_30 = io_ctrl_fun == 4'h1; // @[ALU.scala 39:18:@5497.4]
  assign _T_31 = io_op1 - io_op2; // @[ALU.scala 39:44:@5498.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 39:44:@5499.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 39:44:@5500.4]
  assign _T_34 = io_ctrl_fun == 4'h5; // @[ALU.scala 40:18:@5501.4]
  assign _T_35 = io_op1 & io_op2; // @[ALU.scala 40:44:@5502.4]
  assign _T_36 = io_ctrl_fun == 4'h6; // @[ALU.scala 41:18:@5503.4]
  assign _T_37 = io_op1 | io_op2; // @[ALU.scala 41:44:@5504.4]
  assign _T_38 = io_ctrl_fun == 4'h7; // @[ALU.scala 42:18:@5505.4]
  assign _T_39 = io_op1 ^ io_op2; // @[ALU.scala 42:44:@5506.4]
  assign _T_40 = io_ctrl_fun == 4'h8; // @[ALU.scala 43:18:@5507.4]
  assign _T_41 = $signed(io_op1); // @[ALU.scala 43:44:@5508.4]
  assign _T_42 = $signed(io_op2); // @[ALU.scala 43:60:@5509.4]
  assign _T_43 = $signed(_T_41) < $signed(_T_42); // @[ALU.scala 43:51:@5510.4]
  assign _T_44 = io_ctrl_fun == 4'h9; // @[ALU.scala 44:18:@5511.4]
  assign _T_45 = io_op1 < io_op2; // @[ALU.scala 44:44:@5512.4]
  assign _T_46 = io_ctrl_fun == 4'h2; // @[ALU.scala 45:18:@5513.4]
  assign _GEN_0 = {{31'd0}, io_op1}; // @[ALU.scala 45:44:@5514.4]
  assign _T_47 = _GEN_0 << alu_shamt; // @[ALU.scala 45:44:@5514.4]
  assign _T_48 = _T_47[31:0]; // @[ALU.scala 45:57:@5515.4]
  assign _T_49 = io_ctrl_fun == 4'h4; // @[ALU.scala 46:18:@5516.4]
  assign _T_51 = $signed(_T_41) >>> alu_shamt; // @[ALU.scala 46:51:@5518.4]
  assign _T_52 = $unsigned(_T_51); // @[ALU.scala 46:65:@5519.4]
  assign _T_53 = io_ctrl_fun == 4'h3; // @[ALU.scala 47:18:@5520.4]
  assign _T_54 = io_op1 >> alu_shamt; // @[ALU.scala 47:44:@5521.4]
  assign _T_55 = io_ctrl_fun == 4'ha; // @[ALU.scala 48:18:@5522.4]
  assign _T_56 = io_ctrl_fun == 4'hb; // @[ALU.scala 49:18:@5523.4]
  assign _T_57 = _T_56 ? io_op2 : 32'h0; // @[Mux.scala 61:16:@5524.4]
  assign _T_58 = _T_55 ? io_op1 : _T_57; // @[Mux.scala 61:16:@5525.4]
  assign _T_59 = _T_53 ? _T_54 : _T_58; // @[Mux.scala 61:16:@5526.4]
  assign _T_60 = _T_49 ? _T_52 : _T_59; // @[Mux.scala 61:16:@5527.4]
  assign _T_61 = _T_46 ? _T_48 : _T_60; // @[Mux.scala 61:16:@5528.4]
  assign _T_62 = _T_44 ? {{31'd0}, _T_45} : _T_61; // @[Mux.scala 61:16:@5529.4]
  assign _T_63 = _T_40 ? {{31'd0}, _T_43} : _T_62; // @[Mux.scala 61:16:@5530.4]
  assign _T_64 = _T_38 ? _T_39 : _T_63; // @[Mux.scala 61:16:@5531.4]
  assign _T_65 = _T_36 ? _T_37 : _T_64; // @[Mux.scala 61:16:@5532.4]
  assign _T_66 = _T_34 ? _T_35 : _T_65; // @[Mux.scala 61:16:@5533.4]
  assign _T_67 = _T_30 ? _T_33 : _T_66; // @[Mux.scala 61:16:@5534.4]
  assign result = _T_29 ? add_result : _T_67; // @[Mux.scala 61:16:@5535.4]
  assign _T_69 = io_pc + io_op2; // @[ALU.scala 52:31:@5537.4]
  assign _T_71 = add_result[31:1]; // @[ALU.scala 53:39:@5540.4]
  assign _T_75 = io_pc + 32'h4; // @[ALU.scala 54:31:@5543.4]
  assign _T_77 = io_ctrl_wb_sel == 2'h2; // @[ALU.scala 55:40:@5546.4]
  assign br_eq = io_op1 == io_rs2_data; // @[ALU.scala 57:29:@5549.4]
  assign _T_80 = $signed(io_rs2_data); // @[ALU.scala 58:50:@5551.4]
  assign br_lt = $signed(_T_41) < $signed(_T_80); // @[ALU.scala 58:36:@5552.4]
  assign br_ltu = io_op1 < io_rs2_data; // @[ALU.scala 59:36:@5553.4]
  assign _T_81 = io_ctrl_br_type == 4'h0; // @[ALU.scala 63:25:@5554.4]
  assign _T_82 = io_ctrl_br_type == 4'h1; // @[ALU.scala 64:25:@5555.4]
  assign _T_84 = br_eq == 1'h0; // @[ALU.scala 64:41:@5556.4]
  assign _T_85 = _T_84 ? 2'h1 : 2'h0; // @[ALU.scala 64:40:@5557.4]
  assign _T_86 = io_ctrl_br_type == 4'h2; // @[ALU.scala 65:25:@5558.4]
  assign _T_87 = br_eq ? 2'h1 : 2'h0; // @[ALU.scala 65:40:@5559.4]
  assign _T_88 = io_ctrl_br_type == 4'h3; // @[ALU.scala 66:25:@5560.4]
  assign _T_90 = br_lt == 1'h0; // @[ALU.scala 66:41:@5561.4]
  assign _T_91 = _T_90 ? 2'h1 : 2'h0; // @[ALU.scala 66:40:@5562.4]
  assign _T_92 = io_ctrl_br_type == 4'h4; // @[ALU.scala 67:25:@5563.4]
  assign _T_94 = br_ltu == 1'h0; // @[ALU.scala 67:41:@5564.4]
  assign _T_95 = _T_94 ? 2'h1 : 2'h0; // @[ALU.scala 67:40:@5565.4]
  assign _T_96 = io_ctrl_br_type == 4'h5; // @[ALU.scala 68:25:@5566.4]
  assign _T_97 = br_lt ? 2'h1 : 2'h0; // @[ALU.scala 68:40:@5567.4]
  assign _T_98 = io_ctrl_br_type == 4'h6; // @[ALU.scala 69:25:@5568.4]
  assign _T_99 = br_ltu ? 2'h1 : 2'h0; // @[ALU.scala 69:40:@5569.4]
  assign _T_100 = io_ctrl_br_type == 4'h7; // @[ALU.scala 70:25:@5570.4]
  assign _T_101 = io_ctrl_br_type == 4'h8; // @[ALU.scala 71:25:@5571.4]
  assign _T_102 = _T_101 ? 2'h2 : 2'h0; // @[ALU.scala 71:8:@5572.4]
  assign _T_103 = _T_100 ? 2'h1 : _T_102; // @[ALU.scala 70:8:@5573.4]
  assign _T_104 = _T_98 ? _T_99 : _T_103; // @[ALU.scala 69:8:@5574.4]
  assign _T_105 = _T_96 ? _T_97 : _T_104; // @[ALU.scala 68:8:@5575.4]
  assign _T_106 = _T_92 ? _T_95 : _T_105; // @[ALU.scala 67:8:@5576.4]
  assign _T_107 = _T_88 ? _T_91 : _T_106; // @[ALU.scala 66:8:@5577.4]
  assign _T_108 = _T_86 ? _T_87 : _T_107; // @[ALU.scala 65:8:@5578.4]
  assign _T_109 = _T_82 ? _T_85 : _T_108; // @[ALU.scala 64:8:@5579.4]
  assign io_ctrl_pc_sel = _T_81 ? 2'h0 : _T_109; // @[ALU.scala 62:18:@5581.4]
  assign io_result = _T_77 ? io_target_conti : result; // @[ALU.scala 55:18:@5548.4]
  assign io_target_brjmp = io_pc + io_op2; // @[ALU.scala 52:22:@5539.4]
  assign io_target_jpreg = {_T_71,1'h0}; // @[ALU.scala 53:22:@5542.4]
  assign io_target_conti = io_pc + 32'h4; // @[ALU.scala 54:22:@5545.4]
endmodule
module BackEnd( // @[:@5583.2]
  input         clock, // @[:@5584.4]
  input         reset, // @[:@5585.4]
  output        io_mem_req_valid, // @[:@5586.4]
  output [31:0] io_mem_req_bits_addr, // @[:@5586.4]
  output [31:0] io_mem_req_bits_data, // @[:@5586.4]
  output        io_mem_req_bits_fcn, // @[:@5586.4]
  output [2:0]  io_mem_req_bits_typ, // @[:@5586.4]
  input         io_mem_resp_valid, // @[:@5586.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@5586.4]
  output [31:0] io_cyc, // @[:@5586.4]
  output        io_front_xcpt_valid, // @[:@5586.4]
  output [31:0] io_front_xcpt_bits, // @[:@5586.4]
  output        io_front_kill, // @[:@5586.4]
  output        io_front_forward, // @[:@5586.4]
  input         io_front_inst_valid, // @[:@5586.4]
  input  [31:0] io_front_inst_bits, // @[:@5586.4]
  input  [31:0] io_front_pc, // @[:@5586.4]
  input  [9:0]  io_front_pred_history, // @[:@5586.4]
  input         io_front_pred_diff, // @[:@5586.4]
  input  [31:0] io_front_pred_tgt, // @[:@5586.4]
  output        io_front_ras_pop, // @[:@5586.4]
  output        io_front_ras_push_valid, // @[:@5586.4]
  output [31:0] io_front_ras_push_bits, // @[:@5586.4]
  output [31:0] io_front_fb_pc, // @[:@5586.4]
  output [1:0]  io_front_fb_type, // @[:@5586.4]
  output        io_front_feedBack_redirect, // @[:@5586.4]
  output [9:0]  io_front_feedBack_history, // @[:@5586.4]
  output        io_front_feedBack_diff, // @[:@5586.4]
  output [31:0] io_front_feedBack_tgt, // @[:@5586.4]
  output        io_front_feedBack_valid // @[:@5586.4]
);
  wire  csr_clock; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_reset; // @[BackEnd.scala 81:19:@5588.4]
  wire [2:0] csr_io_rw_cmd; // @[BackEnd.scala 81:19:@5588.4]
  wire [11:0] csr_io_rw_addr; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_rw_rdata; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_rw_wdata; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_eret; // @[BackEnd.scala 81:19:@5588.4]
  wire [1:0] csr_io_status_prv; // @[BackEnd.scala 81:19:@5588.4]
  wire [13:0] csr_io_status_unimp5; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_status_mprv; // @[BackEnd.scala 81:19:@5588.4]
  wire [1:0] csr_io_status_unimp4; // @[BackEnd.scala 81:19:@5588.4]
  wire [1:0] csr_io_status_mpp; // @[BackEnd.scala 81:19:@5588.4]
  wire [2:0] csr_io_status_unimp3; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_status_mpie; // @[BackEnd.scala 81:19:@5588.4]
  wire [2:0] csr_io_status_unimp2; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_status_mie; // @[BackEnd.scala 81:19:@5588.4]
  wire [2:0] csr_io_status_unimp1; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_xcpt; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_cause; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_tval; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_evec; // @[BackEnd.scala 81:19:@5588.4]
  wire  csr_io_illegal; // @[BackEnd.scala 81:19:@5588.4]
  wire [1:0] csr_io_retire; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_pc; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] csr_io_time; // @[BackEnd.scala 81:19:@5588.4]
  wire [31:0] InstDecoder_io_inst; // @[BackEnd.scala 86:25:@5594.4]
  wire [3:0] InstDecoder_io_cinfo_br_type; // @[BackEnd.scala 86:25:@5594.4]
  wire [1:0] InstDecoder_io_cinfo_op1_sel; // @[BackEnd.scala 86:25:@5594.4]
  wire [2:0] InstDecoder_io_cinfo_op2_sel; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 86:25:@5594.4]
  wire [3:0] InstDecoder_io_cinfo_alu_fun; // @[BackEnd.scala 86:25:@5594.4]
  wire [1:0] InstDecoder_io_cinfo_wb_sel; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_mem_en; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_mem_fcn; // @[BackEnd.scala 86:25:@5594.4]
  wire [2:0] InstDecoder_io_cinfo_mem_typ; // @[BackEnd.scala 86:25:@5594.4]
  wire [2:0] InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_illegal; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_is_branch; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_jal; // @[BackEnd.scala 86:25:@5594.4]
  wire  InstDecoder_io_cinfo_ret; // @[BackEnd.scala 86:25:@5594.4]
  wire [4:0] InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 86:25:@5594.4]
  wire [4:0] InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 86:25:@5594.4]
  wire [4:0] InstDecoder_io_cinfo_wbaddr; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_i; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_s; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_sb; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_u; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_uj; // @[BackEnd.scala 86:25:@5594.4]
  wire [31:0] InstDecoder_io_dinfo_imm_z; // @[BackEnd.scala 86:25:@5594.4]
  wire  regfile_clock; // @[BackEnd.scala 115:23:@5621.4]
  wire [4:0] regfile_io_rs1_addr; // @[BackEnd.scala 115:23:@5621.4]
  wire [31:0] regfile_io_rs1_data; // @[BackEnd.scala 115:23:@5621.4]
  wire [4:0] regfile_io_rs2_addr; // @[BackEnd.scala 115:23:@5621.4]
  wire [31:0] regfile_io_rs2_data; // @[BackEnd.scala 115:23:@5621.4]
  wire [4:0] regfile_io_waddr; // @[BackEnd.scala 115:23:@5621.4]
  wire [31:0] regfile_io_wdata; // @[BackEnd.scala 115:23:@5621.4]
  wire  regfile_io_wen; // @[BackEnd.scala 115:23:@5621.4]
  wire [31:0] ALU_io_op1; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_op2; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_pc; // @[BackEnd.scala 184:19:@5729.4]
  wire [3:0] ALU_io_ctrl_fun; // @[BackEnd.scala 184:19:@5729.4]
  wire [3:0] ALU_io_ctrl_br_type; // @[BackEnd.scala 184:19:@5729.4]
  wire [1:0] ALU_io_ctrl_wb_sel; // @[BackEnd.scala 184:19:@5729.4]
  wire [1:0] ALU_io_ctrl_pc_sel; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_rs2_data; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_result; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_target_brjmp; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_target_jpreg; // @[BackEnd.scala 184:19:@5729.4]
  wire [31:0] ALU_io_target_conti; // @[BackEnd.scala 184:19:@5729.4]
  reg  exe_rf_wen; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_0;
  reg [4:0] exe_wbaddr; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_1;
  reg  exe_mem_en; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_2;
  reg [2:0] exe_csr_cmd; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_3;
  reg  exe_illegal; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_4;
  reg [31:0] exe_pc; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_5;
  reg [31:0] exe_inst; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_6;
  reg [31:0] exe_rs2_data; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_7;
  reg [1:0] exe_wb_sel; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_8;
  reg  exe_mem_fcn; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_9;
  reg [2:0] exe_mem_typ; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_10;
  reg [3:0] exe_br_type; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_11;
  reg  exe_branch; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_12;
  reg  exe_jal; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_13;
  reg  exe_ret; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_14;
  reg [9:0] exe_pred_history; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_15;
  reg  exe_pred_diff; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_16;
  reg [31:0] exe_pred_tgt; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_17;
  reg [31:0] exe_op1_data; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_18;
  reg [31:0] exe_op2_data; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_19;
  reg [3:0] exe_alu_fun; // @[BackEnd.scala 89:22:@5599.4]
  reg [31:0] _RAND_20;
  reg  exe_valid; // @[BackEnd.scala 90:26:@5600.4]
  reg [31:0] _RAND_21;
  reg  mem_rf_wen; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_22;
  reg [4:0] mem_wbaddr; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_23;
  reg  mem_mem_en; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_24;
  reg [2:0] mem_csr_cmd; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_25;
  reg  mem_illegal; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_26;
  reg [31:0] mem_pc; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_27;
  reg [31:0] mem_inst; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_28;
  reg [1:0] mem_wb_sel; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_29;
  reg  mem_mem_fcn; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_30;
  reg [2:0] mem_mem_typ; // @[BackEnd.scala 92:22:@5602.4]
  reg [31:0] _RAND_31;
  reg  mem_valid; // @[BackEnd.scala 93:26:@5603.4]
  reg [31:0] _RAND_32;
  reg  wb_rf_wen; // @[BackEnd.scala 95:22:@5605.4]
  reg [31:0] _RAND_33;
  reg [4:0] wb_wbaddr; // @[BackEnd.scala 95:22:@5605.4]
  reg [31:0] _RAND_34;
  reg  wb_valid; // @[BackEnd.scala 96:26:@5606.4]
  reg [31:0] _RAND_35;
  reg [31:0] wb_wbdata; // @[BackEnd.scala 101:23:@5610.4]
  reg [31:0] _RAND_36;
  wire  dec_wire_rs1_oen; // @[BackEnd.scala 105:33:@5613.4]
  wire  dec_wire_rs2_oen; // @[BackEnd.scala 106:33:@5615.4]
  wire  _T_159; // @[BackEnd.scala 124:18:@5630.4]
  wire  _T_214; // @[BackEnd.scala 175:34:@5711.4]
  wire  _T_216; // @[BackEnd.scala 175:61:@5712.4]
  wire  exe_wire_rf_wen; // @[BackEnd.scala 175:47:@5713.4]
  wire  _T_160; // @[BackEnd.scala 124:42:@5631.4]
  wire  _T_161; // @[BackEnd.scala 125:18:@5632.4]
  wire  _T_286; // @[BackEnd.scala 241:34:@5829.4]
  wire  _T_288; // @[BackEnd.scala 241:61:@5830.4]
  wire  mem_wire_rf_wen; // @[BackEnd.scala 241:47:@5831.4]
  wire  _T_162; // @[BackEnd.scala 125:42:@5633.4]
  wire  _T_163; // @[BackEnd.scala 126:18:@5634.4]
  wire  _T_339; // @[BackEnd.scala 300:33:@5990.4]
  wire  _T_341; // @[BackEnd.scala 300:58:@5991.4]
  wire  wb_wire_rf_wen; // @[BackEnd.scala 300:45:@5992.4]
  wire  _T_164; // @[BackEnd.scala 126:42:@5635.4]
  wire [31:0] rf_rs1_data; // @[BackEnd.scala 116:25:@5624.4 BackEnd.scala 120:15:@5628.4]
  wire [31:0] _T_165; // @[Mux.scala 61:16:@5636.4]
  wire  _T_333; // @[BackEnd.scala 287:17:@5975.4]
  wire  _T_334; // @[BackEnd.scala 288:17:@5976.4]
  reg [31:0] mem_reg_exe_out; // @[BackEnd.scala 217:28:@5794.4]
  reg [31:0] _RAND_37;
  wire [31:0] _T_335; // @[Mux.scala 61:16:@5977.4]
  wire [31:0] mem_wbdata; // @[Mux.scala 61:16:@5978.4]
  wire [31:0] _T_166; // @[Mux.scala 61:16:@5637.4]
  wire [31:0] exe_wbdata; // @[BackEnd.scala 99:24:@5608.4 BackEnd.scala 192:14:@5739.4]
  wire [31:0] dec_rs1_data; // @[Mux.scala 61:16:@5638.4]
  wire  _T_168; // @[BackEnd.scala 130:18:@5640.4]
  wire  _T_169; // @[BackEnd.scala 130:42:@5641.4]
  wire  _T_170; // @[BackEnd.scala 131:18:@5642.4]
  wire  _T_171; // @[BackEnd.scala 131:42:@5643.4]
  wire  _T_172; // @[BackEnd.scala 132:18:@5644.4]
  wire  _T_173; // @[BackEnd.scala 132:42:@5645.4]
  wire [31:0] rf_rs2_data; // @[BackEnd.scala 117:25:@5625.4 BackEnd.scala 121:15:@5629.4]
  wire [31:0] _T_174; // @[Mux.scala 61:16:@5646.4]
  wire [31:0] _T_175; // @[Mux.scala 61:16:@5647.4]
  wire [31:0] dec_rs2_data; // @[Mux.scala 61:16:@5648.4]
  wire  _T_177; // @[BackEnd.scala 136:24:@5650.4]
  wire  _T_178; // @[BackEnd.scala 137:24:@5651.4]
  wire [31:0] _T_179; // @[Mux.scala 61:16:@5652.4]
  wire [31:0] dec_op1_data; // @[Mux.scala 61:16:@5653.4]
  wire  _T_181; // @[BackEnd.scala 140:24:@5655.4]
  wire  _T_182; // @[BackEnd.scala 141:24:@5656.4]
  wire  _T_183; // @[BackEnd.scala 142:24:@5657.4]
  wire  _T_184; // @[BackEnd.scala 143:24:@5658.4]
  wire  _T_185; // @[BackEnd.scala 144:24:@5659.4]
  wire [31:0] _T_186; // @[Mux.scala 61:16:@5660.4]
  wire [31:0] _T_187; // @[Mux.scala 61:16:@5661.4]
  wire [31:0] _T_188; // @[Mux.scala 61:16:@5662.4]
  wire [31:0] _T_189; // @[Mux.scala 61:16:@5663.4]
  wire [31:0] dec_op2_data; // @[Mux.scala 61:16:@5664.4]
  wire  exe_wire_mem_en; // @[BackEnd.scala 176:34:@5715.4]
  wire  _T_403; // @[BackEnd.scala 310:60:@6058.4]
  wire  exe_load_inst; // @[BackEnd.scala 310:45:@6059.4]
  wire  _T_405; // @[BackEnd.scala 313:20:@6061.4]
  wire  _T_407; // @[BackEnd.scala 313:79:@6062.4]
  wire  _T_408; // @[BackEnd.scala 313:57:@6063.4]
  wire  _T_409; // @[BackEnd.scala 313:87:@6064.4]
  wire  _T_411; // @[BackEnd.scala 314:20:@6066.4]
  wire  _T_413; // @[BackEnd.scala 314:79:@6067.4]
  wire  _T_414; // @[BackEnd.scala 314:57:@6068.4]
  wire  _T_415; // @[BackEnd.scala 314:87:@6069.4]
  wire  _T_416; // @[BackEnd.scala 313:108:@6070.4]
  wire [2:0] exe_wire_csr_cmd; // @[BackEnd.scala 177:26:@5717.4]
  wire  _T_417; // @[BackEnd.scala 315:22:@6071.4]
  wire  stall_0; // @[BackEnd.scala 314:108:@6072.4]
  wire  mem_wire_mem_en; // @[BackEnd.scala 242:34:@5833.4]
  wire  _T_423; // @[BackEnd.scala 318:42:@6077.4]
  wire  stall_2; // @[BackEnd.scala 318:39:@6078.4]
  wire  _T_195; // @[BackEnd.scala 146:51:@5668.4]
  wire  _T_196; // @[BackEnd.scala 146:48:@5669.4]
  wire  _T_197; // @[BackEnd.scala 146:70:@5670.4]
  wire  _T_205; // @[BackEnd.scala 150:34:@5679.8]
  wire  _T_206; // @[BackEnd.scala 150:31:@5680.8]
  wire  _T_207; // @[BackEnd.scala 154:44:@5684.8]
  wire  _T_208; // @[BackEnd.scala 154:75:@5685.8]
  wire  _T_209; // @[BackEnd.scala 154:54:@5686.8]
  wire  _T_211; // @[BackEnd.scala 155:26:@5687.8]
  wire  _T_212; // @[BackEnd.scala 154:86:@5688.8]
  wire [2:0] _T_213; // @[BackEnd.scala 154:24:@5689.8]
  wire  _GEN_0; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_1; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_2; // @[BackEnd.scala 149:54:@5678.6]
  wire [2:0] _GEN_3; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_4; // @[BackEnd.scala 149:54:@5678.6]
  wire [3:0] _GEN_5; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_6; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_7; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_8; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_9; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_10; // @[BackEnd.scala 149:54:@5678.6]
  wire [3:0] _GEN_11; // @[BackEnd.scala 149:54:@5678.6]
  wire [1:0] _GEN_12; // @[BackEnd.scala 149:54:@5678.6]
  wire [4:0] _GEN_13; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_14; // @[BackEnd.scala 149:54:@5678.6]
  wire [2:0] _GEN_15; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_16; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_17; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_18; // @[BackEnd.scala 149:54:@5678.6]
  wire [31:0] _GEN_19; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_20; // @[BackEnd.scala 149:54:@5678.6]
  wire [9:0] _GEN_21; // @[BackEnd.scala 149:54:@5678.6]
  wire  _GEN_23; // @[BackEnd.scala 146:94:@5671.4]
  wire [3:0] exe_wire_br_type; // @[BackEnd.scala 178:26:@5719.4]
  wire  exe_wire_branch; // @[BackEnd.scala 179:33:@5721.4]
  wire  exe_wire_jal; // @[BackEnd.scala 180:33:@5723.4]
  wire  exe_wire_ret; // @[BackEnd.scala 181:33:@5725.4]
  reg  _T_229; // @[BackEnd.scala 67:27:@5741.4]
  reg [31:0] _RAND_38;
  wire  _GEN_46; // @[BackEnd.scala 69:20:@5746.6]
  wire  _GEN_47; // @[BackEnd.scala 68:20:@5742.4]
  reg  _T_237; // @[BackEnd.scala 67:27:@5752.4]
  reg [31:0] _RAND_39;
  wire  _GEN_48; // @[BackEnd.scala 69:20:@5757.6]
  wire  _GEN_49; // @[BackEnd.scala 68:20:@5753.4]
  wire  _T_241; // @[BackEnd.scala 199:25:@5763.4]
  wire  _T_242; // @[BackEnd.scala 200:25:@5764.4]
  wire [31:0] _T_243; // @[BackEnd.scala 200:8:@5765.4]
  wire [31:0] next_pc; // @[BackEnd.scala 199:8:@5766.4]
  wire [1:0] _T_247; // @[BackEnd.scala 206:8:@5768.4]
  wire  _T_249; // @[BackEnd.scala 208:53:@5771.4]
  reg  _T_254; // @[BackEnd.scala 67:27:@5773.4]
  reg [31:0] _RAND_40;
  wire  _GEN_50; // @[BackEnd.scala 69:20:@5778.6]
  wire  _GEN_51; // @[BackEnd.scala 68:20:@5774.4]
  wire  _T_262; // @[BackEnd.scala 214:42:@5791.4]
  wire  mispredict; // @[BackEnd.scala 214:59:@5792.4]
  reg [31:0] mem_reg_jpnpc; // @[BackEnd.scala 218:28:@5795.4]
  reg [31:0] _RAND_41;
  wire  _T_269; // @[BackEnd.scala 219:47:@5798.4]
  wire [31:0] _T_277; // @[Bitwise.scala 72:12:@5820.8]
  wire [31:0] _T_278; // @[BackEnd.scala 236:70:@5821.8]
  wire [31:0] _T_283; // @[Bitwise.scala 72:12:@5824.8]
  wire [31:0] _T_284; // @[BackEnd.scala 237:70:@5825.8]
  wire [31:0] _T_285; // @[BackEnd.scala 236:90:@5826.8]
  wire  _GEN_52; // @[BackEnd.scala 221:34:@5804.6]
  wire  _GEN_53; // @[BackEnd.scala 221:34:@5804.6]
  wire  _GEN_54; // @[BackEnd.scala 221:34:@5804.6]
  wire [2:0] _GEN_55; // @[BackEnd.scala 221:34:@5804.6]
  wire  _GEN_56; // @[BackEnd.scala 221:34:@5804.6]
  wire [31:0] _GEN_57; // @[BackEnd.scala 221:34:@5804.6]
  wire [31:0] _GEN_58; // @[BackEnd.scala 221:34:@5804.6]
  wire [1:0] _GEN_59; // @[BackEnd.scala 221:34:@5804.6]
  wire [4:0] _GEN_60; // @[BackEnd.scala 221:34:@5804.6]
  wire  _GEN_62; // @[BackEnd.scala 221:34:@5804.6]
  wire [2:0] _GEN_63; // @[BackEnd.scala 221:34:@5804.6]
  wire [31:0] _GEN_64; // @[BackEnd.scala 221:34:@5804.6]
  wire [31:0] _GEN_65; // @[BackEnd.scala 221:34:@5804.6]
  wire  _GEN_66; // @[BackEnd.scala 219:71:@5799.4]
  wire  mem_wire_illegal; // @[BackEnd.scala 244:35:@5837.4]
  wire [1:0] _T_294; // @[BackEnd.scala 252:47:@5933.4]
  wire  _T_297; // @[BackEnd.scala 253:27:@5934.4]
  wire [1:0] _T_299; // @[BackEnd.scala 254:27:@5935.4]
  wire  _T_301; // @[BackEnd.scala 254:33:@5936.4]
  wire  _T_302; // @[Mux.scala 46:19:@5937.4]
  wire  _T_303; // @[Mux.scala 46:16:@5938.4]
  wire  _T_304; // @[Mux.scala 46:19:@5939.4]
  wire  ls_addr_ma_valid; // @[Mux.scala 46:16:@5940.4]
  wire [1:0] _T_305; // @[BackEnd.scala 256:39:@5941.4]
  wire  _T_307; // @[BackEnd.scala 256:45:@5942.4]
  wire  ma_jump; // @[BackEnd.scala 256:49:@5943.4]
  wire  _T_308; // @[BackEnd.scala 257:57:@5944.4]
  wire  _T_309; // @[BackEnd.scala 257:42:@5945.4]
  wire  ma_load; // @[BackEnd.scala 257:67:@5946.4]
  wire  _T_311; // @[BackEnd.scala 258:42:@5948.4]
  wire  ma_store; // @[BackEnd.scala 258:67:@5949.4]
  wire  _T_312; // @[BackEnd.scala 259:27:@5950.4]
  wire  _T_313; // @[BackEnd.scala 259:39:@5951.4]
  wire [1:0] _T_320; // @[Mux.scala 61:16:@5954.4]
  wire [2:0] _T_321; // @[Mux.scala 61:16:@5955.4]
  wire [2:0] _T_322; // @[Mux.scala 61:16:@5956.4]
  wire [2:0] _T_323; // @[Mux.scala 61:16:@5957.4]
  wire [31:0] _T_325; // @[Mux.scala 61:16:@5959.4]
  wire [31:0] _T_326; // @[Mux.scala 61:16:@5960.4]
  wire [31:0] _T_327; // @[Mux.scala 61:16:@5961.4]
  wire  _T_329; // @[BackEnd.scala 272:34:@5964.4]
  wire  _T_330; // @[BackEnd.scala 272:45:@5965.4]
  wire  _T_331; // @[BackEnd.scala 272:57:@5966.4]
  wire  _GEN_80; // @[BackEnd.scala 290:50:@5981.4]
  reg  _T_429; // @[BackEnd.scala 67:27:@6081.4]
  reg [31:0] _RAND_42;
  wire  _GEN_84; // @[BackEnd.scala 69:20:@6086.6]
  wire  _GEN_85; // @[BackEnd.scala 68:20:@6082.4]
  wire [2:0] _T_434; // @[BackEnd.scala 321:31:@6092.4]
  wire  _T_436; // @[BackEnd.scala 321:38:@6093.4]
  wire [7:0] _T_442; // @[BackEnd.scala 330:10:@6096.4]
  wire [7:0] _T_443; // @[BackEnd.scala 329:10:@6097.4]
  wire  _T_451; // @[BackEnd.scala 333:27:@6100.4]
  wire  _T_454; // @[BackEnd.scala 334:27:@6101.4]
  wire [7:0] _T_457; // @[BackEnd.scala 334:10:@6102.4]
  wire [7:0] _T_458; // @[BackEnd.scala 333:10:@6103.4]
  wire [7:0] _T_459; // @[BackEnd.scala 332:10:@6104.4]
  wire [7:0] _T_460; // @[BackEnd.scala 331:10:@6105.4]
  wire [7:0] _T_463; // @[BackEnd.scala 335:10:@6106.4]
  wire  _T_465; // @[BackEnd.scala 336:34:@6107.4]
  wire  _T_466; // @[BackEnd.scala 336:31:@6108.4]
  wire [31:0] _T_467; // @[BackEnd.scala 336:10:@6109.4]
  wire  _T_470; // @[BackEnd.scala 324:9:@6111.4]
  wire  _T_474; // @[BackEnd.scala 353:24:@6123.6]
  CSRFile csr ( // @[BackEnd.scala 81:19:@5588.4]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_status_prv(csr_io_status_prv),
    .io_status_unimp5(csr_io_status_unimp5),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_unimp4(csr_io_status_unimp4),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_unimp3(csr_io_status_unimp3),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_unimp2(csr_io_status_unimp2),
    .io_status_mie(csr_io_status_mie),
    .io_status_unimp1(csr_io_status_unimp1),
    .io_xcpt(csr_io_xcpt),
    .io_cause(csr_io_cause),
    .io_tval(csr_io_tval),
    .io_evec(csr_io_evec),
    .io_illegal(csr_io_illegal),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    .io_time(csr_io_time)
  );
  InstDecoder InstDecoder ( // @[BackEnd.scala 86:25:@5594.4]
    .io_inst(InstDecoder_io_inst),
    .io_cinfo_br_type(InstDecoder_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_io_cinfo_illegal),
    .io_cinfo_is_branch(InstDecoder_io_cinfo_is_branch),
    .io_cinfo_jal(InstDecoder_io_cinfo_jal),
    .io_cinfo_ret(InstDecoder_io_cinfo_ret),
    .io_cinfo_rs1_addr(InstDecoder_io_cinfo_rs1_addr),
    .io_cinfo_rs2_addr(InstDecoder_io_cinfo_rs2_addr),
    .io_cinfo_wbaddr(InstDecoder_io_cinfo_wbaddr),
    .io_dinfo_imm_i(InstDecoder_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_io_dinfo_imm_z)
  );
  Regfile regfile ( // @[BackEnd.scala 115:23:@5621.4]
    .clock(regfile_clock),
    .io_rs1_addr(regfile_io_rs1_addr),
    .io_rs1_data(regfile_io_rs1_data),
    .io_rs2_addr(regfile_io_rs2_addr),
    .io_rs2_data(regfile_io_rs2_data),
    .io_waddr(regfile_io_waddr),
    .io_wdata(regfile_io_wdata),
    .io_wen(regfile_io_wen)
  );
  ALU ALU ( // @[BackEnd.scala 184:19:@5729.4]
    .io_op1(ALU_io_op1),
    .io_op2(ALU_io_op2),
    .io_pc(ALU_io_pc),
    .io_ctrl_fun(ALU_io_ctrl_fun),
    .io_ctrl_br_type(ALU_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_io_ctrl_pc_sel),
    .io_rs2_data(ALU_io_rs2_data),
    .io_result(ALU_io_result),
    .io_target_brjmp(ALU_io_target_brjmp),
    .io_target_jpreg(ALU_io_target_jpreg),
    .io_target_conti(ALU_io_target_conti)
  );
  assign dec_wire_rs1_oen = io_front_inst_valid & InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 105:33:@5613.4]
  assign dec_wire_rs2_oen = io_front_inst_valid & InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 106:33:@5615.4]
  assign _T_159 = exe_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 124:18:@5630.4]
  assign _T_214 = exe_rf_wen & exe_valid; // @[BackEnd.scala 175:34:@5711.4]
  assign _T_216 = exe_wbaddr != 5'h0; // @[BackEnd.scala 175:61:@5712.4]
  assign exe_wire_rf_wen = _T_214 & _T_216; // @[BackEnd.scala 175:47:@5713.4]
  assign _T_160 = _T_159 & exe_wire_rf_wen; // @[BackEnd.scala 124:42:@5631.4]
  assign _T_161 = mem_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 125:18:@5632.4]
  assign _T_286 = mem_rf_wen & mem_valid; // @[BackEnd.scala 241:34:@5829.4]
  assign _T_288 = mem_wbaddr != 5'h0; // @[BackEnd.scala 241:61:@5830.4]
  assign mem_wire_rf_wen = _T_286 & _T_288; // @[BackEnd.scala 241:47:@5831.4]
  assign _T_162 = _T_161 & mem_wire_rf_wen; // @[BackEnd.scala 125:42:@5633.4]
  assign _T_163 = wb_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 126:18:@5634.4]
  assign _T_339 = wb_rf_wen & wb_valid; // @[BackEnd.scala 300:33:@5990.4]
  assign _T_341 = wb_wbaddr != 5'h0; // @[BackEnd.scala 300:58:@5991.4]
  assign wb_wire_rf_wen = _T_339 & _T_341; // @[BackEnd.scala 300:45:@5992.4]
  assign _T_164 = _T_163 & wb_wire_rf_wen; // @[BackEnd.scala 126:42:@5635.4]
  assign rf_rs1_data = regfile_io_rs1_data; // @[BackEnd.scala 116:25:@5624.4 BackEnd.scala 120:15:@5628.4]
  assign _T_165 = _T_164 ? wb_wbdata : rf_rs1_data; // @[Mux.scala 61:16:@5636.4]
  assign _T_333 = mem_wb_sel == 2'h1; // @[BackEnd.scala 287:17:@5975.4]
  assign _T_334 = mem_wb_sel == 2'h3; // @[BackEnd.scala 288:17:@5976.4]
  assign _T_335 = _T_334 ? csr_io_rw_rdata : mem_reg_exe_out; // @[Mux.scala 61:16:@5977.4]
  assign mem_wbdata = _T_333 ? io_mem_resp_bits_data : _T_335; // @[Mux.scala 61:16:@5978.4]
  assign _T_166 = _T_162 ? mem_wbdata : _T_165; // @[Mux.scala 61:16:@5637.4]
  assign exe_wbdata = ALU_io_result; // @[BackEnd.scala 99:24:@5608.4 BackEnd.scala 192:14:@5739.4]
  assign dec_rs1_data = _T_160 ? exe_wbdata : _T_166; // @[Mux.scala 61:16:@5638.4]
  assign _T_168 = exe_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 130:18:@5640.4]
  assign _T_169 = _T_168 & exe_wire_rf_wen; // @[BackEnd.scala 130:42:@5641.4]
  assign _T_170 = mem_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 131:18:@5642.4]
  assign _T_171 = _T_170 & mem_wire_rf_wen; // @[BackEnd.scala 131:42:@5643.4]
  assign _T_172 = wb_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 132:18:@5644.4]
  assign _T_173 = _T_172 & wb_wire_rf_wen; // @[BackEnd.scala 132:42:@5645.4]
  assign rf_rs2_data = regfile_io_rs2_data; // @[BackEnd.scala 117:25:@5625.4 BackEnd.scala 121:15:@5629.4]
  assign _T_174 = _T_173 ? wb_wbdata : rf_rs2_data; // @[Mux.scala 61:16:@5646.4]
  assign _T_175 = _T_171 ? mem_wbdata : _T_174; // @[Mux.scala 61:16:@5647.4]
  assign dec_rs2_data = _T_169 ? exe_wbdata : _T_175; // @[Mux.scala 61:16:@5648.4]
  assign _T_177 = InstDecoder_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 136:24:@5650.4]
  assign _T_178 = InstDecoder_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 137:24:@5651.4]
  assign _T_179 = _T_178 ? io_front_pc : dec_rs1_data; // @[Mux.scala 61:16:@5652.4]
  assign dec_op1_data = _T_177 ? InstDecoder_io_dinfo_imm_z : _T_179; // @[Mux.scala 61:16:@5653.4]
  assign _T_181 = InstDecoder_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 140:24:@5655.4]
  assign _T_182 = InstDecoder_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 141:24:@5656.4]
  assign _T_183 = InstDecoder_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 142:24:@5657.4]
  assign _T_184 = InstDecoder_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 143:24:@5658.4]
  assign _T_185 = InstDecoder_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 144:24:@5659.4]
  assign _T_186 = _T_185 ? InstDecoder_io_dinfo_imm_uj : dec_rs2_data; // @[Mux.scala 61:16:@5660.4]
  assign _T_187 = _T_184 ? InstDecoder_io_dinfo_imm_u : _T_186; // @[Mux.scala 61:16:@5661.4]
  assign _T_188 = _T_183 ? InstDecoder_io_dinfo_imm_sb : _T_187; // @[Mux.scala 61:16:@5662.4]
  assign _T_189 = _T_182 ? InstDecoder_io_dinfo_imm_s : _T_188; // @[Mux.scala 61:16:@5663.4]
  assign dec_op2_data = _T_181 ? InstDecoder_io_dinfo_imm_i : _T_189; // @[Mux.scala 61:16:@5664.4]
  assign exe_wire_mem_en = exe_mem_en & exe_valid; // @[BackEnd.scala 176:34:@5715.4]
  assign _T_403 = exe_mem_fcn == 1'h0; // @[BackEnd.scala 310:60:@6058.4]
  assign exe_load_inst = exe_wire_mem_en & _T_403; // @[BackEnd.scala 310:45:@6059.4]
  assign _T_405 = exe_load_inst & _T_159; // @[BackEnd.scala 313:20:@6061.4]
  assign _T_407 = InstDecoder_io_cinfo_rs1_addr != 5'h0; // @[BackEnd.scala 313:79:@6062.4]
  assign _T_408 = _T_405 & _T_407; // @[BackEnd.scala 313:57:@6063.4]
  assign _T_409 = _T_408 & dec_wire_rs1_oen; // @[BackEnd.scala 313:87:@6064.4]
  assign _T_411 = exe_load_inst & _T_168; // @[BackEnd.scala 314:20:@6066.4]
  assign _T_413 = InstDecoder_io_cinfo_rs2_addr != 5'h0; // @[BackEnd.scala 314:79:@6067.4]
  assign _T_414 = _T_411 & _T_413; // @[BackEnd.scala 314:57:@6068.4]
  assign _T_415 = _T_414 & dec_wire_rs2_oen; // @[BackEnd.scala 314:87:@6069.4]
  assign _T_416 = _T_409 | _T_415; // @[BackEnd.scala 313:108:@6070.4]
  assign exe_wire_csr_cmd = exe_valid ? exe_csr_cmd : 3'h0; // @[BackEnd.scala 177:26:@5717.4]
  assign _T_417 = exe_wire_csr_cmd != 3'h0; // @[BackEnd.scala 315:22:@6071.4]
  assign stall_0 = _T_416 | _T_417; // @[BackEnd.scala 314:108:@6072.4]
  assign mem_wire_mem_en = mem_mem_en & mem_valid; // @[BackEnd.scala 242:34:@5833.4]
  assign _T_423 = io_mem_resp_valid == 1'h0; // @[BackEnd.scala 318:42:@6077.4]
  assign stall_2 = mem_wire_mem_en & _T_423; // @[BackEnd.scala 318:39:@6078.4]
  assign _T_195 = stall_2 == 1'h0; // @[BackEnd.scala 146:51:@5668.4]
  assign _T_196 = stall_0 & _T_195; // @[BackEnd.scala 146:48:@5669.4]
  assign _T_197 = _T_196 | io_front_xcpt_valid; // @[BackEnd.scala 146:70:@5670.4]
  assign _T_205 = io_front_kill == 1'h0; // @[BackEnd.scala 150:34:@5679.8]
  assign _T_206 = io_front_inst_valid & _T_205; // @[BackEnd.scala 150:31:@5680.8]
  assign _T_207 = InstDecoder_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 154:44:@5684.8]
  assign _T_208 = InstDecoder_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 154:75:@5685.8]
  assign _T_209 = _T_207 | _T_208; // @[BackEnd.scala 154:54:@5686.8]
  assign _T_211 = InstDecoder_io_cinfo_rs1_addr == 5'h0; // @[BackEnd.scala 155:26:@5687.8]
  assign _T_212 = _T_209 & _T_211; // @[BackEnd.scala 154:86:@5688.8]
  assign _T_213 = _T_212 ? 3'h5 : InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 154:24:@5689.8]
  assign _GEN_0 = _T_195 ? _T_206 : exe_valid; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_1 = _T_195 ? InstDecoder_io_cinfo_rf_wen : exe_rf_wen; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_2 = _T_195 ? InstDecoder_io_cinfo_mem_en : exe_mem_en; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_3 = _T_195 ? _T_213 : exe_csr_cmd; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_4 = _T_195 ? InstDecoder_io_cinfo_illegal : exe_illegal; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_5 = _T_195 ? InstDecoder_io_cinfo_br_type : exe_br_type; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_6 = _T_195 ? io_front_pc : exe_pc; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_7 = _T_195 ? dec_op1_data : exe_op1_data; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_8 = _T_195 ? dec_op2_data : exe_op2_data; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_9 = _T_195 ? dec_rs2_data : exe_rs2_data; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_10 = _T_195 ? InstDecoder_io_inst : exe_inst; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_11 = _T_195 ? InstDecoder_io_cinfo_alu_fun : exe_alu_fun; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_12 = _T_195 ? InstDecoder_io_cinfo_wb_sel : exe_wb_sel; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_13 = _T_195 ? InstDecoder_io_cinfo_wbaddr : exe_wbaddr; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_14 = _T_195 ? InstDecoder_io_cinfo_mem_fcn : exe_mem_fcn; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_15 = _T_195 ? InstDecoder_io_cinfo_mem_typ : exe_mem_typ; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_16 = _T_195 ? InstDecoder_io_cinfo_is_branch : exe_branch; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_17 = _T_195 ? InstDecoder_io_cinfo_jal : exe_jal; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_18 = _T_195 ? InstDecoder_io_cinfo_ret : exe_ret; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_19 = _T_195 ? io_front_pred_tgt : exe_pred_tgt; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_20 = _T_195 ? io_front_pred_diff : exe_pred_diff; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_21 = _T_195 ? io_front_pred_history : exe_pred_history; // @[BackEnd.scala 149:54:@5678.6]
  assign _GEN_23 = _T_197 ? 1'h0 : _GEN_0; // @[BackEnd.scala 146:94:@5671.4]
  assign exe_wire_br_type = exe_valid ? exe_br_type : 4'h0; // @[BackEnd.scala 178:26:@5719.4]
  assign exe_wire_branch = exe_valid & exe_branch; // @[BackEnd.scala 179:33:@5721.4]
  assign exe_wire_jal = exe_valid & exe_jal; // @[BackEnd.scala 180:33:@5723.4]
  assign exe_wire_ret = exe_valid & exe_ret; // @[BackEnd.scala 181:33:@5725.4]
  assign _GEN_46 = exe_wire_ret ? 1'h0 : _T_229; // @[BackEnd.scala 69:20:@5746.6]
  assign _GEN_47 = _T_195 ? 1'h1 : _GEN_46; // @[BackEnd.scala 68:20:@5742.4]
  assign _GEN_48 = exe_wire_jal ? 1'h0 : _T_237; // @[BackEnd.scala 69:20:@5757.6]
  assign _GEN_49 = _T_195 ? 1'h1 : _GEN_48; // @[BackEnd.scala 68:20:@5753.4]
  assign _T_241 = ALU_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 199:25:@5763.4]
  assign _T_242 = ALU_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 200:25:@5764.4]
  assign _T_243 = _T_242 ? ALU_io_target_jpreg : ALU_io_target_conti; // @[BackEnd.scala 200:8:@5765.4]
  assign next_pc = _T_241 ? ALU_io_target_brjmp : _T_243; // @[BackEnd.scala 199:8:@5766.4]
  assign _T_247 = exe_wire_ret ? 2'h1 : 2'h3; // @[BackEnd.scala 206:8:@5768.4]
  assign _T_249 = exe_wire_br_type != 4'h0; // @[BackEnd.scala 208:53:@5771.4]
  assign _GEN_50 = _T_249 ? 1'h0 : _T_254; // @[BackEnd.scala 69:20:@5778.6]
  assign _GEN_51 = _T_195 ? 1'h1 : _GEN_50; // @[BackEnd.scala 68:20:@5774.4]
  assign _T_262 = next_pc != exe_pred_tgt; // @[BackEnd.scala 214:42:@5791.4]
  assign mispredict = _T_262 & exe_valid; // @[BackEnd.scala 214:59:@5792.4]
  assign _T_269 = stall_2 | io_front_xcpt_valid; // @[BackEnd.scala 219:47:@5798.4]
  assign _T_277 = _T_241 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@5820.8]
  assign _T_278 = _T_277 & ALU_io_target_brjmp; // @[BackEnd.scala 236:70:@5821.8]
  assign _T_283 = _T_242 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@5824.8]
  assign _T_284 = _T_283 & ALU_io_target_jpreg; // @[BackEnd.scala 237:70:@5825.8]
  assign _T_285 = _T_278 | _T_284; // @[BackEnd.scala 236:90:@5826.8]
  assign _GEN_52 = _T_195 ? exe_valid : mem_valid; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_53 = _T_195 ? exe_rf_wen : mem_rf_wen; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_54 = _T_195 ? exe_mem_en : mem_mem_en; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_55 = _T_195 ? exe_csr_cmd : mem_csr_cmd; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_56 = _T_195 ? exe_illegal : mem_illegal; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_57 = _T_195 ? exe_pc : mem_pc; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_58 = _T_195 ? exe_inst : mem_inst; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_59 = _T_195 ? exe_wb_sel : mem_wb_sel; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_60 = _T_195 ? exe_wbaddr : mem_wbaddr; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_62 = _T_195 ? exe_mem_fcn : mem_mem_fcn; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_63 = _T_195 ? exe_mem_typ : mem_mem_typ; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_64 = _T_195 ? exe_wbdata : mem_reg_exe_out; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_65 = _T_195 ? _T_285 : mem_reg_jpnpc; // @[BackEnd.scala 221:34:@5804.6]
  assign _GEN_66 = _T_269 ? 1'h0 : _GEN_52; // @[BackEnd.scala 219:71:@5799.4]
  assign mem_wire_illegal = mem_illegal & mem_valid; // @[BackEnd.scala 244:35:@5837.4]
  assign _T_294 = mem_mem_typ[1:0]; // @[BackEnd.scala 252:47:@5933.4]
  assign _T_297 = mem_reg_exe_out[0]; // @[BackEnd.scala 253:27:@5934.4]
  assign _T_299 = mem_reg_exe_out[1:0]; // @[BackEnd.scala 254:27:@5935.4]
  assign _T_301 = _T_299 != 2'h0; // @[BackEnd.scala 254:33:@5936.4]
  assign _T_302 = 2'h3 == _T_294; // @[Mux.scala 46:19:@5937.4]
  assign _T_303 = _T_302 ? _T_301 : 1'h0; // @[Mux.scala 46:16:@5938.4]
  assign _T_304 = 2'h2 == _T_294; // @[Mux.scala 46:19:@5939.4]
  assign ls_addr_ma_valid = _T_304 ? _T_297 : _T_303; // @[Mux.scala 46:16:@5940.4]
  assign _T_305 = mem_reg_jpnpc[1:0]; // @[BackEnd.scala 256:39:@5941.4]
  assign _T_307 = _T_305 != 2'h0; // @[BackEnd.scala 256:45:@5942.4]
  assign ma_jump = _T_307 & mem_valid; // @[BackEnd.scala 256:49:@5943.4]
  assign _T_308 = mem_mem_fcn == 1'h0; // @[BackEnd.scala 257:57:@5944.4]
  assign _T_309 = mem_wire_mem_en & _T_308; // @[BackEnd.scala 257:42:@5945.4]
  assign ma_load = _T_309 & ls_addr_ma_valid; // @[BackEnd.scala 257:67:@5946.4]
  assign _T_311 = mem_wire_mem_en & mem_mem_fcn; // @[BackEnd.scala 258:42:@5948.4]
  assign ma_store = _T_311 & ls_addr_ma_valid; // @[BackEnd.scala 258:67:@5949.4]
  assign _T_312 = ma_load | ma_store; // @[BackEnd.scala 259:27:@5950.4]
  assign _T_313 = _T_312 | ma_jump; // @[BackEnd.scala 259:39:@5951.4]
  assign _T_320 = mem_wire_illegal ? 2'h2 : 2'h0; // @[Mux.scala 61:16:@5954.4]
  assign _T_321 = ma_store ? 3'h6 : {{1'd0}, _T_320}; // @[Mux.scala 61:16:@5955.4]
  assign _T_322 = ma_load ? 3'h4 : _T_321; // @[Mux.scala 61:16:@5956.4]
  assign _T_323 = ma_jump ? 3'h0 : _T_322; // @[Mux.scala 61:16:@5957.4]
  assign _T_325 = mem_wire_illegal ? mem_inst : 32'h0; // @[Mux.scala 61:16:@5959.4]
  assign _T_326 = ma_store ? mem_reg_exe_out : _T_325; // @[Mux.scala 61:16:@5960.4]
  assign _T_327 = ma_load ? mem_reg_exe_out : _T_326; // @[Mux.scala 61:16:@5961.4]
  assign _T_329 = ma_jump | ma_load; // @[BackEnd.scala 272:34:@5964.4]
  assign _T_330 = _T_329 | ma_store; // @[BackEnd.scala 272:45:@5965.4]
  assign _T_331 = _T_330 | mem_wire_illegal; // @[BackEnd.scala 272:57:@5966.4]
  assign _GEN_80 = _T_269 ? 1'h0 : mem_valid; // @[BackEnd.scala 290:50:@5981.4]
  assign _GEN_84 = mispredict ? 1'h0 : _T_429; // @[BackEnd.scala 69:20:@6086.6]
  assign _GEN_85 = _T_195 ? 1'h1 : _GEN_84; // @[BackEnd.scala 68:20:@6082.4]
  assign _T_434 = {stall_2,1'h0,stall_0}; // @[BackEnd.scala 321:31:@6092.4]
  assign _T_436 = _T_434 != 3'h0; // @[BackEnd.scala 321:38:@6093.4]
  assign _T_442 = stall_0 ? 8'h53 : 8'h20; // @[BackEnd.scala 330:10:@6096.4]
  assign _T_443 = stall_2 ? 8'h46 : _T_442; // @[BackEnd.scala 329:10:@6097.4]
  assign _T_451 = ALU_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 333:27:@6100.4]
  assign _T_454 = ALU_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 334:27:@6101.4]
  assign _T_457 = _T_454 ? 8'h20 : 8'h3f; // @[BackEnd.scala 334:10:@6102.4]
  assign _T_458 = _T_451 ? 8'h45 : _T_457; // @[BackEnd.scala 333:10:@6103.4]
  assign _T_459 = _T_242 ? 8'h4a : _T_458; // @[BackEnd.scala 332:10:@6104.4]
  assign _T_460 = _T_241 ? 8'h42 : _T_459; // @[BackEnd.scala 331:10:@6105.4]
  assign _T_463 = csr_io_illegal ? 8'h58 : 8'h20; // @[BackEnd.scala 335:10:@6106.4]
  assign _T_465 = exe_valid == 1'h0; // @[BackEnd.scala 336:34:@6107.4]
  assign _T_466 = io_front_xcpt_valid | _T_465; // @[BackEnd.scala 336:31:@6108.4]
  assign _T_467 = _T_466 ? 32'h4033 : exe_inst; // @[BackEnd.scala 336:10:@6109.4]
  assign _T_470 = reset == 1'h0; // @[BackEnd.scala 324:9:@6111.4]
  assign _T_474 = ALU_io_target_conti != exe_pred_tgt; // @[BackEnd.scala 353:24:@6123.6]
  assign io_mem_req_valid = exe_mem_en & exe_valid; // @[BackEnd.scala 276:24:@5970.4]
  assign io_mem_req_bits_addr = ALU_io_result; // @[BackEnd.scala 277:24:@5971.4]
  assign io_mem_req_bits_data = exe_rs2_data; // @[BackEnd.scala 280:24:@5974.4]
  assign io_mem_req_bits_fcn = exe_mem_fcn; // @[BackEnd.scala 278:24:@5972.4]
  assign io_mem_req_bits_typ = exe_mem_typ; // @[BackEnd.scala 279:24:@5973.4]
  assign io_cyc = csr_io_time; // @[BackEnd.scala 82:10:@5592.4]
  assign io_front_xcpt_valid = _T_331 | csr_io_eret; // @[BackEnd.scala 272:23:@5968.4]
  assign io_front_xcpt_bits = csr_io_evec; // @[BackEnd.scala 273:23:@5969.4]
  assign io_front_kill = mispredict & _T_429; // @[BackEnd.scala 320:17:@6090.4]
  assign io_front_forward = _T_436 == 1'h0; // @[BackEnd.scala 321:21:@6095.4]
  assign io_front_ras_pop = exe_wire_ret & _T_229; // @[BackEnd.scala 194:27:@5750.4]
  assign io_front_ras_push_valid = exe_wire_jal & _T_237; // @[BackEnd.scala 195:27:@5761.4]
  assign io_front_ras_push_bits = ALU_io_target_conti; // @[BackEnd.scala 196:27:@5762.4]
  assign io_front_fb_pc = exe_pc; // @[BackEnd.scala 203:18:@5767.4]
  assign io_front_fb_type = exe_wire_branch ? 2'h2 : _T_247; // @[BackEnd.scala 204:20:@5770.4]
  assign io_front_feedBack_redirect = _T_241 | _T_242; // @[BackEnd.scala 210:30:@5787.4]
  assign io_front_feedBack_history = exe_pred_history; // @[BackEnd.scala 211:30:@5788.4]
  assign io_front_feedBack_diff = exe_pred_diff; // @[BackEnd.scala 212:30:@5789.4]
  assign io_front_feedBack_tgt = _T_241 ? ALU_io_target_brjmp : _T_243; // @[BackEnd.scala 209:25:@5783.4]
  assign io_front_feedBack_valid = _T_249 & _T_254; // @[BackEnd.scala 208:27:@5782.4]
  assign csr_clock = clock; // @[:@5589.4]
  assign csr_reset = reset; // @[:@5590.4]
  assign csr_io_rw_cmd = mem_valid ? mem_csr_cmd : 3'h0; // @[BackEnd.scala 249:19:@5931.4]
  assign csr_io_rw_addr = mem_inst[31:20]; // @[BackEnd.scala 247:19:@5929.4]
  assign csr_io_rw_wdata = mem_reg_exe_out; // @[BackEnd.scala 248:19:@5930.4]
  assign csr_io_xcpt = _T_313 | mem_wire_illegal; // @[BackEnd.scala 259:16:@5953.4]
  assign csr_io_cause = {{29'd0}, _T_323}; // @[BackEnd.scala 260:16:@5958.4]
  assign csr_io_tval = ma_jump ? mem_reg_jpnpc : _T_327; // @[BackEnd.scala 266:16:@5963.4]
  assign csr_io_illegal = 1'h0;
  assign csr_io_retire = {{1'd0}, wb_valid}; // @[BackEnd.scala 305:20:@5997.4]
  assign csr_io_pc = mem_pc; // @[BackEnd.scala 250:19:@5932.4]
  assign InstDecoder_io_inst = io_front_inst_bits; // @[BackEnd.scala 103:20:@5611.4]
  assign regfile_clock = clock; // @[:@5622.4]
  assign regfile_io_rs1_addr = InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 118:23:@5626.4]
  assign regfile_io_rs2_addr = InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 119:23:@5627.4]
  assign regfile_io_waddr = wb_wbaddr; // @[BackEnd.scala 301:20:@5994.4]
  assign regfile_io_wdata = wb_wbdata; // @[BackEnd.scala 302:20:@5995.4]
  assign regfile_io_wen = _T_339 & _T_341; // @[BackEnd.scala 303:20:@5996.4]
  assign ALU_io_op1 = exe_op1_data; // @[BackEnd.scala 185:20:@5732.4]
  assign ALU_io_op2 = exe_op2_data; // @[BackEnd.scala 186:20:@5733.4]
  assign ALU_io_pc = exe_pc; // @[BackEnd.scala 188:20:@5735.4]
  assign ALU_io_ctrl_fun = exe_alu_fun; // @[BackEnd.scala 189:20:@5736.4]
  assign ALU_io_ctrl_br_type = exe_valid ? exe_br_type : 4'h0; // @[BackEnd.scala 190:20:@5737.4]
  assign ALU_io_ctrl_wb_sel = exe_wb_sel; // @[BackEnd.scala 191:20:@5738.4]
  assign ALU_io_rs2_data = exe_rs2_data; // @[BackEnd.scala 187:20:@5734.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exe_rf_wen = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  exe_wbaddr = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  exe_mem_en = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  exe_csr_cmd = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  exe_illegal = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  exe_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  exe_inst = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  exe_rs2_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  exe_wb_sel = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  exe_mem_fcn = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  exe_mem_typ = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  exe_br_type = _RAND_11[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  exe_branch = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  exe_jal = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  exe_ret = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  exe_pred_history = _RAND_15[9:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  exe_pred_diff = _RAND_16[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  exe_pred_tgt = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  exe_op1_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  exe_op2_data = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  exe_alu_fun = _RAND_20[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  exe_valid = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_rf_wen = _RAND_22[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_wbaddr = _RAND_23[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_mem_en = _RAND_24[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_csr_cmd = _RAND_25[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_illegal = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_pc = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_inst = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_wb_sel = _RAND_29[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  mem_mem_fcn = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  mem_mem_typ = _RAND_31[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  mem_valid = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_rf_wen = _RAND_33[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  wb_wbaddr = _RAND_34[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  wb_valid = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  wb_wbdata = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_reg_exe_out = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_229 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_237 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  _T_254 = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  mem_reg_jpnpc = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  _T_429 = _RAND_42[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_rf_wen <= InstDecoder_io_cinfo_rf_wen;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_wbaddr <= InstDecoder_io_cinfo_wbaddr;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_mem_en <= InstDecoder_io_cinfo_mem_en;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        if (_T_212) begin
          exe_csr_cmd <= 3'h5;
        end else begin
          exe_csr_cmd <= InstDecoder_io_cinfo_csr_cmd;
        end
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_illegal <= InstDecoder_io_cinfo_illegal;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_pc <= io_front_pc;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_inst <= InstDecoder_io_inst;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        if (_T_169) begin
          exe_rs2_data <= exe_wbdata;
        end else begin
          if (_T_171) begin
            if (_T_333) begin
              exe_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_334) begin
                exe_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_rs2_data <= mem_reg_exe_out;
              end
            end
          end else begin
            if (_T_173) begin
              exe_rs2_data <= wb_wbdata;
            end else begin
              exe_rs2_data <= rf_rs2_data;
            end
          end
        end
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_wb_sel <= InstDecoder_io_cinfo_wb_sel;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_mem_fcn <= InstDecoder_io_cinfo_mem_fcn;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_mem_typ <= InstDecoder_io_cinfo_mem_typ;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_br_type <= InstDecoder_io_cinfo_br_type;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_branch <= InstDecoder_io_cinfo_is_branch;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_jal <= InstDecoder_io_cinfo_jal;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_ret <= InstDecoder_io_cinfo_ret;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_pred_history <= io_front_pred_history;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_pred_diff <= io_front_pred_diff;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_pred_tgt <= io_front_pred_tgt;
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        if (_T_177) begin
          exe_op1_data <= InstDecoder_io_dinfo_imm_z;
        end else begin
          if (_T_178) begin
            exe_op1_data <= io_front_pc;
          end else begin
            if (_T_160) begin
              exe_op1_data <= exe_wbdata;
            end else begin
              if (_T_162) begin
                if (_T_333) begin
                  exe_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_334) begin
                    exe_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_op1_data <= mem_reg_exe_out;
                  end
                end
              end else begin
                if (_T_164) begin
                  exe_op1_data <= wb_wbdata;
                end else begin
                  exe_op1_data <= rf_rs1_data;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        if (_T_181) begin
          exe_op2_data <= InstDecoder_io_dinfo_imm_i;
        end else begin
          if (_T_182) begin
            exe_op2_data <= InstDecoder_io_dinfo_imm_s;
          end else begin
            if (_T_183) begin
              exe_op2_data <= InstDecoder_io_dinfo_imm_sb;
            end else begin
              if (_T_184) begin
                exe_op2_data <= InstDecoder_io_dinfo_imm_u;
              end else begin
                if (_T_185) begin
                  exe_op2_data <= InstDecoder_io_dinfo_imm_uj;
                end else begin
                  if (_T_169) begin
                    exe_op2_data <= exe_wbdata;
                  end else begin
                    if (_T_171) begin
                      if (_T_333) begin
                        exe_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_334) begin
                          exe_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_op2_data <= mem_reg_exe_out;
                        end
                      end
                    end else begin
                      if (_T_173) begin
                        exe_op2_data <= wb_wbdata;
                      end else begin
                        exe_op2_data <= rf_rs2_data;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_197)) begin
      if (_T_195) begin
        exe_alu_fun <= InstDecoder_io_cinfo_alu_fun;
      end
    end
    if (reset) begin
      exe_valid <= 1'h0;
    end else begin
      if (_T_197) begin
        exe_valid <= 1'h0;
      end else begin
        if (_T_195) begin
          exe_valid <= _T_206;
        end
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_rf_wen <= exe_rf_wen;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_wbaddr <= exe_wbaddr;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_mem_en <= exe_mem_en;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_csr_cmd <= exe_csr_cmd;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_illegal <= exe_illegal;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_pc <= exe_pc;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_inst <= exe_inst;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_wb_sel <= exe_wb_sel;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_mem_fcn <= exe_mem_fcn;
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_mem_typ <= exe_mem_typ;
      end
    end
    if (reset) begin
      mem_valid <= 1'h0;
    end else begin
      if (_T_269) begin
        mem_valid <= 1'h0;
      end else begin
        if (_T_195) begin
          mem_valid <= exe_valid;
        end
      end
    end
    if (!(_T_269)) begin
      wb_rf_wen <= mem_rf_wen;
    end
    if (!(_T_269)) begin
      wb_wbaddr <= mem_wbaddr;
    end
    if (reset) begin
      wb_valid <= 1'h0;
    end else begin
      if (_T_269) begin
        wb_valid <= 1'h0;
      end else begin
        wb_valid <= mem_valid;
      end
    end
    if (!(_T_269)) begin
      if (_T_333) begin
        wb_wbdata <= io_mem_resp_bits_data;
      end else begin
        if (_T_334) begin
          wb_wbdata <= csr_io_rw_rdata;
        end else begin
          wb_wbdata <= mem_reg_exe_out;
        end
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_reg_exe_out <= exe_wbdata;
      end
    end
    if (reset) begin
      _T_229 <= 1'h1;
    end else begin
      if (_T_195) begin
        _T_229 <= 1'h1;
      end else begin
        if (exe_wire_ret) begin
          _T_229 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_237 <= 1'h1;
    end else begin
      if (_T_195) begin
        _T_237 <= 1'h1;
      end else begin
        if (exe_wire_jal) begin
          _T_237 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_254 <= 1'h1;
    end else begin
      if (_T_195) begin
        _T_254 <= 1'h1;
      end else begin
        if (_T_249) begin
          _T_254 <= 1'h0;
        end
      end
    end
    if (!(_T_269)) begin
      if (_T_195) begin
        mem_reg_jpnpc <= _T_285;
      end
    end
    if (reset) begin
      _T_429 <= 1'h1;
    end else begin
      if (_T_195) begin
        _T_429 <= 1'h1;
      end else begin
        if (mispredict) begin
          _T_429 <= 1'h0;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_470) begin
          $fwrite(32'h80000002,"Core: Cyc= %d (%x, %x, %x) %c %c %c ExeInst: DASM(%x)\n",io_cyc,io_front_pc,exe_pc,mem_pc,_T_443,_T_460,_T_463,_T_467); // @[BackEnd.scala 324:9:@6113.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid & _T_470) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_rf_wen,wb_wbaddr,wb_wbdata); // @[BackEnd.scala 339:11:@6119.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_front_feedBack_valid & _T_470) begin
          $fwrite(32'h80000002,"BranchJump: Cyc= %d kill %x pc %x tgt %x actual %x expect %x inst DASM(%x)\n",io_cyc,mispredict,exe_pc,next_pc,io_front_feedBack_redirect,_T_474,exe_inst); // @[BackEnd.scala 347:11:@6127.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module chiwen( // @[:@6131.2]
  input         clock, // @[:@6132.4]
  input         reset, // @[:@6133.4]
  input  [31:0] io_imem_r_data, // @[:@6134.4]
  input         io_imem_r_valid, // @[:@6134.4]
  input         io_imem_r_last, // @[:@6134.4]
  input         io_imem_ar_ready, // @[:@6134.4]
  output        io_imem_ar_valid, // @[:@6134.4]
  output [31:0] io_imem_ar_addr, // @[:@6134.4]
  output        io_dmem_req_valid, // @[:@6134.4]
  output [31:0] io_dmem_req_bits_addr, // @[:@6134.4]
  output [31:0] io_dmem_req_bits_data, // @[:@6134.4]
  output        io_dmem_req_bits_fcn, // @[:@6134.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:@6134.4]
  input         io_dmem_resp_valid, // @[:@6134.4]
  input  [31:0] io_dmem_resp_bits_data // @[:@6134.4]
);
  wire  frontEnd_clock; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_reset; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_cyc; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_mem_r_data; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_mem_r_valid; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_mem_r_last; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_mem_ar_ready; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_mem_ar_valid; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_mem_ar_addr; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_xcpt_valid; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_xcpt_bits; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_kill; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_forward; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_inst_valid; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_inst_bits; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_pc; // @[Core.scala 29:24:@6136.4]
  wire [9:0] frontEnd_io_back_pred_history; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_pred_diff; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_pred_tgt; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_ras_pop; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_ras_push_valid; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_ras_push_bits; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_fb_pc; // @[Core.scala 29:24:@6136.4]
  wire [1:0] frontEnd_io_back_fb_type; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_feedBack_redirect; // @[Core.scala 29:24:@6136.4]
  wire [9:0] frontEnd_io_back_feedBack_history; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_feedBack_diff; // @[Core.scala 29:24:@6136.4]
  wire [31:0] frontEnd_io_back_feedBack_tgt; // @[Core.scala 29:24:@6136.4]
  wire  frontEnd_io_back_feedBack_valid; // @[Core.scala 29:24:@6136.4]
  wire  backEnd_clock; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_reset; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_mem_req_valid; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_mem_req_bits_addr; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_mem_req_bits_data; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_mem_req_bits_fcn; // @[Core.scala 30:24:@6139.4]
  wire [2:0] backEnd_io_mem_req_bits_typ; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_mem_resp_valid; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_mem_resp_bits_data; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_cyc; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_xcpt_valid; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_xcpt_bits; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_kill; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_forward; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_inst_valid; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_inst_bits; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_pc; // @[Core.scala 30:24:@6139.4]
  wire [9:0] backEnd_io_front_pred_history; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_pred_diff; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_pred_tgt; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_ras_pop; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_ras_push_valid; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_ras_push_bits; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_fb_pc; // @[Core.scala 30:24:@6139.4]
  wire [1:0] backEnd_io_front_fb_type; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_feedBack_redirect; // @[Core.scala 30:24:@6139.4]
  wire [9:0] backEnd_io_front_feedBack_history; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_feedBack_diff; // @[Core.scala 30:24:@6139.4]
  wire [31:0] backEnd_io_front_feedBack_tgt; // @[Core.scala 30:24:@6139.4]
  wire  backEnd_io_front_feedBack_valid; // @[Core.scala 30:24:@6139.4]
  FrontEnd frontEnd ( // @[Core.scala 29:24:@6136.4]
    .clock(frontEnd_clock),
    .reset(frontEnd_reset),
    .io_cyc(frontEnd_io_cyc),
    .io_mem_r_data(frontEnd_io_mem_r_data),
    .io_mem_r_valid(frontEnd_io_mem_r_valid),
    .io_mem_r_last(frontEnd_io_mem_r_last),
    .io_mem_ar_ready(frontEnd_io_mem_ar_ready),
    .io_mem_ar_valid(frontEnd_io_mem_ar_valid),
    .io_mem_ar_addr(frontEnd_io_mem_ar_addr),
    .io_back_xcpt_valid(frontEnd_io_back_xcpt_valid),
    .io_back_xcpt_bits(frontEnd_io_back_xcpt_bits),
    .io_back_kill(frontEnd_io_back_kill),
    .io_back_forward(frontEnd_io_back_forward),
    .io_back_inst_valid(frontEnd_io_back_inst_valid),
    .io_back_inst_bits(frontEnd_io_back_inst_bits),
    .io_back_pc(frontEnd_io_back_pc),
    .io_back_pred_history(frontEnd_io_back_pred_history),
    .io_back_pred_diff(frontEnd_io_back_pred_diff),
    .io_back_pred_tgt(frontEnd_io_back_pred_tgt),
    .io_back_ras_pop(frontEnd_io_back_ras_pop),
    .io_back_ras_push_valid(frontEnd_io_back_ras_push_valid),
    .io_back_ras_push_bits(frontEnd_io_back_ras_push_bits),
    .io_back_fb_pc(frontEnd_io_back_fb_pc),
    .io_back_fb_type(frontEnd_io_back_fb_type),
    .io_back_feedBack_redirect(frontEnd_io_back_feedBack_redirect),
    .io_back_feedBack_history(frontEnd_io_back_feedBack_history),
    .io_back_feedBack_diff(frontEnd_io_back_feedBack_diff),
    .io_back_feedBack_tgt(frontEnd_io_back_feedBack_tgt),
    .io_back_feedBack_valid(frontEnd_io_back_feedBack_valid)
  );
  BackEnd backEnd ( // @[Core.scala 30:24:@6139.4]
    .clock(backEnd_clock),
    .reset(backEnd_reset),
    .io_mem_req_valid(backEnd_io_mem_req_valid),
    .io_mem_req_bits_addr(backEnd_io_mem_req_bits_addr),
    .io_mem_req_bits_data(backEnd_io_mem_req_bits_data),
    .io_mem_req_bits_fcn(backEnd_io_mem_req_bits_fcn),
    .io_mem_req_bits_typ(backEnd_io_mem_req_bits_typ),
    .io_mem_resp_valid(backEnd_io_mem_resp_valid),
    .io_mem_resp_bits_data(backEnd_io_mem_resp_bits_data),
    .io_cyc(backEnd_io_cyc),
    .io_front_xcpt_valid(backEnd_io_front_xcpt_valid),
    .io_front_xcpt_bits(backEnd_io_front_xcpt_bits),
    .io_front_kill(backEnd_io_front_kill),
    .io_front_forward(backEnd_io_front_forward),
    .io_front_inst_valid(backEnd_io_front_inst_valid),
    .io_front_inst_bits(backEnd_io_front_inst_bits),
    .io_front_pc(backEnd_io_front_pc),
    .io_front_pred_history(backEnd_io_front_pred_history),
    .io_front_pred_diff(backEnd_io_front_pred_diff),
    .io_front_pred_tgt(backEnd_io_front_pred_tgt),
    .io_front_ras_pop(backEnd_io_front_ras_pop),
    .io_front_ras_push_valid(backEnd_io_front_ras_push_valid),
    .io_front_ras_push_bits(backEnd_io_front_ras_push_bits),
    .io_front_fb_pc(backEnd_io_front_fb_pc),
    .io_front_fb_type(backEnd_io_front_fb_type),
    .io_front_feedBack_redirect(backEnd_io_front_feedBack_redirect),
    .io_front_feedBack_history(backEnd_io_front_feedBack_history),
    .io_front_feedBack_diff(backEnd_io_front_feedBack_diff),
    .io_front_feedBack_tgt(backEnd_io_front_feedBack_tgt),
    .io_front_feedBack_valid(backEnd_io_front_feedBack_valid)
  );
  assign io_imem_ar_valid = frontEnd_io_mem_ar_valid; // @[Core.scala 31:20:@6147.4]
  assign io_imem_ar_addr = frontEnd_io_mem_ar_addr; // @[Core.scala 31:20:@6145.4]
  assign io_dmem_req_valid = backEnd_io_mem_req_valid; // @[Core.scala 32:20:@6159.4]
  assign io_dmem_req_bits_addr = backEnd_io_mem_req_bits_addr; // @[Core.scala 32:20:@6158.4]
  assign io_dmem_req_bits_data = backEnd_io_mem_req_bits_data; // @[Core.scala 32:20:@6157.4]
  assign io_dmem_req_bits_fcn = backEnd_io_mem_req_bits_fcn; // @[Core.scala 32:20:@6156.4]
  assign io_dmem_req_bits_typ = backEnd_io_mem_req_bits_typ; // @[Core.scala 32:20:@6155.4]
  assign frontEnd_clock = clock; // @[:@6137.4]
  assign frontEnd_reset = reset; // @[:@6138.4]
  assign frontEnd_io_cyc = backEnd_io_cyc; // @[Core.scala 34:20:@6182.4]
  assign frontEnd_io_mem_r_data = io_imem_r_data; // @[Core.scala 31:20:@6152.4]
  assign frontEnd_io_mem_r_valid = io_imem_r_valid; // @[Core.scala 31:20:@6151.4]
  assign frontEnd_io_mem_r_last = io_imem_r_last; // @[Core.scala 31:20:@6150.4]
  assign frontEnd_io_mem_ar_ready = io_imem_ar_ready; // @[Core.scala 31:20:@6148.4]
  assign frontEnd_io_back_xcpt_valid = backEnd_io_front_xcpt_valid; // @[Core.scala 33:20:@6181.4]
  assign frontEnd_io_back_xcpt_bits = backEnd_io_front_xcpt_bits; // @[Core.scala 33:20:@6180.4]
  assign frontEnd_io_back_kill = backEnd_io_front_kill; // @[Core.scala 33:20:@6179.4]
  assign frontEnd_io_back_forward = backEnd_io_front_forward; // @[Core.scala 33:20:@6178.4]
  assign frontEnd_io_back_ras_pop = backEnd_io_front_ras_pop; // @[Core.scala 33:20:@6170.4]
  assign frontEnd_io_back_ras_push_valid = backEnd_io_front_ras_push_valid; // @[Core.scala 33:20:@6169.4]
  assign frontEnd_io_back_ras_push_bits = backEnd_io_front_ras_push_bits; // @[Core.scala 33:20:@6168.4]
  assign frontEnd_io_back_fb_pc = backEnd_io_front_fb_pc; // @[Core.scala 33:20:@6167.4]
  assign frontEnd_io_back_fb_type = backEnd_io_front_fb_type; // @[Core.scala 33:20:@6166.4]
  assign frontEnd_io_back_feedBack_redirect = backEnd_io_front_feedBack_redirect; // @[Core.scala 33:20:@6165.4]
  assign frontEnd_io_back_feedBack_history = backEnd_io_front_feedBack_history; // @[Core.scala 33:20:@6164.4]
  assign frontEnd_io_back_feedBack_diff = backEnd_io_front_feedBack_diff; // @[Core.scala 33:20:@6163.4]
  assign frontEnd_io_back_feedBack_tgt = backEnd_io_front_feedBack_tgt; // @[Core.scala 33:20:@6162.4]
  assign frontEnd_io_back_feedBack_valid = backEnd_io_front_feedBack_valid; // @[Core.scala 33:20:@6161.4]
  assign backEnd_clock = clock; // @[:@6140.4]
  assign backEnd_reset = reset; // @[:@6141.4]
  assign backEnd_io_mem_resp_valid = io_dmem_resp_valid; // @[Core.scala 32:20:@6154.4]
  assign backEnd_io_mem_resp_bits_data = io_dmem_resp_bits_data; // @[Core.scala 32:20:@6153.4]
  assign backEnd_io_front_inst_valid = frontEnd_io_back_inst_valid; // @[Core.scala 33:20:@6177.4]
  assign backEnd_io_front_inst_bits = frontEnd_io_back_inst_bits; // @[Core.scala 33:20:@6176.4]
  assign backEnd_io_front_pc = frontEnd_io_back_pc; // @[Core.scala 33:20:@6175.4]
  assign backEnd_io_front_pred_history = frontEnd_io_back_pred_history; // @[Core.scala 33:20:@6173.4]
  assign backEnd_io_front_pred_diff = frontEnd_io_back_pred_diff; // @[Core.scala 33:20:@6172.4]
  assign backEnd_io_front_pred_tgt = frontEnd_io_back_pred_tgt; // @[Core.scala 33:20:@6171.4]
endmodule
