module FetchInst( // @[:@709.2]
  input         clock, // @[:@710.4]
  input         reset, // @[:@711.4]
  input  [31:0] io_cyc, // @[:@712.4]
  input         io_mem_addr_ready, // @[:@712.4]
  output        io_mem_addr_valid, // @[:@712.4]
  output [31:0] io_mem_addr_bits, // @[:@712.4]
  input         io_mem_inst_0_valid, // @[:@712.4]
  input  [31:0] io_mem_inst_0_bits, // @[:@712.4]
  input         io_mem_inst_1_valid, // @[:@712.4]
  input  [31:0] io_mem_inst_1_bits, // @[:@712.4]
  input         io_if_kill, // @[:@712.4]
  input         io_if_fence, // @[:@712.4]
  input  [31:0] io_if_target, // @[:@712.4]
  input         io_if_split, // @[:@712.4]
  input  [31:0] io_btb_target, // @[:@712.4]
  input         io_dec_forward_0, // @[:@712.4]
  input         io_dec_forward_1, // @[:@712.4]
  input         io_dec_kill_0, // @[:@712.4]
  input         io_dec_kill_1, // @[:@712.4]
  output [31:0] io_if_pc, // @[:@712.4]
  output        io_if_forward_0, // @[:@712.4]
  output        io_if_forward_1, // @[:@712.4]
  output        io_dec_inst_0_valid, // @[:@712.4]
  output [31:0] io_dec_inst_0_bits, // @[:@712.4]
  output        io_dec_inst_1_valid, // @[:@712.4]
  output [31:0] io_dec_inst_1_bits // @[:@712.4]
);
  reg  pc_state; // @[FetchInst.scala 27:25:@714.4]
  reg [31:0] _RAND_0;
  reg [1:0] inst_state_0; // @[FetchInst.scala 29:27:@718.4]
  reg [31:0] _RAND_1;
  reg [1:0] inst_state_1; // @[FetchInst.scala 29:27:@718.4]
  reg [31:0] _RAND_2;
  reg [31:0] if_reg_pc; // @[FetchInst.scala 31:26:@719.4]
  reg [31:0] _RAND_3;
  reg  dec_split; // @[FetchInst.scala 35:27:@722.4]
  reg [31:0] _RAND_4;
  reg  dec_first; // @[FetchInst.scala 36:23:@723.4]
  reg [31:0] _RAND_5;
  reg [31:0] dec_reg_pc; // @[FetchInst.scala 37:23:@724.4]
  reg [31:0] _RAND_6;
  wire  _T_244; // @[FetchInst.scala 40:29:@727.6]
  wire  _T_247; // @[FetchInst.scala 40:19:@729.6]
  wire  _GEN_0; // @[FetchInst.scala 38:27:@725.4]
  wire  _T_250; // @[FetchInst.scala 44:42:@734.4]
  wire  _T_251; // @[FetchInst.scala 44:39:@735.4]
  wire  _T_252; // @[FetchInst.scala 44:64:@736.4]
  wire  _T_254; // @[FetchInst.scala 44:80:@737.4]
  wire  serial; // @[FetchInst.scala 44:77:@738.4]
  reg  _T_257; // @[BackEnd.scala 66:27:@739.4]
  reg [31:0] _RAND_7;
  wire  _GEN_3; // @[BackEnd.scala 68:20:@744.6]
  wire  _GEN_4; // @[BackEnd.scala 67:20:@740.4]
  wire  dec_serial; // @[BackEnd.scala 69:8:@747.4]
  wire [28:0] _T_260; // @[FrontEnd.scala 9:13:@748.4]
  wire [31:0] _T_264; // @[Cat.scala 30:58:@750.4]
  wire [31:0] _T_265; // @[FetchInst.scala 48:10:@751.4]
  wire [31:0] if_pc_next; // @[FetchInst.scala 47:8:@752.4]
  wire  _T_266; // @[FetchInst.scala 51:20:@753.4]
  wire  _T_267; // @[FetchInst.scala 51:34:@754.4]
  wire [31:0] _GEN_5; // @[FetchInst.scala 51:55:@755.4]
  wire  _T_272; // @[FetchInst.scala 57:15:@761.4]
  wire  _T_273; // @[FetchInst.scala 57:57:@762.4]
  wire  _T_274; // @[FetchInst.scala 57:40:@763.4]
  wire  _T_275; // @[FetchInst.scala 55:45:@764.4]
  wire  dec_forward; // @[FetchInst.scala 55:39:@765.4]
  wire  inst_ready; // @[FetchInst.scala 59:23:@766.4]
  wire  _T_276; // @[FetchInst.scala 64:70:@767.4]
  wire  _T_277; // @[FetchInst.scala 64:58:@768.4]
  wire  _T_279; // @[FetchInst.scala 62:5:@769.4]
  wire  _T_280; // @[FetchInst.scala 62:18:@770.4]
  wire  _T_281; // @[FetchInst.scala 62:39:@771.4]
  wire  _T_285; // @[FetchInst.scala 66:50:@775.4]
  wire  _T_286; // @[FetchInst.scala 66:62:@776.4]
  wire  _T_291; // @[FetchInst.scala 62:39:@781.4]
  wire  _T_294; // @[FetchInst.scala 69:41:@784.4]
  wire  _T_295; // @[FetchInst.scala 69:38:@785.4]
  wire  _T_298; // @[FetchInst.scala 69:53:@787.4]
  wire  addr_ready; // @[FetchInst.scala 69:69:@788.4]
  wire  _T_299; // @[Conditional.scala 37:30:@789.4]
  wire  _GEN_6; // @[FetchInst.scala 71:40:@791.6]
  wire  _T_303; // @[FetchInst.scala 75:34:@800.10]
  wire  _GEN_7; // @[FetchInst.scala 74:39:@798.8]
  wire  _GEN_8; // @[Conditional.scala 39:67:@797.6]
  wire  _GEN_9; // @[Conditional.scala 40:58:@790.4]
  wire  inst_valid_0; // @[FetchInst.scala 80:43:@807.4]
  wire  _T_315; // @[FetchInst.scala 81:58:@810.4]
  wire  _T_317; // @[FetchInst.scala 81:46:@811.4]
  wire  inst_valid_1; // @[FetchInst.scala 81:43:@812.4]
  wire  inst_vec_1; // @[FetchInst.scala 86:18:@817.4]
  wire  inst_back_0; // @[FetchInst.scala 88:35:@819.4]
  wire  _T_336; // @[Conditional.scala 37:30:@821.4]
  wire  _T_338; // @[FetchInst.scala 92:29:@825.8]
  wire  _T_340; // @[FetchInst.scala 92:58:@826.8]
  wire  _T_341; // @[FetchInst.scala 92:55:@827.8]
  wire [1:0] _GEN_10; // @[FetchInst.scala 92:81:@828.8]
  wire  _T_343; // @[FetchInst.scala 94:45:@833.8]
  wire  _T_344; // @[FetchInst.scala 94:42:@834.8]
  wire [1:0] _GEN_11; // @[FetchInst.scala 94:65:@835.8]
  wire [1:0] _GEN_12; // @[FetchInst.scala 91:31:@823.6]
  wire  _T_345; // @[Conditional.scala 37:30:@841.6]
  wire  _T_346; // @[FetchInst.scala 99:33:@843.8]
  wire [1:0] _GEN_13; // @[FetchInst.scala 99:52:@844.8]
  wire  _T_347; // @[Conditional.scala 37:30:@849.8]
  wire [1:0] _GEN_14; // @[FetchInst.scala 104:37:@851.10]
  wire [1:0] _GEN_15; // @[Conditional.scala 39:67:@850.8]
  wire [1:0] _GEN_16; // @[Conditional.scala 39:67:@842.6]
  wire [1:0] _GEN_17; // @[Conditional.scala 40:58:@822.4]
  wire  inst_back_1; // @[FetchInst.scala 88:35:@855.4]
  wire  _T_349; // @[Conditional.scala 37:30:@857.4]
  wire  _T_351; // @[FetchInst.scala 92:29:@861.8]
  wire  _T_354; // @[FetchInst.scala 92:55:@863.8]
  wire [1:0] _GEN_18; // @[FetchInst.scala 92:81:@864.8]
  wire  _T_356; // @[FetchInst.scala 94:45:@869.8]
  wire  _T_357; // @[FetchInst.scala 94:42:@870.8]
  wire [1:0] _GEN_19; // @[FetchInst.scala 94:65:@871.8]
  wire [1:0] _GEN_20; // @[FetchInst.scala 91:31:@859.6]
  wire  _T_358; // @[Conditional.scala 37:30:@877.6]
  wire  _T_359; // @[FetchInst.scala 99:33:@879.8]
  wire [1:0] _GEN_21; // @[FetchInst.scala 99:52:@880.8]
  wire  _T_360; // @[Conditional.scala 37:30:@885.8]
  wire [1:0] _GEN_22; // @[FetchInst.scala 104:37:@887.10]
  wire [1:0] _GEN_23; // @[Conditional.scala 39:67:@886.8]
  wire [1:0] _GEN_24; // @[Conditional.scala 39:67:@878.6]
  wire [1:0] _GEN_25; // @[Conditional.scala 40:58:@858.4]
  reg [31:0] reg_inst_0; // @[FetchInst.scala 111:21:@891.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_inst_1; // @[FetchInst.scala 111:21:@891.4]
  reg [31:0] _RAND_9;
  wire  _T_368; // @[FetchInst.scala 116:47:@895.4]
  wire  _T_370; // @[FetchInst.scala 117:43:@898.4]
  wire  _T_371; // @[FetchInst.scala 117:53:@899.4]
  wire  _T_374; // @[FetchInst.scala 116:47:@906.4]
  wire  _T_377; // @[FetchInst.scala 117:53:@910.4]
  wire  _T_381; // @[FetchInst.scala 120:18:@914.4]
  wire  _T_383; // @[FetchInst.scala 120:37:@915.4]
  wire  _T_384; // @[FetchInst.scala 120:27:@916.4]
  wire [7:0] _T_388; // @[FetchInst.scala 127:14:@919.6]
  wire  _T_392; // @[FetchInst.scala 135:26:@921.6]
  wire [7:0] _T_394; // @[Mux.scala 61:16:@922.6]
  wire [7:0] _T_395; // @[Mux.scala 61:16:@923.6]
  wire  _T_399; // @[FetchInst.scala 139:26:@925.6]
  wire [7:0] _T_401; // @[Mux.scala 61:16:@926.6]
  wire [7:0] _T_402; // @[Mux.scala 61:16:@927.6]
  wire [31:0] _T_403; // @[FetchInst.scala 145:14:@928.6]
  wire [31:0] _T_404; // @[FetchInst.scala 146:14:@929.6]
  wire  _T_407; // @[FetchInst.scala 121:13:@931.6]
  assign _T_244 = if_reg_pc[2]; // @[FetchInst.scala 40:29:@727.6]
  assign _T_247 = _T_244 == 1'h0; // @[FetchInst.scala 40:19:@729.6]
  assign _GEN_0 = io_if_forward_1 ? io_if_split : dec_split; // @[FetchInst.scala 38:27:@725.4]
  assign _T_250 = io_mem_inst_1_valid == 1'h0; // @[FetchInst.scala 44:42:@734.4]
  assign _T_251 = pc_state & _T_250; // @[FetchInst.scala 44:39:@735.4]
  assign _T_252 = _T_251 & dec_first; // @[FetchInst.scala 44:64:@736.4]
  assign _T_254 = dec_split == 1'h0; // @[FetchInst.scala 44:80:@737.4]
  assign serial = _T_252 & _T_254; // @[FetchInst.scala 44:77:@738.4]
  assign _GEN_3 = serial ? 1'h0 : _T_257; // @[BackEnd.scala 68:20:@744.6]
  assign _GEN_4 = io_mem_inst_0_valid ? 1'h1 : _GEN_3; // @[BackEnd.scala 67:20:@740.4]
  assign dec_serial = serial & _T_257; // @[BackEnd.scala 69:8:@747.4]
  assign _T_260 = dec_reg_pc[31:3]; // @[FrontEnd.scala 9:13:@748.4]
  assign _T_264 = {_T_260,1'h1,2'h0}; // @[Cat.scala 30:58:@750.4]
  assign _T_265 = dec_serial ? _T_264 : io_btb_target; // @[FetchInst.scala 48:10:@751.4]
  assign if_pc_next = io_if_kill ? io_if_target : _T_265; // @[FetchInst.scala 47:8:@752.4]
  assign _T_266 = io_if_kill | dec_serial; // @[FetchInst.scala 51:20:@753.4]
  assign _T_267 = _T_266 | io_if_forward_1; // @[FetchInst.scala 51:34:@754.4]
  assign _GEN_5 = _T_267 ? if_pc_next : if_reg_pc; // @[FetchInst.scala 51:55:@755.4]
  assign _T_272 = dec_first & _T_250; // @[FetchInst.scala 57:15:@761.4]
  assign _T_273 = inst_state_1 == 2'h0; // @[FetchInst.scala 57:57:@762.4]
  assign _T_274 = _T_272 & _T_273; // @[FetchInst.scala 57:40:@763.4]
  assign _T_275 = dec_split ? _T_244 : _T_274; // @[FetchInst.scala 55:45:@764.4]
  assign dec_forward = io_dec_forward_1 | _T_275; // @[FetchInst.scala 55:39:@765.4]
  assign inst_ready = dec_first ? io_mem_inst_0_valid : io_mem_inst_1_valid; // @[FetchInst.scala 59:23:@766.4]
  assign _T_276 = pc_state == 1'h0; // @[FetchInst.scala 64:70:@767.4]
  assign _T_277 = io_mem_inst_0_valid | _T_276; // @[FetchInst.scala 64:58:@768.4]
  assign _T_279 = io_if_fence == 1'h0; // @[FetchInst.scala 62:5:@769.4]
  assign _T_280 = _T_279 & io_mem_addr_ready; // @[FetchInst.scala 62:18:@770.4]
  assign _T_281 = _T_280 & _T_277; // @[FetchInst.scala 62:39:@771.4]
  assign _T_285 = dec_serial == 1'h0; // @[FetchInst.scala 66:50:@775.4]
  assign _T_286 = _T_285 & inst_ready; // @[FetchInst.scala 66:62:@776.4]
  assign _T_291 = _T_280 & io_mem_addr_valid; // @[FetchInst.scala 62:39:@781.4]
  assign _T_294 = io_if_kill == 1'h0; // @[FetchInst.scala 69:41:@784.4]
  assign _T_295 = io_mem_addr_ready & _T_294; // @[FetchInst.scala 69:38:@785.4]
  assign _T_298 = _T_295 & _T_279; // @[FetchInst.scala 69:53:@787.4]
  assign addr_ready = _T_298 & dec_forward; // @[FetchInst.scala 69:69:@788.4]
  assign _T_299 = 1'h0 == pc_state; // @[Conditional.scala 37:30:@789.4]
  assign _GEN_6 = addr_ready ? 1'h1 : pc_state; // @[FetchInst.scala 71:40:@791.6]
  assign _T_303 = addr_ready & _T_285; // @[FetchInst.scala 75:34:@800.10]
  assign _GEN_7 = inst_ready ? _T_303 : pc_state; // @[FetchInst.scala 74:39:@798.8]
  assign _GEN_8 = pc_state ? _GEN_7 : pc_state; // @[Conditional.scala 39:67:@797.6]
  assign _GEN_9 = _T_299 ? _GEN_6 : _GEN_8; // @[Conditional.scala 40:58:@790.4]
  assign inst_valid_0 = pc_state & dec_first; // @[FetchInst.scala 80:43:@807.4]
  assign _T_315 = dec_first & dec_split; // @[FetchInst.scala 81:58:@810.4]
  assign _T_317 = _T_315 == 1'h0; // @[FetchInst.scala 81:46:@811.4]
  assign inst_valid_1 = pc_state & _T_317; // @[FetchInst.scala 81:43:@812.4]
  assign inst_vec_1 = dec_first == 1'h0; // @[FetchInst.scala 86:18:@817.4]
  assign inst_back_0 = inst_valid_0 & io_mem_inst_0_valid; // @[FetchInst.scala 88:35:@819.4]
  assign _T_336 = 2'h0 == inst_state_0; // @[Conditional.scala 37:30:@821.4]
  assign _T_338 = dec_first & pc_state; // @[FetchInst.scala 92:29:@825.8]
  assign _T_340 = io_mem_inst_0_valid == 1'h0; // @[FetchInst.scala 92:58:@826.8]
  assign _T_341 = _T_338 & _T_340; // @[FetchInst.scala 92:55:@827.8]
  assign _GEN_10 = _T_341 ? 2'h2 : inst_state_0; // @[FetchInst.scala 92:81:@828.8]
  assign _T_343 = io_dec_forward_0 == 1'h0; // @[FetchInst.scala 94:45:@833.8]
  assign _T_344 = inst_back_0 & _T_343; // @[FetchInst.scala 94:42:@834.8]
  assign _GEN_11 = _T_344 ? 2'h1 : inst_state_0; // @[FetchInst.scala 94:65:@835.8]
  assign _GEN_12 = io_dec_kill_0 ? _GEN_10 : _GEN_11; // @[FetchInst.scala 91:31:@823.6]
  assign _T_345 = 2'h1 == inst_state_0; // @[Conditional.scala 37:30:@841.6]
  assign _T_346 = io_dec_forward_0 | io_dec_kill_0; // @[FetchInst.scala 99:33:@843.8]
  assign _GEN_13 = _T_346 ? 2'h0 : inst_state_0; // @[FetchInst.scala 99:52:@844.8]
  assign _T_347 = 2'h2 == inst_state_0; // @[Conditional.scala 37:30:@849.8]
  assign _GEN_14 = io_mem_inst_0_valid ? 2'h0 : inst_state_0; // @[FetchInst.scala 104:37:@851.10]
  assign _GEN_15 = _T_347 ? _GEN_14 : inst_state_0; // @[Conditional.scala 39:67:@850.8]
  assign _GEN_16 = _T_345 ? _GEN_13 : _GEN_15; // @[Conditional.scala 39:67:@842.6]
  assign _GEN_17 = _T_336 ? _GEN_12 : _GEN_16; // @[Conditional.scala 40:58:@822.4]
  assign inst_back_1 = inst_valid_1 & io_mem_inst_1_valid; // @[FetchInst.scala 88:35:@855.4]
  assign _T_349 = 2'h0 == inst_state_1; // @[Conditional.scala 37:30:@857.4]
  assign _T_351 = inst_vec_1 & pc_state; // @[FetchInst.scala 92:29:@861.8]
  assign _T_354 = _T_351 & _T_250; // @[FetchInst.scala 92:55:@863.8]
  assign _GEN_18 = _T_354 ? 2'h2 : inst_state_1; // @[FetchInst.scala 92:81:@864.8]
  assign _T_356 = io_dec_forward_1 == 1'h0; // @[FetchInst.scala 94:45:@869.8]
  assign _T_357 = inst_back_1 & _T_356; // @[FetchInst.scala 94:42:@870.8]
  assign _GEN_19 = _T_357 ? 2'h1 : inst_state_1; // @[FetchInst.scala 94:65:@871.8]
  assign _GEN_20 = io_dec_kill_1 ? _GEN_18 : _GEN_19; // @[FetchInst.scala 91:31:@859.6]
  assign _T_358 = 2'h1 == inst_state_1; // @[Conditional.scala 37:30:@877.6]
  assign _T_359 = io_dec_forward_1 | io_dec_kill_1; // @[FetchInst.scala 99:33:@879.8]
  assign _GEN_21 = _T_359 ? 2'h0 : inst_state_1; // @[FetchInst.scala 99:52:@880.8]
  assign _T_360 = 2'h2 == inst_state_1; // @[Conditional.scala 37:30:@885.8]
  assign _GEN_22 = io_mem_inst_1_valid ? 2'h0 : inst_state_1; // @[FetchInst.scala 104:37:@887.10]
  assign _GEN_23 = _T_360 ? _GEN_22 : inst_state_1; // @[Conditional.scala 39:67:@886.8]
  assign _GEN_24 = _T_358 ? _GEN_21 : _GEN_23; // @[Conditional.scala 39:67:@878.6]
  assign _GEN_25 = _T_349 ? _GEN_20 : _GEN_24; // @[Conditional.scala 40:58:@858.4]
  assign _T_368 = inst_state_0 == 2'h1; // @[FetchInst.scala 116:47:@895.4]
  assign _T_370 = inst_state_0 == 2'h0; // @[FetchInst.scala 117:43:@898.4]
  assign _T_371 = _T_370 & inst_back_0; // @[FetchInst.scala 117:53:@899.4]
  assign _T_374 = inst_state_1 == 2'h1; // @[FetchInst.scala 116:47:@906.4]
  assign _T_377 = _T_273 & inst_back_1; // @[FetchInst.scala 117:53:@910.4]
  assign _T_381 = io_cyc <= 32'h186; // @[FetchInst.scala 120:18:@914.4]
  assign _T_383 = io_cyc >= 32'h16c; // @[FetchInst.scala 120:37:@915.4]
  assign _T_384 = _T_381 & _T_383; // @[FetchInst.scala 120:27:@916.4]
  assign _T_388 = _T_276 ? 8'h41 : 8'h49; // @[FetchInst.scala 127:14:@919.6]
  assign _T_392 = inst_state_0 == 2'h2; // @[FetchInst.scala 135:26:@921.6]
  assign _T_394 = _T_392 ? 8'h43 : 8'h57; // @[Mux.scala 61:16:@922.6]
  assign _T_395 = _T_368 ? 8'h52 : _T_394; // @[Mux.scala 61:16:@923.6]
  assign _T_399 = inst_state_1 == 2'h2; // @[FetchInst.scala 139:26:@925.6]
  assign _T_401 = _T_399 ? 8'h43 : 8'h57; // @[Mux.scala 61:16:@926.6]
  assign _T_402 = _T_374 ? 8'h52 : _T_401; // @[Mux.scala 61:16:@927.6]
  assign _T_403 = io_dec_inst_0_valid ? io_dec_inst_0_bits : 32'h4033; // @[FetchInst.scala 145:14:@928.6]
  assign _T_404 = io_dec_inst_1_valid ? io_dec_inst_1_bits : 32'h4033; // @[FetchInst.scala 146:14:@929.6]
  assign _T_407 = reset == 1'h0; // @[FetchInst.scala 121:13:@931.6]
  assign io_mem_addr_valid = _T_276 | _T_286; // @[FetchInst.scala 66:21:@778.4]
  assign io_mem_addr_bits = if_reg_pc; // @[FetchInst.scala 32:21:@720.4]
  assign io_if_pc = if_reg_pc; // @[FetchInst.scala 33:21:@721.4]
  assign io_if_forward_0 = _T_281 & io_dec_forward_1; // @[FetchInst.scala 64:20:@773.4]
  assign io_if_forward_1 = _T_291 & dec_forward; // @[FetchInst.scala 67:20:@783.4]
  assign io_dec_inst_0_valid = _T_371 | _T_368; // @[FetchInst.scala 117:26:@902.4]
  assign io_dec_inst_0_bits = _T_368 ? reg_inst_0 : io_mem_inst_0_bits; // @[FetchInst.scala 116:26:@897.4]
  assign io_dec_inst_1_valid = _T_377 | _T_374; // @[FetchInst.scala 117:26:@913.4]
  assign io_dec_inst_1_bits = _T_374 ? reg_inst_1 : io_mem_inst_1_bits; // @[FetchInst.scala 116:26:@908.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  pc_state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  inst_state_0 = _RAND_1[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inst_state_1 = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  if_reg_pc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  dec_split = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  dec_first = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  dec_reg_pc = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  _T_257 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_inst_0 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_inst_1 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      pc_state <= 1'h0;
    end else begin
      if (_T_299) begin
        if (addr_ready) begin
          pc_state <= 1'h1;
        end
      end else begin
        if (pc_state) begin
          if (inst_ready) begin
            pc_state <= _T_303;
          end
        end
      end
    end
    if (reset) begin
      inst_state_0 <= 2'h0;
    end else begin
      if (_T_336) begin
        if (io_dec_kill_0) begin
          if (_T_341) begin
            inst_state_0 <= 2'h2;
          end
        end else begin
          if (_T_344) begin
            inst_state_0 <= 2'h1;
          end
        end
      end else begin
        if (_T_345) begin
          if (_T_346) begin
            inst_state_0 <= 2'h0;
          end
        end else begin
          if (_T_347) begin
            if (io_mem_inst_0_valid) begin
              inst_state_0 <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      inst_state_1 <= 2'h0;
    end else begin
      if (_T_349) begin
        if (io_dec_kill_1) begin
          if (_T_354) begin
            inst_state_1 <= 2'h2;
          end
        end else begin
          if (_T_357) begin
            inst_state_1 <= 2'h1;
          end
        end
      end else begin
        if (_T_358) begin
          if (_T_359) begin
            inst_state_1 <= 2'h0;
          end
        end else begin
          if (_T_360) begin
            if (io_mem_inst_1_valid) begin
              inst_state_1 <= 2'h0;
            end
          end
        end
      end
    end
    if (reset) begin
      if_reg_pc <= 32'h80000000;
    end else begin
      if (_T_267) begin
        if (io_if_kill) begin
          if_reg_pc <= io_if_target;
        end else begin
          if (dec_serial) begin
            if_reg_pc <= _T_264;
          end else begin
            if_reg_pc <= io_btb_target;
          end
        end
      end
    end
    if (reset) begin
      dec_split <= 1'h0;
    end else begin
      if (io_if_forward_1) begin
        dec_split <= io_if_split;
      end
    end
    if (io_if_forward_1) begin
      dec_first <= _T_247;
    end
    if (io_if_forward_1) begin
      dec_reg_pc <= if_reg_pc;
    end
    if (reset) begin
      _T_257 <= 1'h1;
    end else begin
      if (io_mem_inst_0_valid) begin
        _T_257 <= 1'h1;
      end else begin
        if (serial) begin
          _T_257 <= 1'h0;
        end
      end
    end
    if (inst_back_0) begin
      reg_inst_0 <= io_mem_inst_0_bits;
    end
    if (inst_back_1) begin
      reg_inst_1 <= io_mem_inst_1_bits;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_384 & _T_407) begin
          $fwrite(32'h80000002,"FetchInst: Cyc= %d if_reg_pc %x pc_valid %x pc_ready %x pc_state %c pc_forward %x %x dec_pc %x dec_forward %x %x inst_state %c %c inst_valid %x:%x %x:%x inst = DASM(%x) DASM(%x)\n",io_cyc,if_reg_pc,io_mem_addr_valid,io_mem_addr_ready,_T_388,io_if_forward_0,io_if_forward_1,dec_reg_pc,io_dec_forward_0,io_dec_forward_1,_T_395,_T_402,io_mem_inst_0_valid,io_dec_inst_0_valid,io_mem_inst_1_valid,io_dec_inst_1_valid,_T_403,_T_404); // @[FetchInst.scala 121:13:@933.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module BTB( // @[:@937.2]
  input         clock, // @[:@938.4]
  input         reset, // @[:@939.4]
  input  [31:0] io_if_pc, // @[:@940.4]
  input  [31:0] io_ras_peek, // @[:@940.4]
  output [31:0] io_pred_pc_0, // @[:@940.4]
  output [31:0] io_pred_pc_1, // @[:@940.4]
  output        io_split, // @[:@940.4]
  input  [31:0] io_fb_pc, // @[:@940.4]
  input  [1:0]  io_fb_type, // @[:@940.4]
  input         io_feedBack_valid, // @[:@940.4]
  input         io_feedBack_bits_redirect, // @[:@940.4]
  input  [31:0] io_feedBack_bits_tgt // @[:@940.4]
);
  reg [31:0] btb_pc_0; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_0;
  reg [31:0] btb_pc_1; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_1;
  reg [31:0] btb_pc_2; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_2;
  reg [31:0] btb_pc_3; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_3;
  reg [31:0] btb_pc_4; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_4;
  reg [31:0] btb_pc_5; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_5;
  reg [31:0] btb_pc_6; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_6;
  reg [31:0] btb_pc_7; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_7;
  reg [31:0] btb_pc_8; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_8;
  reg [31:0] btb_pc_9; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_9;
  reg [31:0] btb_pc_10; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_10;
  reg [31:0] btb_pc_11; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_11;
  reg [31:0] btb_pc_12; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_12;
  reg [31:0] btb_pc_13; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_13;
  reg [31:0] btb_pc_14; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_14;
  reg [31:0] btb_pc_15; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_15;
  reg [31:0] btb_pc_16; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_16;
  reg [31:0] btb_pc_17; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_17;
  reg [31:0] btb_pc_18; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_18;
  reg [31:0] btb_pc_19; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_19;
  reg [31:0] btb_pc_20; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_20;
  reg [31:0] btb_pc_21; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_21;
  reg [31:0] btb_pc_22; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_22;
  reg [31:0] btb_pc_23; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_23;
  reg [31:0] btb_pc_24; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_24;
  reg [31:0] btb_pc_25; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_25;
  reg [31:0] btb_pc_26; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_26;
  reg [31:0] btb_pc_27; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_27;
  reg [31:0] btb_pc_28; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_28;
  reg [31:0] btb_pc_29; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_29;
  reg [31:0] btb_pc_30; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_30;
  reg [31:0] btb_pc_31; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_31;
  reg [31:0] btb_pc_32; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_32;
  reg [31:0] btb_pc_33; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_33;
  reg [31:0] btb_pc_34; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_34;
  reg [31:0] btb_pc_35; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_35;
  reg [31:0] btb_pc_36; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_36;
  reg [31:0] btb_pc_37; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_37;
  reg [31:0] btb_pc_38; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_38;
  reg [31:0] btb_pc_39; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_39;
  reg [31:0] btb_pc_40; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_40;
  reg [31:0] btb_pc_41; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_41;
  reg [31:0] btb_pc_42; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_42;
  reg [31:0] btb_pc_43; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_43;
  reg [31:0] btb_pc_44; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_44;
  reg [31:0] btb_pc_45; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_45;
  reg [31:0] btb_pc_46; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_46;
  reg [31:0] btb_pc_47; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_47;
  reg [31:0] btb_pc_48; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_48;
  reg [31:0] btb_pc_49; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_49;
  reg [31:0] btb_pc_50; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_50;
  reg [31:0] btb_pc_51; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_51;
  reg [31:0] btb_pc_52; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_52;
  reg [31:0] btb_pc_53; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_53;
  reg [31:0] btb_pc_54; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_54;
  reg [31:0] btb_pc_55; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_55;
  reg [31:0] btb_pc_56; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_56;
  reg [31:0] btb_pc_57; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_57;
  reg [31:0] btb_pc_58; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_58;
  reg [31:0] btb_pc_59; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_59;
  reg [31:0] btb_pc_60; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_60;
  reg [31:0] btb_pc_61; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_61;
  reg [31:0] btb_pc_62; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_62;
  reg [31:0] btb_pc_63; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_63;
  reg [31:0] btb_target_0; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_64;
  reg [31:0] btb_target_1; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_65;
  reg [31:0] btb_target_2; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_66;
  reg [31:0] btb_target_3; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_67;
  reg [31:0] btb_target_4; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_68;
  reg [31:0] btb_target_5; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_69;
  reg [31:0] btb_target_6; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_70;
  reg [31:0] btb_target_7; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_71;
  reg [31:0] btb_target_8; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_72;
  reg [31:0] btb_target_9; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_73;
  reg [31:0] btb_target_10; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_74;
  reg [31:0] btb_target_11; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_75;
  reg [31:0] btb_target_12; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_76;
  reg [31:0] btb_target_13; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_77;
  reg [31:0] btb_target_14; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_78;
  reg [31:0] btb_target_15; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_79;
  reg [31:0] btb_target_16; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_80;
  reg [31:0] btb_target_17; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_81;
  reg [31:0] btb_target_18; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_82;
  reg [31:0] btb_target_19; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_83;
  reg [31:0] btb_target_20; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_84;
  reg [31:0] btb_target_21; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_85;
  reg [31:0] btb_target_22; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_86;
  reg [31:0] btb_target_23; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_87;
  reg [31:0] btb_target_24; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_88;
  reg [31:0] btb_target_25; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_89;
  reg [31:0] btb_target_26; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_90;
  reg [31:0] btb_target_27; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_91;
  reg [31:0] btb_target_28; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_92;
  reg [31:0] btb_target_29; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_93;
  reg [31:0] btb_target_30; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_94;
  reg [31:0] btb_target_31; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_95;
  reg [31:0] btb_target_32; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_96;
  reg [31:0] btb_target_33; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_97;
  reg [31:0] btb_target_34; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_98;
  reg [31:0] btb_target_35; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_99;
  reg [31:0] btb_target_36; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_100;
  reg [31:0] btb_target_37; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_101;
  reg [31:0] btb_target_38; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_102;
  reg [31:0] btb_target_39; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_103;
  reg [31:0] btb_target_40; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_104;
  reg [31:0] btb_target_41; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_105;
  reg [31:0] btb_target_42; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_106;
  reg [31:0] btb_target_43; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_107;
  reg [31:0] btb_target_44; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_108;
  reg [31:0] btb_target_45; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_109;
  reg [31:0] btb_target_46; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_110;
  reg [31:0] btb_target_47; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_111;
  reg [31:0] btb_target_48; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_112;
  reg [31:0] btb_target_49; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_113;
  reg [31:0] btb_target_50; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_114;
  reg [31:0] btb_target_51; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_115;
  reg [31:0] btb_target_52; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_116;
  reg [31:0] btb_target_53; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_117;
  reg [31:0] btb_target_54; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_118;
  reg [31:0] btb_target_55; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_119;
  reg [31:0] btb_target_56; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_120;
  reg [31:0] btb_target_57; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_121;
  reg [31:0] btb_target_58; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_122;
  reg [31:0] btb_target_59; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_123;
  reg [31:0] btb_target_60; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_124;
  reg [31:0] btb_target_61; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_125;
  reg [31:0] btb_target_62; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_126;
  reg [31:0] btb_target_63; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_127;
  reg [1:0] btb_hcount_0; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_128;
  reg [1:0] btb_hcount_1; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_129;
  reg [1:0] btb_hcount_2; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_130;
  reg [1:0] btb_hcount_3; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_131;
  reg [1:0] btb_hcount_4; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_132;
  reg [1:0] btb_hcount_5; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_133;
  reg [1:0] btb_hcount_6; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_134;
  reg [1:0] btb_hcount_7; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_135;
  reg [1:0] btb_hcount_8; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_136;
  reg [1:0] btb_hcount_9; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_137;
  reg [1:0] btb_hcount_10; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_138;
  reg [1:0] btb_hcount_11; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_139;
  reg [1:0] btb_hcount_12; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_140;
  reg [1:0] btb_hcount_13; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_141;
  reg [1:0] btb_hcount_14; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_142;
  reg [1:0] btb_hcount_15; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_143;
  reg [1:0] btb_hcount_16; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_144;
  reg [1:0] btb_hcount_17; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_145;
  reg [1:0] btb_hcount_18; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_146;
  reg [1:0] btb_hcount_19; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_147;
  reg [1:0] btb_hcount_20; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_148;
  reg [1:0] btb_hcount_21; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_149;
  reg [1:0] btb_hcount_22; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_150;
  reg [1:0] btb_hcount_23; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_151;
  reg [1:0] btb_hcount_24; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_152;
  reg [1:0] btb_hcount_25; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_153;
  reg [1:0] btb_hcount_26; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_154;
  reg [1:0] btb_hcount_27; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_155;
  reg [1:0] btb_hcount_28; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_156;
  reg [1:0] btb_hcount_29; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_157;
  reg [1:0] btb_hcount_30; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_158;
  reg [1:0] btb_hcount_31; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_159;
  reg [1:0] btb_hcount_32; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_160;
  reg [1:0] btb_hcount_33; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_161;
  reg [1:0] btb_hcount_34; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_162;
  reg [1:0] btb_hcount_35; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_163;
  reg [1:0] btb_hcount_36; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_164;
  reg [1:0] btb_hcount_37; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_165;
  reg [1:0] btb_hcount_38; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_166;
  reg [1:0] btb_hcount_39; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_167;
  reg [1:0] btb_hcount_40; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_168;
  reg [1:0] btb_hcount_41; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_169;
  reg [1:0] btb_hcount_42; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_170;
  reg [1:0] btb_hcount_43; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_171;
  reg [1:0] btb_hcount_44; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_172;
  reg [1:0] btb_hcount_45; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_173;
  reg [1:0] btb_hcount_46; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_174;
  reg [1:0] btb_hcount_47; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_175;
  reg [1:0] btb_hcount_48; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_176;
  reg [1:0] btb_hcount_49; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_177;
  reg [1:0] btb_hcount_50; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_178;
  reg [1:0] btb_hcount_51; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_179;
  reg [1:0] btb_hcount_52; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_180;
  reg [1:0] btb_hcount_53; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_181;
  reg [1:0] btb_hcount_54; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_182;
  reg [1:0] btb_hcount_55; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_183;
  reg [1:0] btb_hcount_56; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_184;
  reg [1:0] btb_hcount_57; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_185;
  reg [1:0] btb_hcount_58; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_186;
  reg [1:0] btb_hcount_59; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_187;
  reg [1:0] btb_hcount_60; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_188;
  reg [1:0] btb_hcount_61; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_189;
  reg [1:0] btb_hcount_62; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_190;
  reg [1:0] btb_hcount_63; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_191;
  reg [1:0] btb_btype_0; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_192;
  reg [1:0] btb_btype_1; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_193;
  reg [1:0] btb_btype_2; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_194;
  reg [1:0] btb_btype_3; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_195;
  reg [1:0] btb_btype_4; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_196;
  reg [1:0] btb_btype_5; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_197;
  reg [1:0] btb_btype_6; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_198;
  reg [1:0] btb_btype_7; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_199;
  reg [1:0] btb_btype_8; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_200;
  reg [1:0] btb_btype_9; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_201;
  reg [1:0] btb_btype_10; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_202;
  reg [1:0] btb_btype_11; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_203;
  reg [1:0] btb_btype_12; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_204;
  reg [1:0] btb_btype_13; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_205;
  reg [1:0] btb_btype_14; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_206;
  reg [1:0] btb_btype_15; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_207;
  reg [1:0] btb_btype_16; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_208;
  reg [1:0] btb_btype_17; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_209;
  reg [1:0] btb_btype_18; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_210;
  reg [1:0] btb_btype_19; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_211;
  reg [1:0] btb_btype_20; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_212;
  reg [1:0] btb_btype_21; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_213;
  reg [1:0] btb_btype_22; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_214;
  reg [1:0] btb_btype_23; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_215;
  reg [1:0] btb_btype_24; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_216;
  reg [1:0] btb_btype_25; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_217;
  reg [1:0] btb_btype_26; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_218;
  reg [1:0] btb_btype_27; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_219;
  reg [1:0] btb_btype_28; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_220;
  reg [1:0] btb_btype_29; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_221;
  reg [1:0] btb_btype_30; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_222;
  reg [1:0] btb_btype_31; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_223;
  reg [1:0] btb_btype_32; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_224;
  reg [1:0] btb_btype_33; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_225;
  reg [1:0] btb_btype_34; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_226;
  reg [1:0] btb_btype_35; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_227;
  reg [1:0] btb_btype_36; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_228;
  reg [1:0] btb_btype_37; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_229;
  reg [1:0] btb_btype_38; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_230;
  reg [1:0] btb_btype_39; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_231;
  reg [1:0] btb_btype_40; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_232;
  reg [1:0] btb_btype_41; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_233;
  reg [1:0] btb_btype_42; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_234;
  reg [1:0] btb_btype_43; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_235;
  reg [1:0] btb_btype_44; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_236;
  reg [1:0] btb_btype_45; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_237;
  reg [1:0] btb_btype_46; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_238;
  reg [1:0] btb_btype_47; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_239;
  reg [1:0] btb_btype_48; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_240;
  reg [1:0] btb_btype_49; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_241;
  reg [1:0] btb_btype_50; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_242;
  reg [1:0] btb_btype_51; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_243;
  reg [1:0] btb_btype_52; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_244;
  reg [1:0] btb_btype_53; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_245;
  reg [1:0] btb_btype_54; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_246;
  reg [1:0] btb_btype_55; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_247;
  reg [1:0] btb_btype_56; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_248;
  reg [1:0] btb_btype_57; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_249;
  reg [1:0] btb_btype_58; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_250;
  reg [1:0] btb_btype_59; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_251;
  reg [1:0] btb_btype_60; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_252;
  reg [1:0] btb_btype_61; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_253;
  reg [1:0] btb_btype_62; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_254;
  reg [1:0] btb_btype_63; // @[BTB.scala 46:20:@1199.4]
  reg [31:0] _RAND_255;
  wire [28:0] _T_152; // @[FrontEnd.scala 9:13:@1202.4]
  wire [31:0] if_pc_0; // @[Cat.scala 30:58:@1204.4]
  wire  _T_157; // @[BTB.scala 76:47:@1206.4]
  wire  _T_158; // @[BTB.scala 76:47:@1207.4]
  wire  _T_159; // @[BTB.scala 76:47:@1208.4]
  wire  _T_160; // @[BTB.scala 76:47:@1209.4]
  wire  _T_161; // @[BTB.scala 76:47:@1210.4]
  wire  _T_162; // @[BTB.scala 76:47:@1211.4]
  wire  _T_163; // @[BTB.scala 76:47:@1212.4]
  wire  _T_164; // @[BTB.scala 76:47:@1213.4]
  wire  _T_165; // @[BTB.scala 76:47:@1214.4]
  wire  _T_166; // @[BTB.scala 76:47:@1215.4]
  wire  _T_167; // @[BTB.scala 76:47:@1216.4]
  wire  _T_168; // @[BTB.scala 76:47:@1217.4]
  wire  _T_169; // @[BTB.scala 76:47:@1218.4]
  wire  _T_170; // @[BTB.scala 76:47:@1219.4]
  wire  _T_171; // @[BTB.scala 76:47:@1220.4]
  wire  _T_172; // @[BTB.scala 76:47:@1221.4]
  wire  _T_173; // @[BTB.scala 76:47:@1222.4]
  wire  _T_174; // @[BTB.scala 76:47:@1223.4]
  wire  _T_175; // @[BTB.scala 76:47:@1224.4]
  wire  _T_176; // @[BTB.scala 76:47:@1225.4]
  wire  _T_177; // @[BTB.scala 76:47:@1226.4]
  wire  _T_178; // @[BTB.scala 76:47:@1227.4]
  wire  _T_179; // @[BTB.scala 76:47:@1228.4]
  wire  _T_180; // @[BTB.scala 76:47:@1229.4]
  wire  _T_181; // @[BTB.scala 76:47:@1230.4]
  wire  _T_182; // @[BTB.scala 76:47:@1231.4]
  wire  _T_183; // @[BTB.scala 76:47:@1232.4]
  wire  _T_184; // @[BTB.scala 76:47:@1233.4]
  wire  _T_185; // @[BTB.scala 76:47:@1234.4]
  wire  _T_186; // @[BTB.scala 76:47:@1235.4]
  wire  _T_187; // @[BTB.scala 76:47:@1236.4]
  wire  _T_188; // @[BTB.scala 76:47:@1237.4]
  wire  _T_189; // @[BTB.scala 76:47:@1238.4]
  wire  _T_190; // @[BTB.scala 76:47:@1239.4]
  wire  _T_191; // @[BTB.scala 76:47:@1240.4]
  wire  _T_192; // @[BTB.scala 76:47:@1241.4]
  wire  _T_193; // @[BTB.scala 76:47:@1242.4]
  wire  _T_194; // @[BTB.scala 76:47:@1243.4]
  wire  _T_195; // @[BTB.scala 76:47:@1244.4]
  wire  _T_196; // @[BTB.scala 76:47:@1245.4]
  wire  _T_197; // @[BTB.scala 76:47:@1246.4]
  wire  _T_198; // @[BTB.scala 76:47:@1247.4]
  wire  _T_199; // @[BTB.scala 76:47:@1248.4]
  wire  _T_200; // @[BTB.scala 76:47:@1249.4]
  wire  _T_201; // @[BTB.scala 76:47:@1250.4]
  wire  _T_202; // @[BTB.scala 76:47:@1251.4]
  wire  _T_203; // @[BTB.scala 76:47:@1252.4]
  wire  _T_204; // @[BTB.scala 76:47:@1253.4]
  wire  _T_205; // @[BTB.scala 76:47:@1254.4]
  wire  _T_206; // @[BTB.scala 76:47:@1255.4]
  wire  _T_207; // @[BTB.scala 76:47:@1256.4]
  wire  _T_208; // @[BTB.scala 76:47:@1257.4]
  wire  _T_209; // @[BTB.scala 76:47:@1258.4]
  wire  _T_210; // @[BTB.scala 76:47:@1259.4]
  wire  _T_211; // @[BTB.scala 76:47:@1260.4]
  wire  _T_212; // @[BTB.scala 76:47:@1261.4]
  wire  _T_213; // @[BTB.scala 76:47:@1262.4]
  wire  _T_214; // @[BTB.scala 76:47:@1263.4]
  wire  _T_215; // @[BTB.scala 76:47:@1264.4]
  wire  _T_216; // @[BTB.scala 76:47:@1265.4]
  wire  _T_217; // @[BTB.scala 76:47:@1266.4]
  wire  _T_218; // @[BTB.scala 76:47:@1267.4]
  wire  _T_219; // @[BTB.scala 76:47:@1268.4]
  wire  _T_220; // @[BTB.scala 76:47:@1269.4]
  wire [7:0] _T_297; // @[BTB.scala 76:62:@1341.4]
  wire [15:0] _T_305; // @[BTB.scala 76:62:@1349.4]
  wire [7:0] _T_312; // @[BTB.scala 76:62:@1356.4]
  wire [31:0] _T_321; // @[BTB.scala 76:62:@1365.4]
  wire [7:0] _T_328; // @[BTB.scala 76:62:@1372.4]
  wire [15:0] _T_336; // @[BTB.scala 76:62:@1380.4]
  wire [7:0] _T_343; // @[BTB.scala 76:62:@1387.4]
  wire [31:0] _T_352; // @[BTB.scala 76:62:@1396.4]
  wire [63:0] _T_353; // @[BTB.scala 76:62:@1397.4]
  wire  _T_355; // @[BTB.scala 52:66:@1398.4]
  wire  _T_357; // @[BTB.scala 52:66:@1399.4]
  wire  _T_359; // @[BTB.scala 52:66:@1400.4]
  wire  _T_361; // @[BTB.scala 52:66:@1401.4]
  wire  _T_363; // @[BTB.scala 52:66:@1402.4]
  wire  _T_365; // @[BTB.scala 52:66:@1403.4]
  wire  _T_367; // @[BTB.scala 52:66:@1404.4]
  wire  _T_369; // @[BTB.scala 52:66:@1405.4]
  wire  _T_371; // @[BTB.scala 52:66:@1406.4]
  wire  _T_373; // @[BTB.scala 52:66:@1407.4]
  wire  _T_375; // @[BTB.scala 52:66:@1408.4]
  wire  _T_377; // @[BTB.scala 52:66:@1409.4]
  wire  _T_379; // @[BTB.scala 52:66:@1410.4]
  wire  _T_381; // @[BTB.scala 52:66:@1411.4]
  wire  _T_383; // @[BTB.scala 52:66:@1412.4]
  wire  _T_385; // @[BTB.scala 52:66:@1413.4]
  wire  _T_387; // @[BTB.scala 52:66:@1414.4]
  wire  _T_389; // @[BTB.scala 52:66:@1415.4]
  wire  _T_391; // @[BTB.scala 52:66:@1416.4]
  wire  _T_393; // @[BTB.scala 52:66:@1417.4]
  wire  _T_395; // @[BTB.scala 52:66:@1418.4]
  wire  _T_397; // @[BTB.scala 52:66:@1419.4]
  wire  _T_399; // @[BTB.scala 52:66:@1420.4]
  wire  _T_401; // @[BTB.scala 52:66:@1421.4]
  wire  _T_403; // @[BTB.scala 52:66:@1422.4]
  wire  _T_405; // @[BTB.scala 52:66:@1423.4]
  wire  _T_407; // @[BTB.scala 52:66:@1424.4]
  wire  _T_409; // @[BTB.scala 52:66:@1425.4]
  wire  _T_411; // @[BTB.scala 52:66:@1426.4]
  wire  _T_413; // @[BTB.scala 52:66:@1427.4]
  wire  _T_415; // @[BTB.scala 52:66:@1428.4]
  wire  _T_417; // @[BTB.scala 52:66:@1429.4]
  wire  _T_419; // @[BTB.scala 52:66:@1430.4]
  wire  _T_421; // @[BTB.scala 52:66:@1431.4]
  wire  _T_423; // @[BTB.scala 52:66:@1432.4]
  wire  _T_425; // @[BTB.scala 52:66:@1433.4]
  wire  _T_427; // @[BTB.scala 52:66:@1434.4]
  wire  _T_429; // @[BTB.scala 52:66:@1435.4]
  wire  _T_431; // @[BTB.scala 52:66:@1436.4]
  wire  _T_433; // @[BTB.scala 52:66:@1437.4]
  wire  _T_435; // @[BTB.scala 52:66:@1438.4]
  wire  _T_437; // @[BTB.scala 52:66:@1439.4]
  wire  _T_439; // @[BTB.scala 52:66:@1440.4]
  wire  _T_441; // @[BTB.scala 52:66:@1441.4]
  wire  _T_443; // @[BTB.scala 52:66:@1442.4]
  wire  _T_445; // @[BTB.scala 52:66:@1443.4]
  wire  _T_447; // @[BTB.scala 52:66:@1444.4]
  wire  _T_449; // @[BTB.scala 52:66:@1445.4]
  wire  _T_451; // @[BTB.scala 52:66:@1446.4]
  wire  _T_453; // @[BTB.scala 52:66:@1447.4]
  wire  _T_455; // @[BTB.scala 52:66:@1448.4]
  wire  _T_457; // @[BTB.scala 52:66:@1449.4]
  wire  _T_459; // @[BTB.scala 52:66:@1450.4]
  wire  _T_461; // @[BTB.scala 52:66:@1451.4]
  wire  _T_463; // @[BTB.scala 52:66:@1452.4]
  wire  _T_465; // @[BTB.scala 52:66:@1453.4]
  wire  _T_467; // @[BTB.scala 52:66:@1454.4]
  wire  _T_469; // @[BTB.scala 52:66:@1455.4]
  wire  _T_471; // @[BTB.scala 52:66:@1456.4]
  wire  _T_473; // @[BTB.scala 52:66:@1457.4]
  wire  _T_475; // @[BTB.scala 52:66:@1458.4]
  wire  _T_477; // @[BTB.scala 52:66:@1459.4]
  wire  _T_479; // @[BTB.scala 52:66:@1460.4]
  wire  _T_481; // @[BTB.scala 52:66:@1461.4]
  wire [7:0] _T_558; // @[BTB.scala 52:72:@1533.4]
  wire [15:0] _T_566; // @[BTB.scala 52:72:@1541.4]
  wire [7:0] _T_573; // @[BTB.scala 52:72:@1548.4]
  wire [31:0] _T_582; // @[BTB.scala 52:72:@1557.4]
  wire [7:0] _T_589; // @[BTB.scala 52:72:@1564.4]
  wire [15:0] _T_597; // @[BTB.scala 52:72:@1572.4]
  wire [7:0] _T_604; // @[BTB.scala 52:72:@1579.4]
  wire [31:0] _T_613; // @[BTB.scala 52:72:@1588.4]
  wire [63:0] _T_614; // @[BTB.scala 52:72:@1589.4]
  wire [63:0] predict_0_lookup; // @[BTB.scala 76:69:@1590.4]
  wire  _T_616; // @[Mux.scala 21:36:@1592.4]
  wire  _T_617; // @[Mux.scala 21:36:@1593.4]
  wire  _T_618; // @[Mux.scala 21:36:@1594.4]
  wire  _T_619; // @[Mux.scala 21:36:@1595.4]
  wire  _T_620; // @[Mux.scala 21:36:@1596.4]
  wire  _T_621; // @[Mux.scala 21:36:@1597.4]
  wire  _T_622; // @[Mux.scala 21:36:@1598.4]
  wire  _T_623; // @[Mux.scala 21:36:@1599.4]
  wire  _T_624; // @[Mux.scala 21:36:@1600.4]
  wire  _T_625; // @[Mux.scala 21:36:@1601.4]
  wire  _T_626; // @[Mux.scala 21:36:@1602.4]
  wire  _T_627; // @[Mux.scala 21:36:@1603.4]
  wire  _T_628; // @[Mux.scala 21:36:@1604.4]
  wire  _T_629; // @[Mux.scala 21:36:@1605.4]
  wire  _T_630; // @[Mux.scala 21:36:@1606.4]
  wire  _T_631; // @[Mux.scala 21:36:@1607.4]
  wire  _T_632; // @[Mux.scala 21:36:@1608.4]
  wire  _T_633; // @[Mux.scala 21:36:@1609.4]
  wire  _T_634; // @[Mux.scala 21:36:@1610.4]
  wire  _T_635; // @[Mux.scala 21:36:@1611.4]
  wire  _T_636; // @[Mux.scala 21:36:@1612.4]
  wire  _T_637; // @[Mux.scala 21:36:@1613.4]
  wire  _T_638; // @[Mux.scala 21:36:@1614.4]
  wire  _T_639; // @[Mux.scala 21:36:@1615.4]
  wire  _T_640; // @[Mux.scala 21:36:@1616.4]
  wire  _T_641; // @[Mux.scala 21:36:@1617.4]
  wire  _T_642; // @[Mux.scala 21:36:@1618.4]
  wire  _T_643; // @[Mux.scala 21:36:@1619.4]
  wire  _T_644; // @[Mux.scala 21:36:@1620.4]
  wire  _T_645; // @[Mux.scala 21:36:@1621.4]
  wire  _T_646; // @[Mux.scala 21:36:@1622.4]
  wire  _T_647; // @[Mux.scala 21:36:@1623.4]
  wire  _T_648; // @[Mux.scala 21:36:@1624.4]
  wire  _T_649; // @[Mux.scala 21:36:@1625.4]
  wire  _T_650; // @[Mux.scala 21:36:@1626.4]
  wire  _T_651; // @[Mux.scala 21:36:@1627.4]
  wire  _T_652; // @[Mux.scala 21:36:@1628.4]
  wire  _T_653; // @[Mux.scala 21:36:@1629.4]
  wire  _T_654; // @[Mux.scala 21:36:@1630.4]
  wire  _T_655; // @[Mux.scala 21:36:@1631.4]
  wire  _T_656; // @[Mux.scala 21:36:@1632.4]
  wire  _T_657; // @[Mux.scala 21:36:@1633.4]
  wire  _T_658; // @[Mux.scala 21:36:@1634.4]
  wire  _T_659; // @[Mux.scala 21:36:@1635.4]
  wire  _T_660; // @[Mux.scala 21:36:@1636.4]
  wire  _T_661; // @[Mux.scala 21:36:@1637.4]
  wire  _T_662; // @[Mux.scala 21:36:@1638.4]
  wire  _T_663; // @[Mux.scala 21:36:@1639.4]
  wire  _T_664; // @[Mux.scala 21:36:@1640.4]
  wire  _T_665; // @[Mux.scala 21:36:@1641.4]
  wire  _T_666; // @[Mux.scala 21:36:@1642.4]
  wire  _T_667; // @[Mux.scala 21:36:@1643.4]
  wire  _T_668; // @[Mux.scala 21:36:@1644.4]
  wire  _T_669; // @[Mux.scala 21:36:@1645.4]
  wire  _T_670; // @[Mux.scala 21:36:@1646.4]
  wire  _T_671; // @[Mux.scala 21:36:@1647.4]
  wire  _T_672; // @[Mux.scala 21:36:@1648.4]
  wire  _T_673; // @[Mux.scala 21:36:@1649.4]
  wire  _T_674; // @[Mux.scala 21:36:@1650.4]
  wire  _T_675; // @[Mux.scala 21:36:@1651.4]
  wire  _T_676; // @[Mux.scala 21:36:@1652.4]
  wire  _T_677; // @[Mux.scala 21:36:@1653.4]
  wire  _T_678; // @[Mux.scala 21:36:@1654.4]
  wire  _T_679; // @[Mux.scala 21:36:@1655.4]
  wire [31:0] _T_682; // @[Mux.scala 19:72:@1656.4]
  wire [31:0] _T_684; // @[Mux.scala 19:72:@1657.4]
  wire [31:0] _T_686; // @[Mux.scala 19:72:@1658.4]
  wire [31:0] _T_688; // @[Mux.scala 19:72:@1659.4]
  wire [31:0] _T_690; // @[Mux.scala 19:72:@1660.4]
  wire [31:0] _T_692; // @[Mux.scala 19:72:@1661.4]
  wire [31:0] _T_694; // @[Mux.scala 19:72:@1662.4]
  wire [31:0] _T_696; // @[Mux.scala 19:72:@1663.4]
  wire [31:0] _T_698; // @[Mux.scala 19:72:@1664.4]
  wire [31:0] _T_700; // @[Mux.scala 19:72:@1665.4]
  wire [31:0] _T_702; // @[Mux.scala 19:72:@1666.4]
  wire [31:0] _T_704; // @[Mux.scala 19:72:@1667.4]
  wire [31:0] _T_706; // @[Mux.scala 19:72:@1668.4]
  wire [31:0] _T_708; // @[Mux.scala 19:72:@1669.4]
  wire [31:0] _T_710; // @[Mux.scala 19:72:@1670.4]
  wire [31:0] _T_712; // @[Mux.scala 19:72:@1671.4]
  wire [31:0] _T_714; // @[Mux.scala 19:72:@1672.4]
  wire [31:0] _T_716; // @[Mux.scala 19:72:@1673.4]
  wire [31:0] _T_718; // @[Mux.scala 19:72:@1674.4]
  wire [31:0] _T_720; // @[Mux.scala 19:72:@1675.4]
  wire [31:0] _T_722; // @[Mux.scala 19:72:@1676.4]
  wire [31:0] _T_724; // @[Mux.scala 19:72:@1677.4]
  wire [31:0] _T_726; // @[Mux.scala 19:72:@1678.4]
  wire [31:0] _T_728; // @[Mux.scala 19:72:@1679.4]
  wire [31:0] _T_730; // @[Mux.scala 19:72:@1680.4]
  wire [31:0] _T_732; // @[Mux.scala 19:72:@1681.4]
  wire [31:0] _T_734; // @[Mux.scala 19:72:@1682.4]
  wire [31:0] _T_736; // @[Mux.scala 19:72:@1683.4]
  wire [31:0] _T_738; // @[Mux.scala 19:72:@1684.4]
  wire [31:0] _T_740; // @[Mux.scala 19:72:@1685.4]
  wire [31:0] _T_742; // @[Mux.scala 19:72:@1686.4]
  wire [31:0] _T_744; // @[Mux.scala 19:72:@1687.4]
  wire [31:0] _T_746; // @[Mux.scala 19:72:@1688.4]
  wire [31:0] _T_748; // @[Mux.scala 19:72:@1689.4]
  wire [31:0] _T_750; // @[Mux.scala 19:72:@1690.4]
  wire [31:0] _T_752; // @[Mux.scala 19:72:@1691.4]
  wire [31:0] _T_754; // @[Mux.scala 19:72:@1692.4]
  wire [31:0] _T_756; // @[Mux.scala 19:72:@1693.4]
  wire [31:0] _T_758; // @[Mux.scala 19:72:@1694.4]
  wire [31:0] _T_760; // @[Mux.scala 19:72:@1695.4]
  wire [31:0] _T_762; // @[Mux.scala 19:72:@1696.4]
  wire [31:0] _T_764; // @[Mux.scala 19:72:@1697.4]
  wire [31:0] _T_766; // @[Mux.scala 19:72:@1698.4]
  wire [31:0] _T_768; // @[Mux.scala 19:72:@1699.4]
  wire [31:0] _T_770; // @[Mux.scala 19:72:@1700.4]
  wire [31:0] _T_772; // @[Mux.scala 19:72:@1701.4]
  wire [31:0] _T_774; // @[Mux.scala 19:72:@1702.4]
  wire [31:0] _T_776; // @[Mux.scala 19:72:@1703.4]
  wire [31:0] _T_778; // @[Mux.scala 19:72:@1704.4]
  wire [31:0] _T_780; // @[Mux.scala 19:72:@1705.4]
  wire [31:0] _T_782; // @[Mux.scala 19:72:@1706.4]
  wire [31:0] _T_784; // @[Mux.scala 19:72:@1707.4]
  wire [31:0] _T_786; // @[Mux.scala 19:72:@1708.4]
  wire [31:0] _T_788; // @[Mux.scala 19:72:@1709.4]
  wire [31:0] _T_790; // @[Mux.scala 19:72:@1710.4]
  wire [31:0] _T_792; // @[Mux.scala 19:72:@1711.4]
  wire [31:0] _T_794; // @[Mux.scala 19:72:@1712.4]
  wire [31:0] _T_796; // @[Mux.scala 19:72:@1713.4]
  wire [31:0] _T_798; // @[Mux.scala 19:72:@1714.4]
  wire [31:0] _T_800; // @[Mux.scala 19:72:@1715.4]
  wire [31:0] _T_802; // @[Mux.scala 19:72:@1716.4]
  wire [31:0] _T_804; // @[Mux.scala 19:72:@1717.4]
  wire [31:0] _T_806; // @[Mux.scala 19:72:@1718.4]
  wire [31:0] _T_808; // @[Mux.scala 19:72:@1719.4]
  wire [31:0] _T_809; // @[Mux.scala 19:72:@1720.4]
  wire [31:0] _T_810; // @[Mux.scala 19:72:@1721.4]
  wire [31:0] _T_811; // @[Mux.scala 19:72:@1722.4]
  wire [31:0] _T_812; // @[Mux.scala 19:72:@1723.4]
  wire [31:0] _T_813; // @[Mux.scala 19:72:@1724.4]
  wire [31:0] _T_814; // @[Mux.scala 19:72:@1725.4]
  wire [31:0] _T_815; // @[Mux.scala 19:72:@1726.4]
  wire [31:0] _T_816; // @[Mux.scala 19:72:@1727.4]
  wire [31:0] _T_817; // @[Mux.scala 19:72:@1728.4]
  wire [31:0] _T_818; // @[Mux.scala 19:72:@1729.4]
  wire [31:0] _T_819; // @[Mux.scala 19:72:@1730.4]
  wire [31:0] _T_820; // @[Mux.scala 19:72:@1731.4]
  wire [31:0] _T_821; // @[Mux.scala 19:72:@1732.4]
  wire [31:0] _T_822; // @[Mux.scala 19:72:@1733.4]
  wire [31:0] _T_823; // @[Mux.scala 19:72:@1734.4]
  wire [31:0] _T_824; // @[Mux.scala 19:72:@1735.4]
  wire [31:0] _T_825; // @[Mux.scala 19:72:@1736.4]
  wire [31:0] _T_826; // @[Mux.scala 19:72:@1737.4]
  wire [31:0] _T_827; // @[Mux.scala 19:72:@1738.4]
  wire [31:0] _T_828; // @[Mux.scala 19:72:@1739.4]
  wire [31:0] _T_829; // @[Mux.scala 19:72:@1740.4]
  wire [31:0] _T_830; // @[Mux.scala 19:72:@1741.4]
  wire [31:0] _T_831; // @[Mux.scala 19:72:@1742.4]
  wire [31:0] _T_832; // @[Mux.scala 19:72:@1743.4]
  wire [31:0] _T_833; // @[Mux.scala 19:72:@1744.4]
  wire [31:0] _T_834; // @[Mux.scala 19:72:@1745.4]
  wire [31:0] _T_835; // @[Mux.scala 19:72:@1746.4]
  wire [31:0] _T_836; // @[Mux.scala 19:72:@1747.4]
  wire [31:0] _T_837; // @[Mux.scala 19:72:@1748.4]
  wire [31:0] _T_838; // @[Mux.scala 19:72:@1749.4]
  wire [31:0] _T_839; // @[Mux.scala 19:72:@1750.4]
  wire [31:0] _T_840; // @[Mux.scala 19:72:@1751.4]
  wire [31:0] _T_841; // @[Mux.scala 19:72:@1752.4]
  wire [31:0] _T_842; // @[Mux.scala 19:72:@1753.4]
  wire [31:0] _T_843; // @[Mux.scala 19:72:@1754.4]
  wire [31:0] _T_844; // @[Mux.scala 19:72:@1755.4]
  wire [31:0] _T_845; // @[Mux.scala 19:72:@1756.4]
  wire [31:0] _T_846; // @[Mux.scala 19:72:@1757.4]
  wire [31:0] _T_847; // @[Mux.scala 19:72:@1758.4]
  wire [31:0] _T_848; // @[Mux.scala 19:72:@1759.4]
  wire [31:0] _T_849; // @[Mux.scala 19:72:@1760.4]
  wire [31:0] _T_850; // @[Mux.scala 19:72:@1761.4]
  wire [31:0] _T_851; // @[Mux.scala 19:72:@1762.4]
  wire [31:0] _T_852; // @[Mux.scala 19:72:@1763.4]
  wire [31:0] _T_853; // @[Mux.scala 19:72:@1764.4]
  wire [31:0] _T_854; // @[Mux.scala 19:72:@1765.4]
  wire [31:0] _T_855; // @[Mux.scala 19:72:@1766.4]
  wire [31:0] _T_856; // @[Mux.scala 19:72:@1767.4]
  wire [31:0] _T_857; // @[Mux.scala 19:72:@1768.4]
  wire [31:0] _T_858; // @[Mux.scala 19:72:@1769.4]
  wire [31:0] _T_859; // @[Mux.scala 19:72:@1770.4]
  wire [31:0] _T_860; // @[Mux.scala 19:72:@1771.4]
  wire [31:0] _T_861; // @[Mux.scala 19:72:@1772.4]
  wire [31:0] _T_862; // @[Mux.scala 19:72:@1773.4]
  wire [31:0] _T_863; // @[Mux.scala 19:72:@1774.4]
  wire [31:0] _T_864; // @[Mux.scala 19:72:@1775.4]
  wire [31:0] _T_865; // @[Mux.scala 19:72:@1776.4]
  wire [31:0] _T_866; // @[Mux.scala 19:72:@1777.4]
  wire [31:0] _T_867; // @[Mux.scala 19:72:@1778.4]
  wire [31:0] _T_868; // @[Mux.scala 19:72:@1779.4]
  wire [31:0] _T_869; // @[Mux.scala 19:72:@1780.4]
  wire [31:0] _T_870; // @[Mux.scala 19:72:@1781.4]
  wire [31:0] predict_0_jump_tgt; // @[Mux.scala 19:72:@1782.4]
  wire [1:0] _T_940; // @[Mux.scala 19:72:@1850.4]
  wire [1:0] _T_942; // @[Mux.scala 19:72:@1851.4]
  wire [1:0] _T_944; // @[Mux.scala 19:72:@1852.4]
  wire [1:0] _T_946; // @[Mux.scala 19:72:@1853.4]
  wire [1:0] _T_948; // @[Mux.scala 19:72:@1854.4]
  wire [1:0] _T_950; // @[Mux.scala 19:72:@1855.4]
  wire [1:0] _T_952; // @[Mux.scala 19:72:@1856.4]
  wire [1:0] _T_954; // @[Mux.scala 19:72:@1857.4]
  wire [1:0] _T_956; // @[Mux.scala 19:72:@1858.4]
  wire [1:0] _T_958; // @[Mux.scala 19:72:@1859.4]
  wire [1:0] _T_960; // @[Mux.scala 19:72:@1860.4]
  wire [1:0] _T_962; // @[Mux.scala 19:72:@1861.4]
  wire [1:0] _T_964; // @[Mux.scala 19:72:@1862.4]
  wire [1:0] _T_966; // @[Mux.scala 19:72:@1863.4]
  wire [1:0] _T_968; // @[Mux.scala 19:72:@1864.4]
  wire [1:0] _T_970; // @[Mux.scala 19:72:@1865.4]
  wire [1:0] _T_972; // @[Mux.scala 19:72:@1866.4]
  wire [1:0] _T_974; // @[Mux.scala 19:72:@1867.4]
  wire [1:0] _T_976; // @[Mux.scala 19:72:@1868.4]
  wire [1:0] _T_978; // @[Mux.scala 19:72:@1869.4]
  wire [1:0] _T_980; // @[Mux.scala 19:72:@1870.4]
  wire [1:0] _T_982; // @[Mux.scala 19:72:@1871.4]
  wire [1:0] _T_984; // @[Mux.scala 19:72:@1872.4]
  wire [1:0] _T_986; // @[Mux.scala 19:72:@1873.4]
  wire [1:0] _T_988; // @[Mux.scala 19:72:@1874.4]
  wire [1:0] _T_990; // @[Mux.scala 19:72:@1875.4]
  wire [1:0] _T_992; // @[Mux.scala 19:72:@1876.4]
  wire [1:0] _T_994; // @[Mux.scala 19:72:@1877.4]
  wire [1:0] _T_996; // @[Mux.scala 19:72:@1878.4]
  wire [1:0] _T_998; // @[Mux.scala 19:72:@1879.4]
  wire [1:0] _T_1000; // @[Mux.scala 19:72:@1880.4]
  wire [1:0] _T_1002; // @[Mux.scala 19:72:@1881.4]
  wire [1:0] _T_1004; // @[Mux.scala 19:72:@1882.4]
  wire [1:0] _T_1006; // @[Mux.scala 19:72:@1883.4]
  wire [1:0] _T_1008; // @[Mux.scala 19:72:@1884.4]
  wire [1:0] _T_1010; // @[Mux.scala 19:72:@1885.4]
  wire [1:0] _T_1012; // @[Mux.scala 19:72:@1886.4]
  wire [1:0] _T_1014; // @[Mux.scala 19:72:@1887.4]
  wire [1:0] _T_1016; // @[Mux.scala 19:72:@1888.4]
  wire [1:0] _T_1018; // @[Mux.scala 19:72:@1889.4]
  wire [1:0] _T_1020; // @[Mux.scala 19:72:@1890.4]
  wire [1:0] _T_1022; // @[Mux.scala 19:72:@1891.4]
  wire [1:0] _T_1024; // @[Mux.scala 19:72:@1892.4]
  wire [1:0] _T_1026; // @[Mux.scala 19:72:@1893.4]
  wire [1:0] _T_1028; // @[Mux.scala 19:72:@1894.4]
  wire [1:0] _T_1030; // @[Mux.scala 19:72:@1895.4]
  wire [1:0] _T_1032; // @[Mux.scala 19:72:@1896.4]
  wire [1:0] _T_1034; // @[Mux.scala 19:72:@1897.4]
  wire [1:0] _T_1036; // @[Mux.scala 19:72:@1898.4]
  wire [1:0] _T_1038; // @[Mux.scala 19:72:@1899.4]
  wire [1:0] _T_1040; // @[Mux.scala 19:72:@1900.4]
  wire [1:0] _T_1042; // @[Mux.scala 19:72:@1901.4]
  wire [1:0] _T_1044; // @[Mux.scala 19:72:@1902.4]
  wire [1:0] _T_1046; // @[Mux.scala 19:72:@1903.4]
  wire [1:0] _T_1048; // @[Mux.scala 19:72:@1904.4]
  wire [1:0] _T_1050; // @[Mux.scala 19:72:@1905.4]
  wire [1:0] _T_1052; // @[Mux.scala 19:72:@1906.4]
  wire [1:0] _T_1054; // @[Mux.scala 19:72:@1907.4]
  wire [1:0] _T_1056; // @[Mux.scala 19:72:@1908.4]
  wire [1:0] _T_1058; // @[Mux.scala 19:72:@1909.4]
  wire [1:0] _T_1060; // @[Mux.scala 19:72:@1910.4]
  wire [1:0] _T_1062; // @[Mux.scala 19:72:@1911.4]
  wire [1:0] _T_1064; // @[Mux.scala 19:72:@1912.4]
  wire [1:0] _T_1066; // @[Mux.scala 19:72:@1913.4]
  wire [1:0] _T_1067; // @[Mux.scala 19:72:@1914.4]
  wire [1:0] _T_1068; // @[Mux.scala 19:72:@1915.4]
  wire [1:0] _T_1069; // @[Mux.scala 19:72:@1916.4]
  wire [1:0] _T_1070; // @[Mux.scala 19:72:@1917.4]
  wire [1:0] _T_1071; // @[Mux.scala 19:72:@1918.4]
  wire [1:0] _T_1072; // @[Mux.scala 19:72:@1919.4]
  wire [1:0] _T_1073; // @[Mux.scala 19:72:@1920.4]
  wire [1:0] _T_1074; // @[Mux.scala 19:72:@1921.4]
  wire [1:0] _T_1075; // @[Mux.scala 19:72:@1922.4]
  wire [1:0] _T_1076; // @[Mux.scala 19:72:@1923.4]
  wire [1:0] _T_1077; // @[Mux.scala 19:72:@1924.4]
  wire [1:0] _T_1078; // @[Mux.scala 19:72:@1925.4]
  wire [1:0] _T_1079; // @[Mux.scala 19:72:@1926.4]
  wire [1:0] _T_1080; // @[Mux.scala 19:72:@1927.4]
  wire [1:0] _T_1081; // @[Mux.scala 19:72:@1928.4]
  wire [1:0] _T_1082; // @[Mux.scala 19:72:@1929.4]
  wire [1:0] _T_1083; // @[Mux.scala 19:72:@1930.4]
  wire [1:0] _T_1084; // @[Mux.scala 19:72:@1931.4]
  wire [1:0] _T_1085; // @[Mux.scala 19:72:@1932.4]
  wire [1:0] _T_1086; // @[Mux.scala 19:72:@1933.4]
  wire [1:0] _T_1087; // @[Mux.scala 19:72:@1934.4]
  wire [1:0] _T_1088; // @[Mux.scala 19:72:@1935.4]
  wire [1:0] _T_1089; // @[Mux.scala 19:72:@1936.4]
  wire [1:0] _T_1090; // @[Mux.scala 19:72:@1937.4]
  wire [1:0] _T_1091; // @[Mux.scala 19:72:@1938.4]
  wire [1:0] _T_1092; // @[Mux.scala 19:72:@1939.4]
  wire [1:0] _T_1093; // @[Mux.scala 19:72:@1940.4]
  wire [1:0] _T_1094; // @[Mux.scala 19:72:@1941.4]
  wire [1:0] _T_1095; // @[Mux.scala 19:72:@1942.4]
  wire [1:0] _T_1096; // @[Mux.scala 19:72:@1943.4]
  wire [1:0] _T_1097; // @[Mux.scala 19:72:@1944.4]
  wire [1:0] _T_1098; // @[Mux.scala 19:72:@1945.4]
  wire [1:0] _T_1099; // @[Mux.scala 19:72:@1946.4]
  wire [1:0] _T_1100; // @[Mux.scala 19:72:@1947.4]
  wire [1:0] _T_1101; // @[Mux.scala 19:72:@1948.4]
  wire [1:0] _T_1102; // @[Mux.scala 19:72:@1949.4]
  wire [1:0] _T_1103; // @[Mux.scala 19:72:@1950.4]
  wire [1:0] _T_1104; // @[Mux.scala 19:72:@1951.4]
  wire [1:0] _T_1105; // @[Mux.scala 19:72:@1952.4]
  wire [1:0] _T_1106; // @[Mux.scala 19:72:@1953.4]
  wire [1:0] _T_1107; // @[Mux.scala 19:72:@1954.4]
  wire [1:0] _T_1108; // @[Mux.scala 19:72:@1955.4]
  wire [1:0] _T_1109; // @[Mux.scala 19:72:@1956.4]
  wire [1:0] _T_1110; // @[Mux.scala 19:72:@1957.4]
  wire [1:0] _T_1111; // @[Mux.scala 19:72:@1958.4]
  wire [1:0] _T_1112; // @[Mux.scala 19:72:@1959.4]
  wire [1:0] _T_1113; // @[Mux.scala 19:72:@1960.4]
  wire [1:0] _T_1114; // @[Mux.scala 19:72:@1961.4]
  wire [1:0] _T_1115; // @[Mux.scala 19:72:@1962.4]
  wire [1:0] _T_1116; // @[Mux.scala 19:72:@1963.4]
  wire [1:0] _T_1117; // @[Mux.scala 19:72:@1964.4]
  wire [1:0] _T_1118; // @[Mux.scala 19:72:@1965.4]
  wire [1:0] _T_1119; // @[Mux.scala 19:72:@1966.4]
  wire [1:0] _T_1120; // @[Mux.scala 19:72:@1967.4]
  wire [1:0] _T_1121; // @[Mux.scala 19:72:@1968.4]
  wire [1:0] _T_1122; // @[Mux.scala 19:72:@1969.4]
  wire [1:0] _T_1123; // @[Mux.scala 19:72:@1970.4]
  wire [1:0] _T_1124; // @[Mux.scala 19:72:@1971.4]
  wire [1:0] _T_1125; // @[Mux.scala 19:72:@1972.4]
  wire [1:0] _T_1126; // @[Mux.scala 19:72:@1973.4]
  wire [1:0] _T_1127; // @[Mux.scala 19:72:@1974.4]
  wire [1:0] _T_1128; // @[Mux.scala 19:72:@1975.4]
  wire [1:0] predict_0_btype; // @[Mux.scala 19:72:@1976.4]
  wire [1:0] _T_1198; // @[Mux.scala 19:72:@2044.4]
  wire [1:0] _T_1200; // @[Mux.scala 19:72:@2045.4]
  wire [1:0] _T_1202; // @[Mux.scala 19:72:@2046.4]
  wire [1:0] _T_1204; // @[Mux.scala 19:72:@2047.4]
  wire [1:0] _T_1206; // @[Mux.scala 19:72:@2048.4]
  wire [1:0] _T_1208; // @[Mux.scala 19:72:@2049.4]
  wire [1:0] _T_1210; // @[Mux.scala 19:72:@2050.4]
  wire [1:0] _T_1212; // @[Mux.scala 19:72:@2051.4]
  wire [1:0] _T_1214; // @[Mux.scala 19:72:@2052.4]
  wire [1:0] _T_1216; // @[Mux.scala 19:72:@2053.4]
  wire [1:0] _T_1218; // @[Mux.scala 19:72:@2054.4]
  wire [1:0] _T_1220; // @[Mux.scala 19:72:@2055.4]
  wire [1:0] _T_1222; // @[Mux.scala 19:72:@2056.4]
  wire [1:0] _T_1224; // @[Mux.scala 19:72:@2057.4]
  wire [1:0] _T_1226; // @[Mux.scala 19:72:@2058.4]
  wire [1:0] _T_1228; // @[Mux.scala 19:72:@2059.4]
  wire [1:0] _T_1230; // @[Mux.scala 19:72:@2060.4]
  wire [1:0] _T_1232; // @[Mux.scala 19:72:@2061.4]
  wire [1:0] _T_1234; // @[Mux.scala 19:72:@2062.4]
  wire [1:0] _T_1236; // @[Mux.scala 19:72:@2063.4]
  wire [1:0] _T_1238; // @[Mux.scala 19:72:@2064.4]
  wire [1:0] _T_1240; // @[Mux.scala 19:72:@2065.4]
  wire [1:0] _T_1242; // @[Mux.scala 19:72:@2066.4]
  wire [1:0] _T_1244; // @[Mux.scala 19:72:@2067.4]
  wire [1:0] _T_1246; // @[Mux.scala 19:72:@2068.4]
  wire [1:0] _T_1248; // @[Mux.scala 19:72:@2069.4]
  wire [1:0] _T_1250; // @[Mux.scala 19:72:@2070.4]
  wire [1:0] _T_1252; // @[Mux.scala 19:72:@2071.4]
  wire [1:0] _T_1254; // @[Mux.scala 19:72:@2072.4]
  wire [1:0] _T_1256; // @[Mux.scala 19:72:@2073.4]
  wire [1:0] _T_1258; // @[Mux.scala 19:72:@2074.4]
  wire [1:0] _T_1260; // @[Mux.scala 19:72:@2075.4]
  wire [1:0] _T_1262; // @[Mux.scala 19:72:@2076.4]
  wire [1:0] _T_1264; // @[Mux.scala 19:72:@2077.4]
  wire [1:0] _T_1266; // @[Mux.scala 19:72:@2078.4]
  wire [1:0] _T_1268; // @[Mux.scala 19:72:@2079.4]
  wire [1:0] _T_1270; // @[Mux.scala 19:72:@2080.4]
  wire [1:0] _T_1272; // @[Mux.scala 19:72:@2081.4]
  wire [1:0] _T_1274; // @[Mux.scala 19:72:@2082.4]
  wire [1:0] _T_1276; // @[Mux.scala 19:72:@2083.4]
  wire [1:0] _T_1278; // @[Mux.scala 19:72:@2084.4]
  wire [1:0] _T_1280; // @[Mux.scala 19:72:@2085.4]
  wire [1:0] _T_1282; // @[Mux.scala 19:72:@2086.4]
  wire [1:0] _T_1284; // @[Mux.scala 19:72:@2087.4]
  wire [1:0] _T_1286; // @[Mux.scala 19:72:@2088.4]
  wire [1:0] _T_1288; // @[Mux.scala 19:72:@2089.4]
  wire [1:0] _T_1290; // @[Mux.scala 19:72:@2090.4]
  wire [1:0] _T_1292; // @[Mux.scala 19:72:@2091.4]
  wire [1:0] _T_1294; // @[Mux.scala 19:72:@2092.4]
  wire [1:0] _T_1296; // @[Mux.scala 19:72:@2093.4]
  wire [1:0] _T_1298; // @[Mux.scala 19:72:@2094.4]
  wire [1:0] _T_1300; // @[Mux.scala 19:72:@2095.4]
  wire [1:0] _T_1302; // @[Mux.scala 19:72:@2096.4]
  wire [1:0] _T_1304; // @[Mux.scala 19:72:@2097.4]
  wire [1:0] _T_1306; // @[Mux.scala 19:72:@2098.4]
  wire [1:0] _T_1308; // @[Mux.scala 19:72:@2099.4]
  wire [1:0] _T_1310; // @[Mux.scala 19:72:@2100.4]
  wire [1:0] _T_1312; // @[Mux.scala 19:72:@2101.4]
  wire [1:0] _T_1314; // @[Mux.scala 19:72:@2102.4]
  wire [1:0] _T_1316; // @[Mux.scala 19:72:@2103.4]
  wire [1:0] _T_1318; // @[Mux.scala 19:72:@2104.4]
  wire [1:0] _T_1320; // @[Mux.scala 19:72:@2105.4]
  wire [1:0] _T_1322; // @[Mux.scala 19:72:@2106.4]
  wire [1:0] _T_1324; // @[Mux.scala 19:72:@2107.4]
  wire [1:0] _T_1325; // @[Mux.scala 19:72:@2108.4]
  wire [1:0] _T_1326; // @[Mux.scala 19:72:@2109.4]
  wire [1:0] _T_1327; // @[Mux.scala 19:72:@2110.4]
  wire [1:0] _T_1328; // @[Mux.scala 19:72:@2111.4]
  wire [1:0] _T_1329; // @[Mux.scala 19:72:@2112.4]
  wire [1:0] _T_1330; // @[Mux.scala 19:72:@2113.4]
  wire [1:0] _T_1331; // @[Mux.scala 19:72:@2114.4]
  wire [1:0] _T_1332; // @[Mux.scala 19:72:@2115.4]
  wire [1:0] _T_1333; // @[Mux.scala 19:72:@2116.4]
  wire [1:0] _T_1334; // @[Mux.scala 19:72:@2117.4]
  wire [1:0] _T_1335; // @[Mux.scala 19:72:@2118.4]
  wire [1:0] _T_1336; // @[Mux.scala 19:72:@2119.4]
  wire [1:0] _T_1337; // @[Mux.scala 19:72:@2120.4]
  wire [1:0] _T_1338; // @[Mux.scala 19:72:@2121.4]
  wire [1:0] _T_1339; // @[Mux.scala 19:72:@2122.4]
  wire [1:0] _T_1340; // @[Mux.scala 19:72:@2123.4]
  wire [1:0] _T_1341; // @[Mux.scala 19:72:@2124.4]
  wire [1:0] _T_1342; // @[Mux.scala 19:72:@2125.4]
  wire [1:0] _T_1343; // @[Mux.scala 19:72:@2126.4]
  wire [1:0] _T_1344; // @[Mux.scala 19:72:@2127.4]
  wire [1:0] _T_1345; // @[Mux.scala 19:72:@2128.4]
  wire [1:0] _T_1346; // @[Mux.scala 19:72:@2129.4]
  wire [1:0] _T_1347; // @[Mux.scala 19:72:@2130.4]
  wire [1:0] _T_1348; // @[Mux.scala 19:72:@2131.4]
  wire [1:0] _T_1349; // @[Mux.scala 19:72:@2132.4]
  wire [1:0] _T_1350; // @[Mux.scala 19:72:@2133.4]
  wire [1:0] _T_1351; // @[Mux.scala 19:72:@2134.4]
  wire [1:0] _T_1352; // @[Mux.scala 19:72:@2135.4]
  wire [1:0] _T_1353; // @[Mux.scala 19:72:@2136.4]
  wire [1:0] _T_1354; // @[Mux.scala 19:72:@2137.4]
  wire [1:0] _T_1355; // @[Mux.scala 19:72:@2138.4]
  wire [1:0] _T_1356; // @[Mux.scala 19:72:@2139.4]
  wire [1:0] _T_1357; // @[Mux.scala 19:72:@2140.4]
  wire [1:0] _T_1358; // @[Mux.scala 19:72:@2141.4]
  wire [1:0] _T_1359; // @[Mux.scala 19:72:@2142.4]
  wire [1:0] _T_1360; // @[Mux.scala 19:72:@2143.4]
  wire [1:0] _T_1361; // @[Mux.scala 19:72:@2144.4]
  wire [1:0] _T_1362; // @[Mux.scala 19:72:@2145.4]
  wire [1:0] _T_1363; // @[Mux.scala 19:72:@2146.4]
  wire [1:0] _T_1364; // @[Mux.scala 19:72:@2147.4]
  wire [1:0] _T_1365; // @[Mux.scala 19:72:@2148.4]
  wire [1:0] _T_1366; // @[Mux.scala 19:72:@2149.4]
  wire [1:0] _T_1367; // @[Mux.scala 19:72:@2150.4]
  wire [1:0] _T_1368; // @[Mux.scala 19:72:@2151.4]
  wire [1:0] _T_1369; // @[Mux.scala 19:72:@2152.4]
  wire [1:0] _T_1370; // @[Mux.scala 19:72:@2153.4]
  wire [1:0] _T_1371; // @[Mux.scala 19:72:@2154.4]
  wire [1:0] _T_1372; // @[Mux.scala 19:72:@2155.4]
  wire [1:0] _T_1373; // @[Mux.scala 19:72:@2156.4]
  wire [1:0] _T_1374; // @[Mux.scala 19:72:@2157.4]
  wire [1:0] _T_1375; // @[Mux.scala 19:72:@2158.4]
  wire [1:0] _T_1376; // @[Mux.scala 19:72:@2159.4]
  wire [1:0] _T_1377; // @[Mux.scala 19:72:@2160.4]
  wire [1:0] _T_1378; // @[Mux.scala 19:72:@2161.4]
  wire [1:0] _T_1379; // @[Mux.scala 19:72:@2162.4]
  wire [1:0] _T_1380; // @[Mux.scala 19:72:@2163.4]
  wire [1:0] _T_1381; // @[Mux.scala 19:72:@2164.4]
  wire [1:0] _T_1382; // @[Mux.scala 19:72:@2165.4]
  wire [1:0] _T_1383; // @[Mux.scala 19:72:@2166.4]
  wire [1:0] _T_1384; // @[Mux.scala 19:72:@2167.4]
  wire [1:0] _T_1385; // @[Mux.scala 19:72:@2168.4]
  wire [1:0] _T_1386; // @[Mux.scala 19:72:@2169.4]
  wire [1:0] predict_0_hcount; // @[Mux.scala 19:72:@2170.4]
  wire  _T_1391; // @[BTB.scala 80:44:@2174.4]
  wire  _T_1393; // @[BTB.scala 69:34:@2175.4]
  wire  _T_1394; // @[BTB.scala 69:65:@2176.4]
  wire  _T_1396; // @[BTB.scala 69:58:@2177.4]
  wire  _T_1397; // @[BTB.scala 69:55:@2178.4]
  wire  _T_1399; // @[BTB.scala 69:26:@2179.4]
  wire  _T_1401; // @[BTB.scala 69:80:@2180.4]
  wire  _T_1402; // @[BTB.scala 69:70:@2181.4]
  wire [31:0] if_pc_1; // @[Cat.scala 30:58:@2187.4]
  wire [31:0] _T_1403; // @[BTB.scala 70:27:@2182.4]
  wire  _T_1410; // @[BTB.scala 76:47:@2189.4]
  wire  _T_1411; // @[BTB.scala 76:47:@2190.4]
  wire  _T_1412; // @[BTB.scala 76:47:@2191.4]
  wire  _T_1413; // @[BTB.scala 76:47:@2192.4]
  wire  _T_1414; // @[BTB.scala 76:47:@2193.4]
  wire  _T_1415; // @[BTB.scala 76:47:@2194.4]
  wire  _T_1416; // @[BTB.scala 76:47:@2195.4]
  wire  _T_1417; // @[BTB.scala 76:47:@2196.4]
  wire  _T_1418; // @[BTB.scala 76:47:@2197.4]
  wire  _T_1419; // @[BTB.scala 76:47:@2198.4]
  wire  _T_1420; // @[BTB.scala 76:47:@2199.4]
  wire  _T_1421; // @[BTB.scala 76:47:@2200.4]
  wire  _T_1422; // @[BTB.scala 76:47:@2201.4]
  wire  _T_1423; // @[BTB.scala 76:47:@2202.4]
  wire  _T_1424; // @[BTB.scala 76:47:@2203.4]
  wire  _T_1425; // @[BTB.scala 76:47:@2204.4]
  wire  _T_1426; // @[BTB.scala 76:47:@2205.4]
  wire  _T_1427; // @[BTB.scala 76:47:@2206.4]
  wire  _T_1428; // @[BTB.scala 76:47:@2207.4]
  wire  _T_1429; // @[BTB.scala 76:47:@2208.4]
  wire  _T_1430; // @[BTB.scala 76:47:@2209.4]
  wire  _T_1431; // @[BTB.scala 76:47:@2210.4]
  wire  _T_1432; // @[BTB.scala 76:47:@2211.4]
  wire  _T_1433; // @[BTB.scala 76:47:@2212.4]
  wire  _T_1434; // @[BTB.scala 76:47:@2213.4]
  wire  _T_1435; // @[BTB.scala 76:47:@2214.4]
  wire  _T_1436; // @[BTB.scala 76:47:@2215.4]
  wire  _T_1437; // @[BTB.scala 76:47:@2216.4]
  wire  _T_1438; // @[BTB.scala 76:47:@2217.4]
  wire  _T_1439; // @[BTB.scala 76:47:@2218.4]
  wire  _T_1440; // @[BTB.scala 76:47:@2219.4]
  wire  _T_1441; // @[BTB.scala 76:47:@2220.4]
  wire  _T_1442; // @[BTB.scala 76:47:@2221.4]
  wire  _T_1443; // @[BTB.scala 76:47:@2222.4]
  wire  _T_1444; // @[BTB.scala 76:47:@2223.4]
  wire  _T_1445; // @[BTB.scala 76:47:@2224.4]
  wire  _T_1446; // @[BTB.scala 76:47:@2225.4]
  wire  _T_1447; // @[BTB.scala 76:47:@2226.4]
  wire  _T_1448; // @[BTB.scala 76:47:@2227.4]
  wire  _T_1449; // @[BTB.scala 76:47:@2228.4]
  wire  _T_1450; // @[BTB.scala 76:47:@2229.4]
  wire  _T_1451; // @[BTB.scala 76:47:@2230.4]
  wire  _T_1452; // @[BTB.scala 76:47:@2231.4]
  wire  _T_1453; // @[BTB.scala 76:47:@2232.4]
  wire  _T_1454; // @[BTB.scala 76:47:@2233.4]
  wire  _T_1455; // @[BTB.scala 76:47:@2234.4]
  wire  _T_1456; // @[BTB.scala 76:47:@2235.4]
  wire  _T_1457; // @[BTB.scala 76:47:@2236.4]
  wire  _T_1458; // @[BTB.scala 76:47:@2237.4]
  wire  _T_1459; // @[BTB.scala 76:47:@2238.4]
  wire  _T_1460; // @[BTB.scala 76:47:@2239.4]
  wire  _T_1461; // @[BTB.scala 76:47:@2240.4]
  wire  _T_1462; // @[BTB.scala 76:47:@2241.4]
  wire  _T_1463; // @[BTB.scala 76:47:@2242.4]
  wire  _T_1464; // @[BTB.scala 76:47:@2243.4]
  wire  _T_1465; // @[BTB.scala 76:47:@2244.4]
  wire  _T_1466; // @[BTB.scala 76:47:@2245.4]
  wire  _T_1467; // @[BTB.scala 76:47:@2246.4]
  wire  _T_1468; // @[BTB.scala 76:47:@2247.4]
  wire  _T_1469; // @[BTB.scala 76:47:@2248.4]
  wire  _T_1470; // @[BTB.scala 76:47:@2249.4]
  wire  _T_1471; // @[BTB.scala 76:47:@2250.4]
  wire  _T_1472; // @[BTB.scala 76:47:@2251.4]
  wire  _T_1473; // @[BTB.scala 76:47:@2252.4]
  wire [7:0] _T_1550; // @[BTB.scala 76:62:@2324.4]
  wire [15:0] _T_1558; // @[BTB.scala 76:62:@2332.4]
  wire [7:0] _T_1565; // @[BTB.scala 76:62:@2339.4]
  wire [31:0] _T_1574; // @[BTB.scala 76:62:@2348.4]
  wire [7:0] _T_1581; // @[BTB.scala 76:62:@2355.4]
  wire [15:0] _T_1589; // @[BTB.scala 76:62:@2363.4]
  wire [7:0] _T_1596; // @[BTB.scala 76:62:@2370.4]
  wire [31:0] _T_1605; // @[BTB.scala 76:62:@2379.4]
  wire [63:0] _T_1606; // @[BTB.scala 76:62:@2380.4]
  wire [63:0] predict_1_lookup; // @[BTB.scala 76:69:@2573.4]
  wire  _T_1869; // @[Mux.scala 21:36:@2575.4]
  wire  _T_1870; // @[Mux.scala 21:36:@2576.4]
  wire  _T_1871; // @[Mux.scala 21:36:@2577.4]
  wire  _T_1872; // @[Mux.scala 21:36:@2578.4]
  wire  _T_1873; // @[Mux.scala 21:36:@2579.4]
  wire  _T_1874; // @[Mux.scala 21:36:@2580.4]
  wire  _T_1875; // @[Mux.scala 21:36:@2581.4]
  wire  _T_1876; // @[Mux.scala 21:36:@2582.4]
  wire  _T_1877; // @[Mux.scala 21:36:@2583.4]
  wire  _T_1878; // @[Mux.scala 21:36:@2584.4]
  wire  _T_1879; // @[Mux.scala 21:36:@2585.4]
  wire  _T_1880; // @[Mux.scala 21:36:@2586.4]
  wire  _T_1881; // @[Mux.scala 21:36:@2587.4]
  wire  _T_1882; // @[Mux.scala 21:36:@2588.4]
  wire  _T_1883; // @[Mux.scala 21:36:@2589.4]
  wire  _T_1884; // @[Mux.scala 21:36:@2590.4]
  wire  _T_1885; // @[Mux.scala 21:36:@2591.4]
  wire  _T_1886; // @[Mux.scala 21:36:@2592.4]
  wire  _T_1887; // @[Mux.scala 21:36:@2593.4]
  wire  _T_1888; // @[Mux.scala 21:36:@2594.4]
  wire  _T_1889; // @[Mux.scala 21:36:@2595.4]
  wire  _T_1890; // @[Mux.scala 21:36:@2596.4]
  wire  _T_1891; // @[Mux.scala 21:36:@2597.4]
  wire  _T_1892; // @[Mux.scala 21:36:@2598.4]
  wire  _T_1893; // @[Mux.scala 21:36:@2599.4]
  wire  _T_1894; // @[Mux.scala 21:36:@2600.4]
  wire  _T_1895; // @[Mux.scala 21:36:@2601.4]
  wire  _T_1896; // @[Mux.scala 21:36:@2602.4]
  wire  _T_1897; // @[Mux.scala 21:36:@2603.4]
  wire  _T_1898; // @[Mux.scala 21:36:@2604.4]
  wire  _T_1899; // @[Mux.scala 21:36:@2605.4]
  wire  _T_1900; // @[Mux.scala 21:36:@2606.4]
  wire  _T_1901; // @[Mux.scala 21:36:@2607.4]
  wire  _T_1902; // @[Mux.scala 21:36:@2608.4]
  wire  _T_1903; // @[Mux.scala 21:36:@2609.4]
  wire  _T_1904; // @[Mux.scala 21:36:@2610.4]
  wire  _T_1905; // @[Mux.scala 21:36:@2611.4]
  wire  _T_1906; // @[Mux.scala 21:36:@2612.4]
  wire  _T_1907; // @[Mux.scala 21:36:@2613.4]
  wire  _T_1908; // @[Mux.scala 21:36:@2614.4]
  wire  _T_1909; // @[Mux.scala 21:36:@2615.4]
  wire  _T_1910; // @[Mux.scala 21:36:@2616.4]
  wire  _T_1911; // @[Mux.scala 21:36:@2617.4]
  wire  _T_1912; // @[Mux.scala 21:36:@2618.4]
  wire  _T_1913; // @[Mux.scala 21:36:@2619.4]
  wire  _T_1914; // @[Mux.scala 21:36:@2620.4]
  wire  _T_1915; // @[Mux.scala 21:36:@2621.4]
  wire  _T_1916; // @[Mux.scala 21:36:@2622.4]
  wire  _T_1917; // @[Mux.scala 21:36:@2623.4]
  wire  _T_1918; // @[Mux.scala 21:36:@2624.4]
  wire  _T_1919; // @[Mux.scala 21:36:@2625.4]
  wire  _T_1920; // @[Mux.scala 21:36:@2626.4]
  wire  _T_1921; // @[Mux.scala 21:36:@2627.4]
  wire  _T_1922; // @[Mux.scala 21:36:@2628.4]
  wire  _T_1923; // @[Mux.scala 21:36:@2629.4]
  wire  _T_1924; // @[Mux.scala 21:36:@2630.4]
  wire  _T_1925; // @[Mux.scala 21:36:@2631.4]
  wire  _T_1926; // @[Mux.scala 21:36:@2632.4]
  wire  _T_1927; // @[Mux.scala 21:36:@2633.4]
  wire  _T_1928; // @[Mux.scala 21:36:@2634.4]
  wire  _T_1929; // @[Mux.scala 21:36:@2635.4]
  wire  _T_1930; // @[Mux.scala 21:36:@2636.4]
  wire  _T_1931; // @[Mux.scala 21:36:@2637.4]
  wire  _T_1932; // @[Mux.scala 21:36:@2638.4]
  wire [31:0] _T_1935; // @[Mux.scala 19:72:@2639.4]
  wire [31:0] _T_1937; // @[Mux.scala 19:72:@2640.4]
  wire [31:0] _T_1939; // @[Mux.scala 19:72:@2641.4]
  wire [31:0] _T_1941; // @[Mux.scala 19:72:@2642.4]
  wire [31:0] _T_1943; // @[Mux.scala 19:72:@2643.4]
  wire [31:0] _T_1945; // @[Mux.scala 19:72:@2644.4]
  wire [31:0] _T_1947; // @[Mux.scala 19:72:@2645.4]
  wire [31:0] _T_1949; // @[Mux.scala 19:72:@2646.4]
  wire [31:0] _T_1951; // @[Mux.scala 19:72:@2647.4]
  wire [31:0] _T_1953; // @[Mux.scala 19:72:@2648.4]
  wire [31:0] _T_1955; // @[Mux.scala 19:72:@2649.4]
  wire [31:0] _T_1957; // @[Mux.scala 19:72:@2650.4]
  wire [31:0] _T_1959; // @[Mux.scala 19:72:@2651.4]
  wire [31:0] _T_1961; // @[Mux.scala 19:72:@2652.4]
  wire [31:0] _T_1963; // @[Mux.scala 19:72:@2653.4]
  wire [31:0] _T_1965; // @[Mux.scala 19:72:@2654.4]
  wire [31:0] _T_1967; // @[Mux.scala 19:72:@2655.4]
  wire [31:0] _T_1969; // @[Mux.scala 19:72:@2656.4]
  wire [31:0] _T_1971; // @[Mux.scala 19:72:@2657.4]
  wire [31:0] _T_1973; // @[Mux.scala 19:72:@2658.4]
  wire [31:0] _T_1975; // @[Mux.scala 19:72:@2659.4]
  wire [31:0] _T_1977; // @[Mux.scala 19:72:@2660.4]
  wire [31:0] _T_1979; // @[Mux.scala 19:72:@2661.4]
  wire [31:0] _T_1981; // @[Mux.scala 19:72:@2662.4]
  wire [31:0] _T_1983; // @[Mux.scala 19:72:@2663.4]
  wire [31:0] _T_1985; // @[Mux.scala 19:72:@2664.4]
  wire [31:0] _T_1987; // @[Mux.scala 19:72:@2665.4]
  wire [31:0] _T_1989; // @[Mux.scala 19:72:@2666.4]
  wire [31:0] _T_1991; // @[Mux.scala 19:72:@2667.4]
  wire [31:0] _T_1993; // @[Mux.scala 19:72:@2668.4]
  wire [31:0] _T_1995; // @[Mux.scala 19:72:@2669.4]
  wire [31:0] _T_1997; // @[Mux.scala 19:72:@2670.4]
  wire [31:0] _T_1999; // @[Mux.scala 19:72:@2671.4]
  wire [31:0] _T_2001; // @[Mux.scala 19:72:@2672.4]
  wire [31:0] _T_2003; // @[Mux.scala 19:72:@2673.4]
  wire [31:0] _T_2005; // @[Mux.scala 19:72:@2674.4]
  wire [31:0] _T_2007; // @[Mux.scala 19:72:@2675.4]
  wire [31:0] _T_2009; // @[Mux.scala 19:72:@2676.4]
  wire [31:0] _T_2011; // @[Mux.scala 19:72:@2677.4]
  wire [31:0] _T_2013; // @[Mux.scala 19:72:@2678.4]
  wire [31:0] _T_2015; // @[Mux.scala 19:72:@2679.4]
  wire [31:0] _T_2017; // @[Mux.scala 19:72:@2680.4]
  wire [31:0] _T_2019; // @[Mux.scala 19:72:@2681.4]
  wire [31:0] _T_2021; // @[Mux.scala 19:72:@2682.4]
  wire [31:0] _T_2023; // @[Mux.scala 19:72:@2683.4]
  wire [31:0] _T_2025; // @[Mux.scala 19:72:@2684.4]
  wire [31:0] _T_2027; // @[Mux.scala 19:72:@2685.4]
  wire [31:0] _T_2029; // @[Mux.scala 19:72:@2686.4]
  wire [31:0] _T_2031; // @[Mux.scala 19:72:@2687.4]
  wire [31:0] _T_2033; // @[Mux.scala 19:72:@2688.4]
  wire [31:0] _T_2035; // @[Mux.scala 19:72:@2689.4]
  wire [31:0] _T_2037; // @[Mux.scala 19:72:@2690.4]
  wire [31:0] _T_2039; // @[Mux.scala 19:72:@2691.4]
  wire [31:0] _T_2041; // @[Mux.scala 19:72:@2692.4]
  wire [31:0] _T_2043; // @[Mux.scala 19:72:@2693.4]
  wire [31:0] _T_2045; // @[Mux.scala 19:72:@2694.4]
  wire [31:0] _T_2047; // @[Mux.scala 19:72:@2695.4]
  wire [31:0] _T_2049; // @[Mux.scala 19:72:@2696.4]
  wire [31:0] _T_2051; // @[Mux.scala 19:72:@2697.4]
  wire [31:0] _T_2053; // @[Mux.scala 19:72:@2698.4]
  wire [31:0] _T_2055; // @[Mux.scala 19:72:@2699.4]
  wire [31:0] _T_2057; // @[Mux.scala 19:72:@2700.4]
  wire [31:0] _T_2059; // @[Mux.scala 19:72:@2701.4]
  wire [31:0] _T_2061; // @[Mux.scala 19:72:@2702.4]
  wire [31:0] _T_2062; // @[Mux.scala 19:72:@2703.4]
  wire [31:0] _T_2063; // @[Mux.scala 19:72:@2704.4]
  wire [31:0] _T_2064; // @[Mux.scala 19:72:@2705.4]
  wire [31:0] _T_2065; // @[Mux.scala 19:72:@2706.4]
  wire [31:0] _T_2066; // @[Mux.scala 19:72:@2707.4]
  wire [31:0] _T_2067; // @[Mux.scala 19:72:@2708.4]
  wire [31:0] _T_2068; // @[Mux.scala 19:72:@2709.4]
  wire [31:0] _T_2069; // @[Mux.scala 19:72:@2710.4]
  wire [31:0] _T_2070; // @[Mux.scala 19:72:@2711.4]
  wire [31:0] _T_2071; // @[Mux.scala 19:72:@2712.4]
  wire [31:0] _T_2072; // @[Mux.scala 19:72:@2713.4]
  wire [31:0] _T_2073; // @[Mux.scala 19:72:@2714.4]
  wire [31:0] _T_2074; // @[Mux.scala 19:72:@2715.4]
  wire [31:0] _T_2075; // @[Mux.scala 19:72:@2716.4]
  wire [31:0] _T_2076; // @[Mux.scala 19:72:@2717.4]
  wire [31:0] _T_2077; // @[Mux.scala 19:72:@2718.4]
  wire [31:0] _T_2078; // @[Mux.scala 19:72:@2719.4]
  wire [31:0] _T_2079; // @[Mux.scala 19:72:@2720.4]
  wire [31:0] _T_2080; // @[Mux.scala 19:72:@2721.4]
  wire [31:0] _T_2081; // @[Mux.scala 19:72:@2722.4]
  wire [31:0] _T_2082; // @[Mux.scala 19:72:@2723.4]
  wire [31:0] _T_2083; // @[Mux.scala 19:72:@2724.4]
  wire [31:0] _T_2084; // @[Mux.scala 19:72:@2725.4]
  wire [31:0] _T_2085; // @[Mux.scala 19:72:@2726.4]
  wire [31:0] _T_2086; // @[Mux.scala 19:72:@2727.4]
  wire [31:0] _T_2087; // @[Mux.scala 19:72:@2728.4]
  wire [31:0] _T_2088; // @[Mux.scala 19:72:@2729.4]
  wire [31:0] _T_2089; // @[Mux.scala 19:72:@2730.4]
  wire [31:0] _T_2090; // @[Mux.scala 19:72:@2731.4]
  wire [31:0] _T_2091; // @[Mux.scala 19:72:@2732.4]
  wire [31:0] _T_2092; // @[Mux.scala 19:72:@2733.4]
  wire [31:0] _T_2093; // @[Mux.scala 19:72:@2734.4]
  wire [31:0] _T_2094; // @[Mux.scala 19:72:@2735.4]
  wire [31:0] _T_2095; // @[Mux.scala 19:72:@2736.4]
  wire [31:0] _T_2096; // @[Mux.scala 19:72:@2737.4]
  wire [31:0] _T_2097; // @[Mux.scala 19:72:@2738.4]
  wire [31:0] _T_2098; // @[Mux.scala 19:72:@2739.4]
  wire [31:0] _T_2099; // @[Mux.scala 19:72:@2740.4]
  wire [31:0] _T_2100; // @[Mux.scala 19:72:@2741.4]
  wire [31:0] _T_2101; // @[Mux.scala 19:72:@2742.4]
  wire [31:0] _T_2102; // @[Mux.scala 19:72:@2743.4]
  wire [31:0] _T_2103; // @[Mux.scala 19:72:@2744.4]
  wire [31:0] _T_2104; // @[Mux.scala 19:72:@2745.4]
  wire [31:0] _T_2105; // @[Mux.scala 19:72:@2746.4]
  wire [31:0] _T_2106; // @[Mux.scala 19:72:@2747.4]
  wire [31:0] _T_2107; // @[Mux.scala 19:72:@2748.4]
  wire [31:0] _T_2108; // @[Mux.scala 19:72:@2749.4]
  wire [31:0] _T_2109; // @[Mux.scala 19:72:@2750.4]
  wire [31:0] _T_2110; // @[Mux.scala 19:72:@2751.4]
  wire [31:0] _T_2111; // @[Mux.scala 19:72:@2752.4]
  wire [31:0] _T_2112; // @[Mux.scala 19:72:@2753.4]
  wire [31:0] _T_2113; // @[Mux.scala 19:72:@2754.4]
  wire [31:0] _T_2114; // @[Mux.scala 19:72:@2755.4]
  wire [31:0] _T_2115; // @[Mux.scala 19:72:@2756.4]
  wire [31:0] _T_2116; // @[Mux.scala 19:72:@2757.4]
  wire [31:0] _T_2117; // @[Mux.scala 19:72:@2758.4]
  wire [31:0] _T_2118; // @[Mux.scala 19:72:@2759.4]
  wire [31:0] _T_2119; // @[Mux.scala 19:72:@2760.4]
  wire [31:0] _T_2120; // @[Mux.scala 19:72:@2761.4]
  wire [31:0] _T_2121; // @[Mux.scala 19:72:@2762.4]
  wire [31:0] _T_2122; // @[Mux.scala 19:72:@2763.4]
  wire [31:0] _T_2123; // @[Mux.scala 19:72:@2764.4]
  wire [31:0] predict_1_jump_tgt; // @[Mux.scala 19:72:@2765.4]
  wire [1:0] _T_2193; // @[Mux.scala 19:72:@2833.4]
  wire [1:0] _T_2195; // @[Mux.scala 19:72:@2834.4]
  wire [1:0] _T_2197; // @[Mux.scala 19:72:@2835.4]
  wire [1:0] _T_2199; // @[Mux.scala 19:72:@2836.4]
  wire [1:0] _T_2201; // @[Mux.scala 19:72:@2837.4]
  wire [1:0] _T_2203; // @[Mux.scala 19:72:@2838.4]
  wire [1:0] _T_2205; // @[Mux.scala 19:72:@2839.4]
  wire [1:0] _T_2207; // @[Mux.scala 19:72:@2840.4]
  wire [1:0] _T_2209; // @[Mux.scala 19:72:@2841.4]
  wire [1:0] _T_2211; // @[Mux.scala 19:72:@2842.4]
  wire [1:0] _T_2213; // @[Mux.scala 19:72:@2843.4]
  wire [1:0] _T_2215; // @[Mux.scala 19:72:@2844.4]
  wire [1:0] _T_2217; // @[Mux.scala 19:72:@2845.4]
  wire [1:0] _T_2219; // @[Mux.scala 19:72:@2846.4]
  wire [1:0] _T_2221; // @[Mux.scala 19:72:@2847.4]
  wire [1:0] _T_2223; // @[Mux.scala 19:72:@2848.4]
  wire [1:0] _T_2225; // @[Mux.scala 19:72:@2849.4]
  wire [1:0] _T_2227; // @[Mux.scala 19:72:@2850.4]
  wire [1:0] _T_2229; // @[Mux.scala 19:72:@2851.4]
  wire [1:0] _T_2231; // @[Mux.scala 19:72:@2852.4]
  wire [1:0] _T_2233; // @[Mux.scala 19:72:@2853.4]
  wire [1:0] _T_2235; // @[Mux.scala 19:72:@2854.4]
  wire [1:0] _T_2237; // @[Mux.scala 19:72:@2855.4]
  wire [1:0] _T_2239; // @[Mux.scala 19:72:@2856.4]
  wire [1:0] _T_2241; // @[Mux.scala 19:72:@2857.4]
  wire [1:0] _T_2243; // @[Mux.scala 19:72:@2858.4]
  wire [1:0] _T_2245; // @[Mux.scala 19:72:@2859.4]
  wire [1:0] _T_2247; // @[Mux.scala 19:72:@2860.4]
  wire [1:0] _T_2249; // @[Mux.scala 19:72:@2861.4]
  wire [1:0] _T_2251; // @[Mux.scala 19:72:@2862.4]
  wire [1:0] _T_2253; // @[Mux.scala 19:72:@2863.4]
  wire [1:0] _T_2255; // @[Mux.scala 19:72:@2864.4]
  wire [1:0] _T_2257; // @[Mux.scala 19:72:@2865.4]
  wire [1:0] _T_2259; // @[Mux.scala 19:72:@2866.4]
  wire [1:0] _T_2261; // @[Mux.scala 19:72:@2867.4]
  wire [1:0] _T_2263; // @[Mux.scala 19:72:@2868.4]
  wire [1:0] _T_2265; // @[Mux.scala 19:72:@2869.4]
  wire [1:0] _T_2267; // @[Mux.scala 19:72:@2870.4]
  wire [1:0] _T_2269; // @[Mux.scala 19:72:@2871.4]
  wire [1:0] _T_2271; // @[Mux.scala 19:72:@2872.4]
  wire [1:0] _T_2273; // @[Mux.scala 19:72:@2873.4]
  wire [1:0] _T_2275; // @[Mux.scala 19:72:@2874.4]
  wire [1:0] _T_2277; // @[Mux.scala 19:72:@2875.4]
  wire [1:0] _T_2279; // @[Mux.scala 19:72:@2876.4]
  wire [1:0] _T_2281; // @[Mux.scala 19:72:@2877.4]
  wire [1:0] _T_2283; // @[Mux.scala 19:72:@2878.4]
  wire [1:0] _T_2285; // @[Mux.scala 19:72:@2879.4]
  wire [1:0] _T_2287; // @[Mux.scala 19:72:@2880.4]
  wire [1:0] _T_2289; // @[Mux.scala 19:72:@2881.4]
  wire [1:0] _T_2291; // @[Mux.scala 19:72:@2882.4]
  wire [1:0] _T_2293; // @[Mux.scala 19:72:@2883.4]
  wire [1:0] _T_2295; // @[Mux.scala 19:72:@2884.4]
  wire [1:0] _T_2297; // @[Mux.scala 19:72:@2885.4]
  wire [1:0] _T_2299; // @[Mux.scala 19:72:@2886.4]
  wire [1:0] _T_2301; // @[Mux.scala 19:72:@2887.4]
  wire [1:0] _T_2303; // @[Mux.scala 19:72:@2888.4]
  wire [1:0] _T_2305; // @[Mux.scala 19:72:@2889.4]
  wire [1:0] _T_2307; // @[Mux.scala 19:72:@2890.4]
  wire [1:0] _T_2309; // @[Mux.scala 19:72:@2891.4]
  wire [1:0] _T_2311; // @[Mux.scala 19:72:@2892.4]
  wire [1:0] _T_2313; // @[Mux.scala 19:72:@2893.4]
  wire [1:0] _T_2315; // @[Mux.scala 19:72:@2894.4]
  wire [1:0] _T_2317; // @[Mux.scala 19:72:@2895.4]
  wire [1:0] _T_2319; // @[Mux.scala 19:72:@2896.4]
  wire [1:0] _T_2320; // @[Mux.scala 19:72:@2897.4]
  wire [1:0] _T_2321; // @[Mux.scala 19:72:@2898.4]
  wire [1:0] _T_2322; // @[Mux.scala 19:72:@2899.4]
  wire [1:0] _T_2323; // @[Mux.scala 19:72:@2900.4]
  wire [1:0] _T_2324; // @[Mux.scala 19:72:@2901.4]
  wire [1:0] _T_2325; // @[Mux.scala 19:72:@2902.4]
  wire [1:0] _T_2326; // @[Mux.scala 19:72:@2903.4]
  wire [1:0] _T_2327; // @[Mux.scala 19:72:@2904.4]
  wire [1:0] _T_2328; // @[Mux.scala 19:72:@2905.4]
  wire [1:0] _T_2329; // @[Mux.scala 19:72:@2906.4]
  wire [1:0] _T_2330; // @[Mux.scala 19:72:@2907.4]
  wire [1:0] _T_2331; // @[Mux.scala 19:72:@2908.4]
  wire [1:0] _T_2332; // @[Mux.scala 19:72:@2909.4]
  wire [1:0] _T_2333; // @[Mux.scala 19:72:@2910.4]
  wire [1:0] _T_2334; // @[Mux.scala 19:72:@2911.4]
  wire [1:0] _T_2335; // @[Mux.scala 19:72:@2912.4]
  wire [1:0] _T_2336; // @[Mux.scala 19:72:@2913.4]
  wire [1:0] _T_2337; // @[Mux.scala 19:72:@2914.4]
  wire [1:0] _T_2338; // @[Mux.scala 19:72:@2915.4]
  wire [1:0] _T_2339; // @[Mux.scala 19:72:@2916.4]
  wire [1:0] _T_2340; // @[Mux.scala 19:72:@2917.4]
  wire [1:0] _T_2341; // @[Mux.scala 19:72:@2918.4]
  wire [1:0] _T_2342; // @[Mux.scala 19:72:@2919.4]
  wire [1:0] _T_2343; // @[Mux.scala 19:72:@2920.4]
  wire [1:0] _T_2344; // @[Mux.scala 19:72:@2921.4]
  wire [1:0] _T_2345; // @[Mux.scala 19:72:@2922.4]
  wire [1:0] _T_2346; // @[Mux.scala 19:72:@2923.4]
  wire [1:0] _T_2347; // @[Mux.scala 19:72:@2924.4]
  wire [1:0] _T_2348; // @[Mux.scala 19:72:@2925.4]
  wire [1:0] _T_2349; // @[Mux.scala 19:72:@2926.4]
  wire [1:0] _T_2350; // @[Mux.scala 19:72:@2927.4]
  wire [1:0] _T_2351; // @[Mux.scala 19:72:@2928.4]
  wire [1:0] _T_2352; // @[Mux.scala 19:72:@2929.4]
  wire [1:0] _T_2353; // @[Mux.scala 19:72:@2930.4]
  wire [1:0] _T_2354; // @[Mux.scala 19:72:@2931.4]
  wire [1:0] _T_2355; // @[Mux.scala 19:72:@2932.4]
  wire [1:0] _T_2356; // @[Mux.scala 19:72:@2933.4]
  wire [1:0] _T_2357; // @[Mux.scala 19:72:@2934.4]
  wire [1:0] _T_2358; // @[Mux.scala 19:72:@2935.4]
  wire [1:0] _T_2359; // @[Mux.scala 19:72:@2936.4]
  wire [1:0] _T_2360; // @[Mux.scala 19:72:@2937.4]
  wire [1:0] _T_2361; // @[Mux.scala 19:72:@2938.4]
  wire [1:0] _T_2362; // @[Mux.scala 19:72:@2939.4]
  wire [1:0] _T_2363; // @[Mux.scala 19:72:@2940.4]
  wire [1:0] _T_2364; // @[Mux.scala 19:72:@2941.4]
  wire [1:0] _T_2365; // @[Mux.scala 19:72:@2942.4]
  wire [1:0] _T_2366; // @[Mux.scala 19:72:@2943.4]
  wire [1:0] _T_2367; // @[Mux.scala 19:72:@2944.4]
  wire [1:0] _T_2368; // @[Mux.scala 19:72:@2945.4]
  wire [1:0] _T_2369; // @[Mux.scala 19:72:@2946.4]
  wire [1:0] _T_2370; // @[Mux.scala 19:72:@2947.4]
  wire [1:0] _T_2371; // @[Mux.scala 19:72:@2948.4]
  wire [1:0] _T_2372; // @[Mux.scala 19:72:@2949.4]
  wire [1:0] _T_2373; // @[Mux.scala 19:72:@2950.4]
  wire [1:0] _T_2374; // @[Mux.scala 19:72:@2951.4]
  wire [1:0] _T_2375; // @[Mux.scala 19:72:@2952.4]
  wire [1:0] _T_2376; // @[Mux.scala 19:72:@2953.4]
  wire [1:0] _T_2377; // @[Mux.scala 19:72:@2954.4]
  wire [1:0] _T_2378; // @[Mux.scala 19:72:@2955.4]
  wire [1:0] _T_2379; // @[Mux.scala 19:72:@2956.4]
  wire [1:0] _T_2380; // @[Mux.scala 19:72:@2957.4]
  wire [1:0] _T_2381; // @[Mux.scala 19:72:@2958.4]
  wire [1:0] predict_1_btype; // @[Mux.scala 19:72:@2959.4]
  wire [1:0] _T_2451; // @[Mux.scala 19:72:@3027.4]
  wire [1:0] _T_2453; // @[Mux.scala 19:72:@3028.4]
  wire [1:0] _T_2455; // @[Mux.scala 19:72:@3029.4]
  wire [1:0] _T_2457; // @[Mux.scala 19:72:@3030.4]
  wire [1:0] _T_2459; // @[Mux.scala 19:72:@3031.4]
  wire [1:0] _T_2461; // @[Mux.scala 19:72:@3032.4]
  wire [1:0] _T_2463; // @[Mux.scala 19:72:@3033.4]
  wire [1:0] _T_2465; // @[Mux.scala 19:72:@3034.4]
  wire [1:0] _T_2467; // @[Mux.scala 19:72:@3035.4]
  wire [1:0] _T_2469; // @[Mux.scala 19:72:@3036.4]
  wire [1:0] _T_2471; // @[Mux.scala 19:72:@3037.4]
  wire [1:0] _T_2473; // @[Mux.scala 19:72:@3038.4]
  wire [1:0] _T_2475; // @[Mux.scala 19:72:@3039.4]
  wire [1:0] _T_2477; // @[Mux.scala 19:72:@3040.4]
  wire [1:0] _T_2479; // @[Mux.scala 19:72:@3041.4]
  wire [1:0] _T_2481; // @[Mux.scala 19:72:@3042.4]
  wire [1:0] _T_2483; // @[Mux.scala 19:72:@3043.4]
  wire [1:0] _T_2485; // @[Mux.scala 19:72:@3044.4]
  wire [1:0] _T_2487; // @[Mux.scala 19:72:@3045.4]
  wire [1:0] _T_2489; // @[Mux.scala 19:72:@3046.4]
  wire [1:0] _T_2491; // @[Mux.scala 19:72:@3047.4]
  wire [1:0] _T_2493; // @[Mux.scala 19:72:@3048.4]
  wire [1:0] _T_2495; // @[Mux.scala 19:72:@3049.4]
  wire [1:0] _T_2497; // @[Mux.scala 19:72:@3050.4]
  wire [1:0] _T_2499; // @[Mux.scala 19:72:@3051.4]
  wire [1:0] _T_2501; // @[Mux.scala 19:72:@3052.4]
  wire [1:0] _T_2503; // @[Mux.scala 19:72:@3053.4]
  wire [1:0] _T_2505; // @[Mux.scala 19:72:@3054.4]
  wire [1:0] _T_2507; // @[Mux.scala 19:72:@3055.4]
  wire [1:0] _T_2509; // @[Mux.scala 19:72:@3056.4]
  wire [1:0] _T_2511; // @[Mux.scala 19:72:@3057.4]
  wire [1:0] _T_2513; // @[Mux.scala 19:72:@3058.4]
  wire [1:0] _T_2515; // @[Mux.scala 19:72:@3059.4]
  wire [1:0] _T_2517; // @[Mux.scala 19:72:@3060.4]
  wire [1:0] _T_2519; // @[Mux.scala 19:72:@3061.4]
  wire [1:0] _T_2521; // @[Mux.scala 19:72:@3062.4]
  wire [1:0] _T_2523; // @[Mux.scala 19:72:@3063.4]
  wire [1:0] _T_2525; // @[Mux.scala 19:72:@3064.4]
  wire [1:0] _T_2527; // @[Mux.scala 19:72:@3065.4]
  wire [1:0] _T_2529; // @[Mux.scala 19:72:@3066.4]
  wire [1:0] _T_2531; // @[Mux.scala 19:72:@3067.4]
  wire [1:0] _T_2533; // @[Mux.scala 19:72:@3068.4]
  wire [1:0] _T_2535; // @[Mux.scala 19:72:@3069.4]
  wire [1:0] _T_2537; // @[Mux.scala 19:72:@3070.4]
  wire [1:0] _T_2539; // @[Mux.scala 19:72:@3071.4]
  wire [1:0] _T_2541; // @[Mux.scala 19:72:@3072.4]
  wire [1:0] _T_2543; // @[Mux.scala 19:72:@3073.4]
  wire [1:0] _T_2545; // @[Mux.scala 19:72:@3074.4]
  wire [1:0] _T_2547; // @[Mux.scala 19:72:@3075.4]
  wire [1:0] _T_2549; // @[Mux.scala 19:72:@3076.4]
  wire [1:0] _T_2551; // @[Mux.scala 19:72:@3077.4]
  wire [1:0] _T_2553; // @[Mux.scala 19:72:@3078.4]
  wire [1:0] _T_2555; // @[Mux.scala 19:72:@3079.4]
  wire [1:0] _T_2557; // @[Mux.scala 19:72:@3080.4]
  wire [1:0] _T_2559; // @[Mux.scala 19:72:@3081.4]
  wire [1:0] _T_2561; // @[Mux.scala 19:72:@3082.4]
  wire [1:0] _T_2563; // @[Mux.scala 19:72:@3083.4]
  wire [1:0] _T_2565; // @[Mux.scala 19:72:@3084.4]
  wire [1:0] _T_2567; // @[Mux.scala 19:72:@3085.4]
  wire [1:0] _T_2569; // @[Mux.scala 19:72:@3086.4]
  wire [1:0] _T_2571; // @[Mux.scala 19:72:@3087.4]
  wire [1:0] _T_2573; // @[Mux.scala 19:72:@3088.4]
  wire [1:0] _T_2575; // @[Mux.scala 19:72:@3089.4]
  wire [1:0] _T_2577; // @[Mux.scala 19:72:@3090.4]
  wire [1:0] _T_2578; // @[Mux.scala 19:72:@3091.4]
  wire [1:0] _T_2579; // @[Mux.scala 19:72:@3092.4]
  wire [1:0] _T_2580; // @[Mux.scala 19:72:@3093.4]
  wire [1:0] _T_2581; // @[Mux.scala 19:72:@3094.4]
  wire [1:0] _T_2582; // @[Mux.scala 19:72:@3095.4]
  wire [1:0] _T_2583; // @[Mux.scala 19:72:@3096.4]
  wire [1:0] _T_2584; // @[Mux.scala 19:72:@3097.4]
  wire [1:0] _T_2585; // @[Mux.scala 19:72:@3098.4]
  wire [1:0] _T_2586; // @[Mux.scala 19:72:@3099.4]
  wire [1:0] _T_2587; // @[Mux.scala 19:72:@3100.4]
  wire [1:0] _T_2588; // @[Mux.scala 19:72:@3101.4]
  wire [1:0] _T_2589; // @[Mux.scala 19:72:@3102.4]
  wire [1:0] _T_2590; // @[Mux.scala 19:72:@3103.4]
  wire [1:0] _T_2591; // @[Mux.scala 19:72:@3104.4]
  wire [1:0] _T_2592; // @[Mux.scala 19:72:@3105.4]
  wire [1:0] _T_2593; // @[Mux.scala 19:72:@3106.4]
  wire [1:0] _T_2594; // @[Mux.scala 19:72:@3107.4]
  wire [1:0] _T_2595; // @[Mux.scala 19:72:@3108.4]
  wire [1:0] _T_2596; // @[Mux.scala 19:72:@3109.4]
  wire [1:0] _T_2597; // @[Mux.scala 19:72:@3110.4]
  wire [1:0] _T_2598; // @[Mux.scala 19:72:@3111.4]
  wire [1:0] _T_2599; // @[Mux.scala 19:72:@3112.4]
  wire [1:0] _T_2600; // @[Mux.scala 19:72:@3113.4]
  wire [1:0] _T_2601; // @[Mux.scala 19:72:@3114.4]
  wire [1:0] _T_2602; // @[Mux.scala 19:72:@3115.4]
  wire [1:0] _T_2603; // @[Mux.scala 19:72:@3116.4]
  wire [1:0] _T_2604; // @[Mux.scala 19:72:@3117.4]
  wire [1:0] _T_2605; // @[Mux.scala 19:72:@3118.4]
  wire [1:0] _T_2606; // @[Mux.scala 19:72:@3119.4]
  wire [1:0] _T_2607; // @[Mux.scala 19:72:@3120.4]
  wire [1:0] _T_2608; // @[Mux.scala 19:72:@3121.4]
  wire [1:0] _T_2609; // @[Mux.scala 19:72:@3122.4]
  wire [1:0] _T_2610; // @[Mux.scala 19:72:@3123.4]
  wire [1:0] _T_2611; // @[Mux.scala 19:72:@3124.4]
  wire [1:0] _T_2612; // @[Mux.scala 19:72:@3125.4]
  wire [1:0] _T_2613; // @[Mux.scala 19:72:@3126.4]
  wire [1:0] _T_2614; // @[Mux.scala 19:72:@3127.4]
  wire [1:0] _T_2615; // @[Mux.scala 19:72:@3128.4]
  wire [1:0] _T_2616; // @[Mux.scala 19:72:@3129.4]
  wire [1:0] _T_2617; // @[Mux.scala 19:72:@3130.4]
  wire [1:0] _T_2618; // @[Mux.scala 19:72:@3131.4]
  wire [1:0] _T_2619; // @[Mux.scala 19:72:@3132.4]
  wire [1:0] _T_2620; // @[Mux.scala 19:72:@3133.4]
  wire [1:0] _T_2621; // @[Mux.scala 19:72:@3134.4]
  wire [1:0] _T_2622; // @[Mux.scala 19:72:@3135.4]
  wire [1:0] _T_2623; // @[Mux.scala 19:72:@3136.4]
  wire [1:0] _T_2624; // @[Mux.scala 19:72:@3137.4]
  wire [1:0] _T_2625; // @[Mux.scala 19:72:@3138.4]
  wire [1:0] _T_2626; // @[Mux.scala 19:72:@3139.4]
  wire [1:0] _T_2627; // @[Mux.scala 19:72:@3140.4]
  wire [1:0] _T_2628; // @[Mux.scala 19:72:@3141.4]
  wire [1:0] _T_2629; // @[Mux.scala 19:72:@3142.4]
  wire [1:0] _T_2630; // @[Mux.scala 19:72:@3143.4]
  wire [1:0] _T_2631; // @[Mux.scala 19:72:@3144.4]
  wire [1:0] _T_2632; // @[Mux.scala 19:72:@3145.4]
  wire [1:0] _T_2633; // @[Mux.scala 19:72:@3146.4]
  wire [1:0] _T_2634; // @[Mux.scala 19:72:@3147.4]
  wire [1:0] _T_2635; // @[Mux.scala 19:72:@3148.4]
  wire [1:0] _T_2636; // @[Mux.scala 19:72:@3149.4]
  wire [1:0] _T_2637; // @[Mux.scala 19:72:@3150.4]
  wire [1:0] _T_2638; // @[Mux.scala 19:72:@3151.4]
  wire [1:0] _T_2639; // @[Mux.scala 19:72:@3152.4]
  wire [1:0] predict_1_hcount; // @[Mux.scala 19:72:@3153.4]
  wire  _T_2644; // @[BTB.scala 80:44:@3157.4]
  wire  _T_2646; // @[BTB.scala 69:34:@3158.4]
  wire  _T_2647; // @[BTB.scala 69:65:@3159.4]
  wire  _T_2649; // @[BTB.scala 69:58:@3160.4]
  wire  _T_2650; // @[BTB.scala 69:55:@3161.4]
  wire  _T_2652; // @[BTB.scala 69:26:@3162.4]
  wire  _T_2654; // @[BTB.scala 69:80:@3163.4]
  wire  _T_2655; // @[BTB.scala 69:70:@3164.4]
  wire [32:0] _T_2659; // @[BTB.scala 84:35:@3169.4]
  wire [31:0] predict_1_cont_tgt; // @[BTB.scala 84:35:@3170.4]
  wire [31:0] _T_2656; // @[BTB.scala 70:27:@3165.4]
  wire  _T_2672; // @[BTB.scala 85:47:@3179.4]
  wire  _T_2675; // @[BTB.scala 85:38:@3181.4]
  reg  fb_reg_valid; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_256;
  reg  fb_reg_redirect; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_257;
  reg [5:0] fb_reg_lfsr; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_258;
  reg [31:0] fb_reg_pc; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_259;
  reg [31:0] fb_reg_target; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_260;
  reg [1:0] fb_reg_btype; // @[BTB.scala 87:23:@3191.4]
  reg [31:0] _RAND_261;
  wire  _T_2683; // @[BTB.scala 99:36:@3197.4]
  wire  _T_2684; // @[BTB.scala 99:46:@3198.4]
  wire  _T_2685; // @[BTB.scala 99:40:@3199.4]
  wire [4:0] _T_2686; // @[BTB.scala 99:55:@3200.4]
  wire [5:0] _T_2687; // @[Cat.scala 30:58:@3201.4]
  wire  _T_2689; // @[BTB.scala 123:42:@3204.4]
  wire  _T_2690; // @[BTB.scala 123:42:@3205.4]
  wire  _T_2691; // @[BTB.scala 123:42:@3206.4]
  wire  _T_2692; // @[BTB.scala 123:42:@3207.4]
  wire  _T_2693; // @[BTB.scala 123:42:@3208.4]
  wire  _T_2694; // @[BTB.scala 123:42:@3209.4]
  wire  _T_2695; // @[BTB.scala 123:42:@3210.4]
  wire  _T_2696; // @[BTB.scala 123:42:@3211.4]
  wire  _T_2697; // @[BTB.scala 123:42:@3212.4]
  wire  _T_2698; // @[BTB.scala 123:42:@3213.4]
  wire  _T_2699; // @[BTB.scala 123:42:@3214.4]
  wire  _T_2700; // @[BTB.scala 123:42:@3215.4]
  wire  _T_2701; // @[BTB.scala 123:42:@3216.4]
  wire  _T_2702; // @[BTB.scala 123:42:@3217.4]
  wire  _T_2703; // @[BTB.scala 123:42:@3218.4]
  wire  _T_2704; // @[BTB.scala 123:42:@3219.4]
  wire  _T_2705; // @[BTB.scala 123:42:@3220.4]
  wire  _T_2706; // @[BTB.scala 123:42:@3221.4]
  wire  _T_2707; // @[BTB.scala 123:42:@3222.4]
  wire  _T_2708; // @[BTB.scala 123:42:@3223.4]
  wire  _T_2709; // @[BTB.scala 123:42:@3224.4]
  wire  _T_2710; // @[BTB.scala 123:42:@3225.4]
  wire  _T_2711; // @[BTB.scala 123:42:@3226.4]
  wire  _T_2712; // @[BTB.scala 123:42:@3227.4]
  wire  _T_2713; // @[BTB.scala 123:42:@3228.4]
  wire  _T_2714; // @[BTB.scala 123:42:@3229.4]
  wire  _T_2715; // @[BTB.scala 123:42:@3230.4]
  wire  _T_2716; // @[BTB.scala 123:42:@3231.4]
  wire  _T_2717; // @[BTB.scala 123:42:@3232.4]
  wire  _T_2718; // @[BTB.scala 123:42:@3233.4]
  wire  _T_2719; // @[BTB.scala 123:42:@3234.4]
  wire  _T_2720; // @[BTB.scala 123:42:@3235.4]
  wire  _T_2721; // @[BTB.scala 123:42:@3236.4]
  wire  _T_2722; // @[BTB.scala 123:42:@3237.4]
  wire  _T_2723; // @[BTB.scala 123:42:@3238.4]
  wire  _T_2724; // @[BTB.scala 123:42:@3239.4]
  wire  _T_2725; // @[BTB.scala 123:42:@3240.4]
  wire  _T_2726; // @[BTB.scala 123:42:@3241.4]
  wire  _T_2727; // @[BTB.scala 123:42:@3242.4]
  wire  _T_2728; // @[BTB.scala 123:42:@3243.4]
  wire  _T_2729; // @[BTB.scala 123:42:@3244.4]
  wire  _T_2730; // @[BTB.scala 123:42:@3245.4]
  wire  _T_2731; // @[BTB.scala 123:42:@3246.4]
  wire  _T_2732; // @[BTB.scala 123:42:@3247.4]
  wire  _T_2733; // @[BTB.scala 123:42:@3248.4]
  wire  _T_2734; // @[BTB.scala 123:42:@3249.4]
  wire  _T_2735; // @[BTB.scala 123:42:@3250.4]
  wire  _T_2736; // @[BTB.scala 123:42:@3251.4]
  wire  _T_2737; // @[BTB.scala 123:42:@3252.4]
  wire  _T_2738; // @[BTB.scala 123:42:@3253.4]
  wire  _T_2739; // @[BTB.scala 123:42:@3254.4]
  wire  _T_2740; // @[BTB.scala 123:42:@3255.4]
  wire  _T_2741; // @[BTB.scala 123:42:@3256.4]
  wire  _T_2742; // @[BTB.scala 123:42:@3257.4]
  wire  _T_2743; // @[BTB.scala 123:42:@3258.4]
  wire  _T_2744; // @[BTB.scala 123:42:@3259.4]
  wire  _T_2745; // @[BTB.scala 123:42:@3260.4]
  wire  _T_2746; // @[BTB.scala 123:42:@3261.4]
  wire  _T_2747; // @[BTB.scala 123:42:@3262.4]
  wire  _T_2748; // @[BTB.scala 123:42:@3263.4]
  wire  _T_2749; // @[BTB.scala 123:42:@3264.4]
  wire  _T_2750; // @[BTB.scala 123:42:@3265.4]
  wire  _T_2751; // @[BTB.scala 123:42:@3266.4]
  wire  _T_2752; // @[BTB.scala 123:42:@3267.4]
  wire [7:0] _T_2829; // @[BTB.scala 123:58:@3339.4]
  wire [15:0] _T_2837; // @[BTB.scala 123:58:@3347.4]
  wire [7:0] _T_2844; // @[BTB.scala 123:58:@3354.4]
  wire [31:0] _T_2853; // @[BTB.scala 123:58:@3363.4]
  wire [7:0] _T_2860; // @[BTB.scala 123:58:@3370.4]
  wire [15:0] _T_2868; // @[BTB.scala 123:58:@3378.4]
  wire [7:0] _T_2875; // @[BTB.scala 123:58:@3385.4]
  wire [31:0] _T_2884; // @[BTB.scala 123:58:@3394.4]
  wire [63:0] _T_2885; // @[BTB.scala 123:58:@3395.4]
  wire [63:0] fb_wire_lookup; // @[BTB.scala 123:65:@3588.4]
  wire  _T_3148; // @[Mux.scala 21:36:@3590.4]
  wire  _T_3149; // @[Mux.scala 21:36:@3591.4]
  wire  _T_3150; // @[Mux.scala 21:36:@3592.4]
  wire  _T_3151; // @[Mux.scala 21:36:@3593.4]
  wire  _T_3152; // @[Mux.scala 21:36:@3594.4]
  wire  _T_3153; // @[Mux.scala 21:36:@3595.4]
  wire  _T_3154; // @[Mux.scala 21:36:@3596.4]
  wire  _T_3155; // @[Mux.scala 21:36:@3597.4]
  wire  _T_3156; // @[Mux.scala 21:36:@3598.4]
  wire  _T_3157; // @[Mux.scala 21:36:@3599.4]
  wire  _T_3158; // @[Mux.scala 21:36:@3600.4]
  wire  _T_3159; // @[Mux.scala 21:36:@3601.4]
  wire  _T_3160; // @[Mux.scala 21:36:@3602.4]
  wire  _T_3161; // @[Mux.scala 21:36:@3603.4]
  wire  _T_3162; // @[Mux.scala 21:36:@3604.4]
  wire  _T_3163; // @[Mux.scala 21:36:@3605.4]
  wire  _T_3164; // @[Mux.scala 21:36:@3606.4]
  wire  _T_3165; // @[Mux.scala 21:36:@3607.4]
  wire  _T_3166; // @[Mux.scala 21:36:@3608.4]
  wire  _T_3167; // @[Mux.scala 21:36:@3609.4]
  wire  _T_3168; // @[Mux.scala 21:36:@3610.4]
  wire  _T_3169; // @[Mux.scala 21:36:@3611.4]
  wire  _T_3170; // @[Mux.scala 21:36:@3612.4]
  wire  _T_3171; // @[Mux.scala 21:36:@3613.4]
  wire  _T_3172; // @[Mux.scala 21:36:@3614.4]
  wire  _T_3173; // @[Mux.scala 21:36:@3615.4]
  wire  _T_3174; // @[Mux.scala 21:36:@3616.4]
  wire  _T_3175; // @[Mux.scala 21:36:@3617.4]
  wire  _T_3176; // @[Mux.scala 21:36:@3618.4]
  wire  _T_3177; // @[Mux.scala 21:36:@3619.4]
  wire  _T_3178; // @[Mux.scala 21:36:@3620.4]
  wire  _T_3179; // @[Mux.scala 21:36:@3621.4]
  wire  _T_3180; // @[Mux.scala 21:36:@3622.4]
  wire  _T_3181; // @[Mux.scala 21:36:@3623.4]
  wire  _T_3182; // @[Mux.scala 21:36:@3624.4]
  wire  _T_3183; // @[Mux.scala 21:36:@3625.4]
  wire  _T_3184; // @[Mux.scala 21:36:@3626.4]
  wire  _T_3185; // @[Mux.scala 21:36:@3627.4]
  wire  _T_3186; // @[Mux.scala 21:36:@3628.4]
  wire  _T_3187; // @[Mux.scala 21:36:@3629.4]
  wire  _T_3188; // @[Mux.scala 21:36:@3630.4]
  wire  _T_3189; // @[Mux.scala 21:36:@3631.4]
  wire  _T_3190; // @[Mux.scala 21:36:@3632.4]
  wire  _T_3191; // @[Mux.scala 21:36:@3633.4]
  wire  _T_3192; // @[Mux.scala 21:36:@3634.4]
  wire  _T_3193; // @[Mux.scala 21:36:@3635.4]
  wire  _T_3194; // @[Mux.scala 21:36:@3636.4]
  wire  _T_3195; // @[Mux.scala 21:36:@3637.4]
  wire  _T_3196; // @[Mux.scala 21:36:@3638.4]
  wire  _T_3197; // @[Mux.scala 21:36:@3639.4]
  wire  _T_3198; // @[Mux.scala 21:36:@3640.4]
  wire  _T_3199; // @[Mux.scala 21:36:@3641.4]
  wire  _T_3200; // @[Mux.scala 21:36:@3642.4]
  wire  _T_3201; // @[Mux.scala 21:36:@3643.4]
  wire  _T_3202; // @[Mux.scala 21:36:@3644.4]
  wire  _T_3203; // @[Mux.scala 21:36:@3645.4]
  wire  _T_3204; // @[Mux.scala 21:36:@3646.4]
  wire  _T_3205; // @[Mux.scala 21:36:@3647.4]
  wire  _T_3206; // @[Mux.scala 21:36:@3648.4]
  wire  _T_3207; // @[Mux.scala 21:36:@3649.4]
  wire  _T_3208; // @[Mux.scala 21:36:@3650.4]
  wire  _T_3209; // @[Mux.scala 21:36:@3651.4]
  wire  _T_3210; // @[Mux.scala 21:36:@3652.4]
  wire  _T_3211; // @[Mux.scala 21:36:@3653.4]
  wire [1:0] _T_3214; // @[Mux.scala 19:72:@3654.4]
  wire [1:0] _T_3216; // @[Mux.scala 19:72:@3655.4]
  wire [1:0] _T_3218; // @[Mux.scala 19:72:@3656.4]
  wire [1:0] _T_3220; // @[Mux.scala 19:72:@3657.4]
  wire [1:0] _T_3222; // @[Mux.scala 19:72:@3658.4]
  wire [1:0] _T_3224; // @[Mux.scala 19:72:@3659.4]
  wire [1:0] _T_3226; // @[Mux.scala 19:72:@3660.4]
  wire [1:0] _T_3228; // @[Mux.scala 19:72:@3661.4]
  wire [1:0] _T_3230; // @[Mux.scala 19:72:@3662.4]
  wire [1:0] _T_3232; // @[Mux.scala 19:72:@3663.4]
  wire [1:0] _T_3234; // @[Mux.scala 19:72:@3664.4]
  wire [1:0] _T_3236; // @[Mux.scala 19:72:@3665.4]
  wire [1:0] _T_3238; // @[Mux.scala 19:72:@3666.4]
  wire [1:0] _T_3240; // @[Mux.scala 19:72:@3667.4]
  wire [1:0] _T_3242; // @[Mux.scala 19:72:@3668.4]
  wire [1:0] _T_3244; // @[Mux.scala 19:72:@3669.4]
  wire [1:0] _T_3246; // @[Mux.scala 19:72:@3670.4]
  wire [1:0] _T_3248; // @[Mux.scala 19:72:@3671.4]
  wire [1:0] _T_3250; // @[Mux.scala 19:72:@3672.4]
  wire [1:0] _T_3252; // @[Mux.scala 19:72:@3673.4]
  wire [1:0] _T_3254; // @[Mux.scala 19:72:@3674.4]
  wire [1:0] _T_3256; // @[Mux.scala 19:72:@3675.4]
  wire [1:0] _T_3258; // @[Mux.scala 19:72:@3676.4]
  wire [1:0] _T_3260; // @[Mux.scala 19:72:@3677.4]
  wire [1:0] _T_3262; // @[Mux.scala 19:72:@3678.4]
  wire [1:0] _T_3264; // @[Mux.scala 19:72:@3679.4]
  wire [1:0] _T_3266; // @[Mux.scala 19:72:@3680.4]
  wire [1:0] _T_3268; // @[Mux.scala 19:72:@3681.4]
  wire [1:0] _T_3270; // @[Mux.scala 19:72:@3682.4]
  wire [1:0] _T_3272; // @[Mux.scala 19:72:@3683.4]
  wire [1:0] _T_3274; // @[Mux.scala 19:72:@3684.4]
  wire [1:0] _T_3276; // @[Mux.scala 19:72:@3685.4]
  wire [1:0] _T_3278; // @[Mux.scala 19:72:@3686.4]
  wire [1:0] _T_3280; // @[Mux.scala 19:72:@3687.4]
  wire [1:0] _T_3282; // @[Mux.scala 19:72:@3688.4]
  wire [1:0] _T_3284; // @[Mux.scala 19:72:@3689.4]
  wire [1:0] _T_3286; // @[Mux.scala 19:72:@3690.4]
  wire [1:0] _T_3288; // @[Mux.scala 19:72:@3691.4]
  wire [1:0] _T_3290; // @[Mux.scala 19:72:@3692.4]
  wire [1:0] _T_3292; // @[Mux.scala 19:72:@3693.4]
  wire [1:0] _T_3294; // @[Mux.scala 19:72:@3694.4]
  wire [1:0] _T_3296; // @[Mux.scala 19:72:@3695.4]
  wire [1:0] _T_3298; // @[Mux.scala 19:72:@3696.4]
  wire [1:0] _T_3300; // @[Mux.scala 19:72:@3697.4]
  wire [1:0] _T_3302; // @[Mux.scala 19:72:@3698.4]
  wire [1:0] _T_3304; // @[Mux.scala 19:72:@3699.4]
  wire [1:0] _T_3306; // @[Mux.scala 19:72:@3700.4]
  wire [1:0] _T_3308; // @[Mux.scala 19:72:@3701.4]
  wire [1:0] _T_3310; // @[Mux.scala 19:72:@3702.4]
  wire [1:0] _T_3312; // @[Mux.scala 19:72:@3703.4]
  wire [1:0] _T_3314; // @[Mux.scala 19:72:@3704.4]
  wire [1:0] _T_3316; // @[Mux.scala 19:72:@3705.4]
  wire [1:0] _T_3318; // @[Mux.scala 19:72:@3706.4]
  wire [1:0] _T_3320; // @[Mux.scala 19:72:@3707.4]
  wire [1:0] _T_3322; // @[Mux.scala 19:72:@3708.4]
  wire [1:0] _T_3324; // @[Mux.scala 19:72:@3709.4]
  wire [1:0] _T_3326; // @[Mux.scala 19:72:@3710.4]
  wire [1:0] _T_3328; // @[Mux.scala 19:72:@3711.4]
  wire [1:0] _T_3330; // @[Mux.scala 19:72:@3712.4]
  wire [1:0] _T_3332; // @[Mux.scala 19:72:@3713.4]
  wire [1:0] _T_3334; // @[Mux.scala 19:72:@3714.4]
  wire [1:0] _T_3336; // @[Mux.scala 19:72:@3715.4]
  wire [1:0] _T_3338; // @[Mux.scala 19:72:@3716.4]
  wire [1:0] _T_3340; // @[Mux.scala 19:72:@3717.4]
  wire [1:0] _T_3341; // @[Mux.scala 19:72:@3718.4]
  wire [1:0] _T_3342; // @[Mux.scala 19:72:@3719.4]
  wire [1:0] _T_3343; // @[Mux.scala 19:72:@3720.4]
  wire [1:0] _T_3344; // @[Mux.scala 19:72:@3721.4]
  wire [1:0] _T_3345; // @[Mux.scala 19:72:@3722.4]
  wire [1:0] _T_3346; // @[Mux.scala 19:72:@3723.4]
  wire [1:0] _T_3347; // @[Mux.scala 19:72:@3724.4]
  wire [1:0] _T_3348; // @[Mux.scala 19:72:@3725.4]
  wire [1:0] _T_3349; // @[Mux.scala 19:72:@3726.4]
  wire [1:0] _T_3350; // @[Mux.scala 19:72:@3727.4]
  wire [1:0] _T_3351; // @[Mux.scala 19:72:@3728.4]
  wire [1:0] _T_3352; // @[Mux.scala 19:72:@3729.4]
  wire [1:0] _T_3353; // @[Mux.scala 19:72:@3730.4]
  wire [1:0] _T_3354; // @[Mux.scala 19:72:@3731.4]
  wire [1:0] _T_3355; // @[Mux.scala 19:72:@3732.4]
  wire [1:0] _T_3356; // @[Mux.scala 19:72:@3733.4]
  wire [1:0] _T_3357; // @[Mux.scala 19:72:@3734.4]
  wire [1:0] _T_3358; // @[Mux.scala 19:72:@3735.4]
  wire [1:0] _T_3359; // @[Mux.scala 19:72:@3736.4]
  wire [1:0] _T_3360; // @[Mux.scala 19:72:@3737.4]
  wire [1:0] _T_3361; // @[Mux.scala 19:72:@3738.4]
  wire [1:0] _T_3362; // @[Mux.scala 19:72:@3739.4]
  wire [1:0] _T_3363; // @[Mux.scala 19:72:@3740.4]
  wire [1:0] _T_3364; // @[Mux.scala 19:72:@3741.4]
  wire [1:0] _T_3365; // @[Mux.scala 19:72:@3742.4]
  wire [1:0] _T_3366; // @[Mux.scala 19:72:@3743.4]
  wire [1:0] _T_3367; // @[Mux.scala 19:72:@3744.4]
  wire [1:0] _T_3368; // @[Mux.scala 19:72:@3745.4]
  wire [1:0] _T_3369; // @[Mux.scala 19:72:@3746.4]
  wire [1:0] _T_3370; // @[Mux.scala 19:72:@3747.4]
  wire [1:0] _T_3371; // @[Mux.scala 19:72:@3748.4]
  wire [1:0] _T_3372; // @[Mux.scala 19:72:@3749.4]
  wire [1:0] _T_3373; // @[Mux.scala 19:72:@3750.4]
  wire [1:0] _T_3374; // @[Mux.scala 19:72:@3751.4]
  wire [1:0] _T_3375; // @[Mux.scala 19:72:@3752.4]
  wire [1:0] _T_3376; // @[Mux.scala 19:72:@3753.4]
  wire [1:0] _T_3377; // @[Mux.scala 19:72:@3754.4]
  wire [1:0] _T_3378; // @[Mux.scala 19:72:@3755.4]
  wire [1:0] _T_3379; // @[Mux.scala 19:72:@3756.4]
  wire [1:0] _T_3380; // @[Mux.scala 19:72:@3757.4]
  wire [1:0] _T_3381; // @[Mux.scala 19:72:@3758.4]
  wire [1:0] _T_3382; // @[Mux.scala 19:72:@3759.4]
  wire [1:0] _T_3383; // @[Mux.scala 19:72:@3760.4]
  wire [1:0] _T_3384; // @[Mux.scala 19:72:@3761.4]
  wire [1:0] _T_3385; // @[Mux.scala 19:72:@3762.4]
  wire [1:0] _T_3386; // @[Mux.scala 19:72:@3763.4]
  wire [1:0] _T_3387; // @[Mux.scala 19:72:@3764.4]
  wire [1:0] _T_3388; // @[Mux.scala 19:72:@3765.4]
  wire [1:0] _T_3389; // @[Mux.scala 19:72:@3766.4]
  wire [1:0] _T_3390; // @[Mux.scala 19:72:@3767.4]
  wire [1:0] _T_3391; // @[Mux.scala 19:72:@3768.4]
  wire [1:0] _T_3392; // @[Mux.scala 19:72:@3769.4]
  wire [1:0] _T_3393; // @[Mux.scala 19:72:@3770.4]
  wire [1:0] _T_3394; // @[Mux.scala 19:72:@3771.4]
  wire [1:0] _T_3395; // @[Mux.scala 19:72:@3772.4]
  wire [1:0] _T_3396; // @[Mux.scala 19:72:@3773.4]
  wire [1:0] _T_3397; // @[Mux.scala 19:72:@3774.4]
  wire [1:0] _T_3398; // @[Mux.scala 19:72:@3775.4]
  wire [1:0] _T_3399; // @[Mux.scala 19:72:@3776.4]
  wire [1:0] _T_3400; // @[Mux.scala 19:72:@3777.4]
  wire [1:0] _T_3401; // @[Mux.scala 19:72:@3778.4]
  wire [1:0] _T_3402; // @[Mux.scala 19:72:@3779.4]
  wire [1:0] fb_wire_hcount; // @[Mux.scala 19:72:@3780.4]
  wire  _T_3407; // @[BTB.scala 121:30:@3784.4]
  wire [31:0] _T_3408; // @[OneHot.scala 26:18:@3785.4]
  wire [31:0] _T_3409; // @[OneHot.scala 27:18:@3786.4]
  wire  _T_3411; // @[OneHot.scala 28:14:@3787.4]
  wire [31:0] _T_3412; // @[OneHot.scala 28:28:@3788.4]
  wire [15:0] _T_3413; // @[OneHot.scala 26:18:@3789.4]
  wire [15:0] _T_3414; // @[OneHot.scala 27:18:@3790.4]
  wire  _T_3416; // @[OneHot.scala 28:14:@3791.4]
  wire [15:0] _T_3417; // @[OneHot.scala 28:28:@3792.4]
  wire [7:0] _T_3418; // @[OneHot.scala 26:18:@3793.4]
  wire [7:0] _T_3419; // @[OneHot.scala 27:18:@3794.4]
  wire  _T_3421; // @[OneHot.scala 28:14:@3795.4]
  wire [7:0] _T_3422; // @[OneHot.scala 28:28:@3796.4]
  wire [3:0] _T_3423; // @[OneHot.scala 26:18:@3797.4]
  wire [3:0] _T_3424; // @[OneHot.scala 27:18:@3798.4]
  wire  _T_3426; // @[OneHot.scala 28:14:@3799.4]
  wire [3:0] _T_3427; // @[OneHot.scala 28:28:@3800.4]
  wire [1:0] _T_3428; // @[OneHot.scala 26:18:@3801.4]
  wire [1:0] _T_3429; // @[OneHot.scala 27:18:@3802.4]
  wire  _T_3431; // @[OneHot.scala 28:14:@3803.4]
  wire [1:0] _T_3432; // @[OneHot.scala 28:28:@3804.4]
  wire  _T_3433; // @[CircuitMath.scala 30:8:@3805.4]
  wire [5:0] _T_3438; // @[Cat.scala 30:58:@3810.4]
  wire [63:0] _T_3700; // @[BTB.scala 127:21:@4003.4]
  wire  _T_3702; // @[BTB.scala 127:21:@4004.4]
  wire  _T_3965; // @[OneHot.scala 39:40:@4198.4]
  wire  _T_3966; // @[OneHot.scala 39:40:@4199.4]
  wire  _T_3967; // @[OneHot.scala 39:40:@4200.4]
  wire  _T_3968; // @[OneHot.scala 39:40:@4201.4]
  wire  _T_3969; // @[OneHot.scala 39:40:@4202.4]
  wire  _T_3970; // @[OneHot.scala 39:40:@4203.4]
  wire  _T_3971; // @[OneHot.scala 39:40:@4204.4]
  wire  _T_3972; // @[OneHot.scala 39:40:@4205.4]
  wire  _T_3973; // @[OneHot.scala 39:40:@4206.4]
  wire  _T_3974; // @[OneHot.scala 39:40:@4207.4]
  wire  _T_3975; // @[OneHot.scala 39:40:@4208.4]
  wire  _T_3976; // @[OneHot.scala 39:40:@4209.4]
  wire  _T_3977; // @[OneHot.scala 39:40:@4210.4]
  wire  _T_3978; // @[OneHot.scala 39:40:@4211.4]
  wire  _T_3979; // @[OneHot.scala 39:40:@4212.4]
  wire  _T_3980; // @[OneHot.scala 39:40:@4213.4]
  wire  _T_3981; // @[OneHot.scala 39:40:@4214.4]
  wire  _T_3982; // @[OneHot.scala 39:40:@4215.4]
  wire  _T_3983; // @[OneHot.scala 39:40:@4216.4]
  wire  _T_3984; // @[OneHot.scala 39:40:@4217.4]
  wire  _T_3985; // @[OneHot.scala 39:40:@4218.4]
  wire  _T_3986; // @[OneHot.scala 39:40:@4219.4]
  wire  _T_3987; // @[OneHot.scala 39:40:@4220.4]
  wire  _T_3988; // @[OneHot.scala 39:40:@4221.4]
  wire  _T_3989; // @[OneHot.scala 39:40:@4222.4]
  wire  _T_3990; // @[OneHot.scala 39:40:@4223.4]
  wire  _T_3991; // @[OneHot.scala 39:40:@4224.4]
  wire  _T_3992; // @[OneHot.scala 39:40:@4225.4]
  wire  _T_3993; // @[OneHot.scala 39:40:@4226.4]
  wire  _T_3994; // @[OneHot.scala 39:40:@4227.4]
  wire  _T_3995; // @[OneHot.scala 39:40:@4228.4]
  wire  _T_3996; // @[OneHot.scala 39:40:@4229.4]
  wire  _T_3997; // @[OneHot.scala 39:40:@4230.4]
  wire  _T_3998; // @[OneHot.scala 39:40:@4231.4]
  wire  _T_3999; // @[OneHot.scala 39:40:@4232.4]
  wire  _T_4000; // @[OneHot.scala 39:40:@4233.4]
  wire  _T_4001; // @[OneHot.scala 39:40:@4234.4]
  wire  _T_4002; // @[OneHot.scala 39:40:@4235.4]
  wire  _T_4003; // @[OneHot.scala 39:40:@4236.4]
  wire  _T_4004; // @[OneHot.scala 39:40:@4237.4]
  wire  _T_4005; // @[OneHot.scala 39:40:@4238.4]
  wire  _T_4006; // @[OneHot.scala 39:40:@4239.4]
  wire  _T_4007; // @[OneHot.scala 39:40:@4240.4]
  wire  _T_4008; // @[OneHot.scala 39:40:@4241.4]
  wire  _T_4009; // @[OneHot.scala 39:40:@4242.4]
  wire  _T_4010; // @[OneHot.scala 39:40:@4243.4]
  wire  _T_4011; // @[OneHot.scala 39:40:@4244.4]
  wire  _T_4012; // @[OneHot.scala 39:40:@4245.4]
  wire  _T_4013; // @[OneHot.scala 39:40:@4246.4]
  wire  _T_4014; // @[OneHot.scala 39:40:@4247.4]
  wire  _T_4015; // @[OneHot.scala 39:40:@4248.4]
  wire  _T_4016; // @[OneHot.scala 39:40:@4249.4]
  wire  _T_4017; // @[OneHot.scala 39:40:@4250.4]
  wire  _T_4018; // @[OneHot.scala 39:40:@4251.4]
  wire  _T_4019; // @[OneHot.scala 39:40:@4252.4]
  wire  _T_4020; // @[OneHot.scala 39:40:@4253.4]
  wire  _T_4021; // @[OneHot.scala 39:40:@4254.4]
  wire  _T_4022; // @[OneHot.scala 39:40:@4255.4]
  wire  _T_4023; // @[OneHot.scala 39:40:@4256.4]
  wire  _T_4024; // @[OneHot.scala 39:40:@4257.4]
  wire  _T_4025; // @[OneHot.scala 39:40:@4258.4]
  wire  _T_4026; // @[OneHot.scala 39:40:@4259.4]
  wire  _T_4027; // @[OneHot.scala 39:40:@4260.4]
  wire [5:0] _T_4093; // @[Mux.scala 31:69:@4262.4]
  wire [5:0] _T_4094; // @[Mux.scala 31:69:@4263.4]
  wire [5:0] _T_4095; // @[Mux.scala 31:69:@4264.4]
  wire [5:0] _T_4096; // @[Mux.scala 31:69:@4265.4]
  wire [5:0] _T_4097; // @[Mux.scala 31:69:@4266.4]
  wire [5:0] _T_4098; // @[Mux.scala 31:69:@4267.4]
  wire [5:0] _T_4099; // @[Mux.scala 31:69:@4268.4]
  wire [5:0] _T_4100; // @[Mux.scala 31:69:@4269.4]
  wire [5:0] _T_4101; // @[Mux.scala 31:69:@4270.4]
  wire [5:0] _T_4102; // @[Mux.scala 31:69:@4271.4]
  wire [5:0] _T_4103; // @[Mux.scala 31:69:@4272.4]
  wire [5:0] _T_4104; // @[Mux.scala 31:69:@4273.4]
  wire [5:0] _T_4105; // @[Mux.scala 31:69:@4274.4]
  wire [5:0] _T_4106; // @[Mux.scala 31:69:@4275.4]
  wire [5:0] _T_4107; // @[Mux.scala 31:69:@4276.4]
  wire [5:0] _T_4108; // @[Mux.scala 31:69:@4277.4]
  wire [5:0] _T_4109; // @[Mux.scala 31:69:@4278.4]
  wire [5:0] _T_4110; // @[Mux.scala 31:69:@4279.4]
  wire [5:0] _T_4111; // @[Mux.scala 31:69:@4280.4]
  wire [5:0] _T_4112; // @[Mux.scala 31:69:@4281.4]
  wire [5:0] _T_4113; // @[Mux.scala 31:69:@4282.4]
  wire [5:0] _T_4114; // @[Mux.scala 31:69:@4283.4]
  wire [5:0] _T_4115; // @[Mux.scala 31:69:@4284.4]
  wire [5:0] _T_4116; // @[Mux.scala 31:69:@4285.4]
  wire [5:0] _T_4117; // @[Mux.scala 31:69:@4286.4]
  wire [5:0] _T_4118; // @[Mux.scala 31:69:@4287.4]
  wire [5:0] _T_4119; // @[Mux.scala 31:69:@4288.4]
  wire [5:0] _T_4120; // @[Mux.scala 31:69:@4289.4]
  wire [5:0] _T_4121; // @[Mux.scala 31:69:@4290.4]
  wire [5:0] _T_4122; // @[Mux.scala 31:69:@4291.4]
  wire [5:0] _T_4123; // @[Mux.scala 31:69:@4292.4]
  wire [5:0] _T_4124; // @[Mux.scala 31:69:@4293.4]
  wire [5:0] _T_4125; // @[Mux.scala 31:69:@4294.4]
  wire [5:0] _T_4126; // @[Mux.scala 31:69:@4295.4]
  wire [5:0] _T_4127; // @[Mux.scala 31:69:@4296.4]
  wire [5:0] _T_4128; // @[Mux.scala 31:69:@4297.4]
  wire [5:0] _T_4129; // @[Mux.scala 31:69:@4298.4]
  wire [5:0] _T_4130; // @[Mux.scala 31:69:@4299.4]
  wire [5:0] _T_4131; // @[Mux.scala 31:69:@4300.4]
  wire [5:0] _T_4132; // @[Mux.scala 31:69:@4301.4]
  wire [5:0] _T_4133; // @[Mux.scala 31:69:@4302.4]
  wire [5:0] _T_4134; // @[Mux.scala 31:69:@4303.4]
  wire [5:0] _T_4135; // @[Mux.scala 31:69:@4304.4]
  wire [5:0] _T_4136; // @[Mux.scala 31:69:@4305.4]
  wire [5:0] _T_4137; // @[Mux.scala 31:69:@4306.4]
  wire [5:0] _T_4138; // @[Mux.scala 31:69:@4307.4]
  wire [5:0] _T_4139; // @[Mux.scala 31:69:@4308.4]
  wire [5:0] _T_4140; // @[Mux.scala 31:69:@4309.4]
  wire [5:0] _T_4141; // @[Mux.scala 31:69:@4310.4]
  wire [5:0] _T_4142; // @[Mux.scala 31:69:@4311.4]
  wire [5:0] _T_4143; // @[Mux.scala 31:69:@4312.4]
  wire [5:0] _T_4144; // @[Mux.scala 31:69:@4313.4]
  wire [5:0] _T_4145; // @[Mux.scala 31:69:@4314.4]
  wire [5:0] _T_4146; // @[Mux.scala 31:69:@4315.4]
  wire [5:0] _T_4147; // @[Mux.scala 31:69:@4316.4]
  wire [5:0] _T_4148; // @[Mux.scala 31:69:@4317.4]
  wire [5:0] _T_4149; // @[Mux.scala 31:69:@4318.4]
  wire [5:0] _T_4150; // @[Mux.scala 31:69:@4319.4]
  wire [5:0] _T_4151; // @[Mux.scala 31:69:@4320.4]
  wire [5:0] _T_4152; // @[Mux.scala 31:69:@4321.4]
  wire [5:0] _T_4153; // @[Mux.scala 31:69:@4322.4]
  wire [5:0] _T_4154; // @[Mux.scala 31:69:@4323.4]
  wire [5:0] _T_4155; // @[Mux.scala 31:69:@4324.4]
  wire [5:0] _T_4156; // @[BTB.scala 127:10:@4325.4]
  wire [5:0] fb_wire_bindex; // @[BTB.scala 126:8:@4326.4]
  wire [31:0] _GEN_0; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_1; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_2; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_3; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_4; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_5; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_6; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_7; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_8; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_9; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_10; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_11; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_12; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_13; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_14; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_15; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_16; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_17; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_18; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_19; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_20; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_21; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_22; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_23; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_24; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_25; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_26; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_27; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_28; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_29; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_30; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_31; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_32; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_33; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_34; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_35; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_36; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_37; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_38; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_39; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_40; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_41; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_42; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_43; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_44; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_45; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_46; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_47; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_48; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_49; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_50; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_51; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_52; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_53; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_54; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_55; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_56; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_57; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_58; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_59; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_60; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_61; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_62; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_63; // @[BTB.scala 132:34:@4330.8]
  wire [31:0] _GEN_64; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_65; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_66; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_67; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_68; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_69; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_70; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_71; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_72; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_73; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_74; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_75; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_76; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_77; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_78; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_79; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_80; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_81; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_82; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_83; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_84; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_85; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_86; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_87; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_88; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_89; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_90; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_91; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_92; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_93; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_94; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_95; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_96; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_97; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_98; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_99; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_100; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_101; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_102; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_103; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_104; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_105; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_106; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_107; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_108; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_109; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_110; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_111; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_112; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_113; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_114; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_115; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_116; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_117; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_118; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_119; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_120; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_121; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_122; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_123; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_124; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_125; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_126; // @[BTB.scala 133:34:@4331.8]
  wire [31:0] _GEN_127; // @[BTB.scala 133:34:@4331.8]
  wire [1:0] _GEN_128; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_129; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_130; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_131; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_132; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_133; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_134; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_135; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_136; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_137; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_138; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_139; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_140; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_141; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_142; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_143; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_144; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_145; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_146; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_147; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_148; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_149; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_150; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_151; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_152; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_153; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_154; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_155; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_156; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_157; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_158; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_159; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_160; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_161; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_162; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_163; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_164; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_165; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_166; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_167; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_168; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_169; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_170; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_171; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_172; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_173; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_174; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_175; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_176; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_177; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_178; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_179; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_180; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_181; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_182; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_183; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_184; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_185; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_186; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_187; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_188; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_189; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_190; // @[BTB.scala 134:34:@4332.8]
  wire [1:0] _GEN_191; // @[BTB.scala 134:34:@4332.8]
  wire [31:0] _GEN_192; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_193; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_194; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_195; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_196; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_197; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_198; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_199; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_200; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_201; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_202; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_203; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_204; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_205; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_206; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_207; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_208; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_209; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_210; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_211; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_212; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_213; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_214; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_215; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_216; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_217; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_218; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_219; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_220; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_221; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_222; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_223; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_224; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_225; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_226; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_227; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_228; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_229; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_230; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_231; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_232; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_233; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_234; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_235; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_236; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_237; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_238; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_239; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_240; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_241; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_242; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_243; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_244; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_245; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_246; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_247; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_248; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_249; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_250; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_251; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_252; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_253; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_254; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_255; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_256; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_257; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_258; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_259; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_260; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_261; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_262; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_263; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_264; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_265; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_266; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_267; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_268; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_269; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_270; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_271; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_272; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_273; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_274; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_275; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_276; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_277; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_278; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_279; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_280; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_281; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_282; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_283; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_284; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_285; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_286; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_287; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_288; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_289; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_290; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_291; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_292; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_293; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_294; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_295; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_296; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_297; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_298; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_299; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_300; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_301; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_302; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_303; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_304; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_305; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_306; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_307; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_308; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_309; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_310; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_311; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_312; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_313; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_314; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_315; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_316; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_317; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_318; // @[BTB.scala 131:28:@4329.6]
  wire [31:0] _GEN_319; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_320; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_321; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_322; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_323; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_324; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_325; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_326; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_327; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_328; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_329; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_330; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_331; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_332; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_333; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_334; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_335; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_336; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_337; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_338; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_339; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_340; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_341; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_342; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_343; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_344; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_345; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_346; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_347; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_348; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_349; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_350; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_351; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_352; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_353; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_354; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_355; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_356; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_357; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_358; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_359; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_360; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_361; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_362; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_363; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_364; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_365; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_366; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_367; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_368; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_369; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_370; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_371; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_372; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_373; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_374; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_375; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_376; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_377; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_378; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_379; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_380; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_381; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_382; // @[BTB.scala 131:28:@4329.6]
  wire [1:0] _GEN_383; // @[BTB.scala 131:28:@4329.6]
  wire  _T_4159; // @[BTB.scala 136:24:@4334.6]
  wire  _T_4163; // @[BTB.scala 53:42:@4339.12]
  wire  _T_4164; // @[BTB.scala 53:49:@4340.12]
  wire  _T_4165; // @[BTB.scala 53:58:@4341.12]
  wire  _T_4167; // @[BTB.scala 53:56:@4342.12]
  wire  _T_4168; // @[BTB.scala 53:53:@4343.12]
  wire [1:0] _T_4169; // @[Cat.scala 30:58:@4344.12]
  wire [1:0] _GEN_384; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_385; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_386; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_387; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_388; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_389; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_390; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_391; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_392; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_393; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_394; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_395; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_396; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_397; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_398; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_399; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_400; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_401; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_402; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_403; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_404; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_405; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_406; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_407; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_408; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_409; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_410; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_411; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_412; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_413; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_414; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_415; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_416; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_417; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_418; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_419; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_420; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_421; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_422; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_423; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_424; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_425; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_426; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_427; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_428; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_429; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_430; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_431; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_432; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_433; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_434; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_435; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_436; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_437; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_438; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_439; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_440; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_441; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_442; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_443; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_444; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_445; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_446; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _GEN_447; // @[BTB.scala 139:38:@4345.12]
  wire [1:0] _T_4170; // @[BTB.scala 54:42:@4348.12]
  wire  _T_4172; // @[BTB.scala 54:42:@4349.12]
  wire  _T_4177; // @[BTB.scala 54:53:@4353.12]
  wire [1:0] _T_4178; // @[Cat.scala 30:58:@4354.12]
  wire [1:0] _GEN_448; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_449; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_450; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_451; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_452; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_453; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_454; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_455; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_456; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_457; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_458; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_459; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_460; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_461; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_462; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_463; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_464; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_465; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_466; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_467; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_468; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_469; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_470; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_471; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_472; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_473; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_474; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_475; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_476; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_477; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_478; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_479; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_480; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_481; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_482; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_483; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_484; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_485; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_486; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_487; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_488; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_489; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_490; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_491; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_492; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_493; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_494; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_495; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_496; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_497; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_498; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_499; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_500; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_501; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_502; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_503; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_504; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_505; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_506; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_507; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_508; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_509; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_510; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_511; // @[BTB.scala 141:38:@4355.12]
  wire [1:0] _GEN_512; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_513; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_514; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_515; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_516; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_517; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_518; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_519; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_520; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_521; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_522; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_523; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_524; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_525; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_526; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_527; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_528; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_529; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_530; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_531; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_532; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_533; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_534; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_535; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_536; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_537; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_538; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_539; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_540; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_541; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_542; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_543; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_544; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_545; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_546; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_547; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_548; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_549; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_550; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_551; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_552; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_553; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_554; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_555; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_556; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_557; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_558; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_559; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_560; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_561; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_562; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_563; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_564; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_565; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_566; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_567; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_568; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_569; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_570; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_571; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_572; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_573; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_574; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_575; // @[BTB.scala 138:32:@4338.10]
  wire [1:0] _GEN_576; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_577; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_578; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_579; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_580; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_581; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_582; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_583; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_584; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_585; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_586; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_587; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_588; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_589; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_590; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_591; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_592; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_593; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_594; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_595; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_596; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_597; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_598; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_599; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_600; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_601; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_602; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_603; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_604; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_605; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_606; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_607; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_608; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_609; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_610; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_611; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_612; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_613; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_614; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_615; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_616; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_617; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_618; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_619; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_620; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_621; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_622; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_623; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_624; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_625; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_626; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_627; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_628; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_629; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_630; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_631; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_632; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_633; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_634; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_635; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_636; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_637; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_638; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_639; // @[BTB.scala 144:36:@4360.12]
  wire [1:0] _GEN_640; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_641; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_642; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_643; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_644; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_645; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_646; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_647; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_648; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_649; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_650; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_651; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_652; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_653; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_654; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_655; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_656; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_657; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_658; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_659; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_660; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_661; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_662; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_663; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_664; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_665; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_666; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_667; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_668; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_669; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_670; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_671; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_672; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_673; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_674; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_675; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_676; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_677; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_678; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_679; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_680; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_681; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_682; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_683; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_684; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_685; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_686; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_687; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_688; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_689; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_690; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_691; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_692; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_693; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_694; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_695; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_696; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_697; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_698; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_699; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_700; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_701; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_702; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_703; // @[BTB.scala 143:35:@4359.10]
  wire [1:0] _GEN_704; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_705; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_706; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_707; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_708; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_709; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_710; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_711; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_712; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_713; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_714; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_715; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_716; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_717; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_718; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_719; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_720; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_721; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_722; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_723; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_724; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_725; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_726; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_727; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_728; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_729; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_730; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_731; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_732; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_733; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_734; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_735; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_736; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_737; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_738; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_739; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_740; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_741; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_742; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_743; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_744; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_745; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_746; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_747; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_748; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_749; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_750; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_751; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_752; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_753; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_754; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_755; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_756; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_757; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_758; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_759; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_760; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_761; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_762; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_763; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_764; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_765; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_766; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_767; // @[BTB.scala 137:28:@4337.8]
  wire [1:0] _GEN_768; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_769; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_770; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_771; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_772; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_773; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_774; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_775; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_776; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_777; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_778; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_779; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_780; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_781; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_782; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_783; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_784; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_785; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_786; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_787; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_788; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_789; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_790; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_791; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_792; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_793; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_794; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_795; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_796; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_797; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_798; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_799; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_800; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_801; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_802; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_803; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_804; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_805; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_806; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_807; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_808; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_809; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_810; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_811; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_812; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_813; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_814; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_815; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_816; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_817; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_818; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_819; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_820; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_821; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_822; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_823; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_824; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_825; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_826; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_827; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_828; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_829; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_830; // @[BTB.scala 136:46:@4335.6]
  wire [1:0] _GEN_831; // @[BTB.scala 136:46:@4335.6]
  wire [31:0] _GEN_832; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_833; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_834; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_835; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_836; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_837; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_838; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_839; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_840; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_841; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_842; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_843; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_844; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_845; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_846; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_847; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_848; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_849; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_850; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_851; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_852; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_853; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_854; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_855; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_856; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_857; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_858; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_859; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_860; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_861; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_862; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_863; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_864; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_865; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_866; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_867; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_868; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_869; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_870; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_871; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_872; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_873; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_874; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_875; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_876; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_877; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_878; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_879; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_880; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_881; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_882; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_883; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_884; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_885; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_886; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_887; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_888; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_889; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_890; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_891; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_892; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_893; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_894; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_895; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_896; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_897; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_898; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_899; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_900; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_901; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_902; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_903; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_904; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_905; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_906; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_907; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_908; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_909; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_910; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_911; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_912; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_913; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_914; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_915; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_916; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_917; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_918; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_919; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_920; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_921; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_922; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_923; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_924; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_925; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_926; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_927; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_928; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_929; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_930; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_931; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_932; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_933; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_934; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_935; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_936; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_937; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_938; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_939; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_940; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_941; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_942; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_943; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_944; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_945; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_946; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_947; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_948; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_949; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_950; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_951; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_952; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_953; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_954; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_955; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_956; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_957; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_958; // @[BTB.scala 130:23:@4328.4]
  wire [31:0] _GEN_959; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_960; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_961; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_962; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_963; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_964; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_965; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_966; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_967; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_968; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_969; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_970; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_971; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_972; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_973; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_974; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_975; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_976; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_977; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_978; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_979; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_980; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_981; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_982; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_983; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_984; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_985; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_986; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_987; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_988; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_989; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_990; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_991; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_992; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_993; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_994; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_995; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_996; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_997; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_998; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_999; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1000; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1001; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1002; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1003; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1004; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1005; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1006; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1007; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1008; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1009; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1010; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1011; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1012; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1013; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1014; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1015; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1016; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1017; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1018; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1019; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1020; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1021; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1022; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1023; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1024; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1025; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1026; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1027; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1028; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1029; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1030; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1031; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1032; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1033; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1034; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1035; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1036; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1037; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1038; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1039; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1040; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1041; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1042; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1043; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1044; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1045; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1046; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1047; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1048; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1049; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1050; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1051; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1052; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1053; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1054; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1055; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1056; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1057; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1058; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1059; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1060; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1061; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1062; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1063; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1064; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1065; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1066; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1067; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1068; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1069; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1070; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1071; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1072; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1073; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1074; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1075; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1076; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1077; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1078; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1079; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1080; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1081; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1082; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1083; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1084; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1085; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1086; // @[BTB.scala 130:23:@4328.4]
  wire [1:0] _GEN_1087; // @[BTB.scala 130:23:@4328.4]
  assign _T_152 = io_if_pc[31:3]; // @[FrontEnd.scala 9:13:@1202.4]
  assign if_pc_0 = {_T_152,1'h0,2'h0}; // @[Cat.scala 30:58:@1204.4]
  assign _T_157 = btb_pc_0 == if_pc_0; // @[BTB.scala 76:47:@1206.4]
  assign _T_158 = btb_pc_1 == if_pc_0; // @[BTB.scala 76:47:@1207.4]
  assign _T_159 = btb_pc_2 == if_pc_0; // @[BTB.scala 76:47:@1208.4]
  assign _T_160 = btb_pc_3 == if_pc_0; // @[BTB.scala 76:47:@1209.4]
  assign _T_161 = btb_pc_4 == if_pc_0; // @[BTB.scala 76:47:@1210.4]
  assign _T_162 = btb_pc_5 == if_pc_0; // @[BTB.scala 76:47:@1211.4]
  assign _T_163 = btb_pc_6 == if_pc_0; // @[BTB.scala 76:47:@1212.4]
  assign _T_164 = btb_pc_7 == if_pc_0; // @[BTB.scala 76:47:@1213.4]
  assign _T_165 = btb_pc_8 == if_pc_0; // @[BTB.scala 76:47:@1214.4]
  assign _T_166 = btb_pc_9 == if_pc_0; // @[BTB.scala 76:47:@1215.4]
  assign _T_167 = btb_pc_10 == if_pc_0; // @[BTB.scala 76:47:@1216.4]
  assign _T_168 = btb_pc_11 == if_pc_0; // @[BTB.scala 76:47:@1217.4]
  assign _T_169 = btb_pc_12 == if_pc_0; // @[BTB.scala 76:47:@1218.4]
  assign _T_170 = btb_pc_13 == if_pc_0; // @[BTB.scala 76:47:@1219.4]
  assign _T_171 = btb_pc_14 == if_pc_0; // @[BTB.scala 76:47:@1220.4]
  assign _T_172 = btb_pc_15 == if_pc_0; // @[BTB.scala 76:47:@1221.4]
  assign _T_173 = btb_pc_16 == if_pc_0; // @[BTB.scala 76:47:@1222.4]
  assign _T_174 = btb_pc_17 == if_pc_0; // @[BTB.scala 76:47:@1223.4]
  assign _T_175 = btb_pc_18 == if_pc_0; // @[BTB.scala 76:47:@1224.4]
  assign _T_176 = btb_pc_19 == if_pc_0; // @[BTB.scala 76:47:@1225.4]
  assign _T_177 = btb_pc_20 == if_pc_0; // @[BTB.scala 76:47:@1226.4]
  assign _T_178 = btb_pc_21 == if_pc_0; // @[BTB.scala 76:47:@1227.4]
  assign _T_179 = btb_pc_22 == if_pc_0; // @[BTB.scala 76:47:@1228.4]
  assign _T_180 = btb_pc_23 == if_pc_0; // @[BTB.scala 76:47:@1229.4]
  assign _T_181 = btb_pc_24 == if_pc_0; // @[BTB.scala 76:47:@1230.4]
  assign _T_182 = btb_pc_25 == if_pc_0; // @[BTB.scala 76:47:@1231.4]
  assign _T_183 = btb_pc_26 == if_pc_0; // @[BTB.scala 76:47:@1232.4]
  assign _T_184 = btb_pc_27 == if_pc_0; // @[BTB.scala 76:47:@1233.4]
  assign _T_185 = btb_pc_28 == if_pc_0; // @[BTB.scala 76:47:@1234.4]
  assign _T_186 = btb_pc_29 == if_pc_0; // @[BTB.scala 76:47:@1235.4]
  assign _T_187 = btb_pc_30 == if_pc_0; // @[BTB.scala 76:47:@1236.4]
  assign _T_188 = btb_pc_31 == if_pc_0; // @[BTB.scala 76:47:@1237.4]
  assign _T_189 = btb_pc_32 == if_pc_0; // @[BTB.scala 76:47:@1238.4]
  assign _T_190 = btb_pc_33 == if_pc_0; // @[BTB.scala 76:47:@1239.4]
  assign _T_191 = btb_pc_34 == if_pc_0; // @[BTB.scala 76:47:@1240.4]
  assign _T_192 = btb_pc_35 == if_pc_0; // @[BTB.scala 76:47:@1241.4]
  assign _T_193 = btb_pc_36 == if_pc_0; // @[BTB.scala 76:47:@1242.4]
  assign _T_194 = btb_pc_37 == if_pc_0; // @[BTB.scala 76:47:@1243.4]
  assign _T_195 = btb_pc_38 == if_pc_0; // @[BTB.scala 76:47:@1244.4]
  assign _T_196 = btb_pc_39 == if_pc_0; // @[BTB.scala 76:47:@1245.4]
  assign _T_197 = btb_pc_40 == if_pc_0; // @[BTB.scala 76:47:@1246.4]
  assign _T_198 = btb_pc_41 == if_pc_0; // @[BTB.scala 76:47:@1247.4]
  assign _T_199 = btb_pc_42 == if_pc_0; // @[BTB.scala 76:47:@1248.4]
  assign _T_200 = btb_pc_43 == if_pc_0; // @[BTB.scala 76:47:@1249.4]
  assign _T_201 = btb_pc_44 == if_pc_0; // @[BTB.scala 76:47:@1250.4]
  assign _T_202 = btb_pc_45 == if_pc_0; // @[BTB.scala 76:47:@1251.4]
  assign _T_203 = btb_pc_46 == if_pc_0; // @[BTB.scala 76:47:@1252.4]
  assign _T_204 = btb_pc_47 == if_pc_0; // @[BTB.scala 76:47:@1253.4]
  assign _T_205 = btb_pc_48 == if_pc_0; // @[BTB.scala 76:47:@1254.4]
  assign _T_206 = btb_pc_49 == if_pc_0; // @[BTB.scala 76:47:@1255.4]
  assign _T_207 = btb_pc_50 == if_pc_0; // @[BTB.scala 76:47:@1256.4]
  assign _T_208 = btb_pc_51 == if_pc_0; // @[BTB.scala 76:47:@1257.4]
  assign _T_209 = btb_pc_52 == if_pc_0; // @[BTB.scala 76:47:@1258.4]
  assign _T_210 = btb_pc_53 == if_pc_0; // @[BTB.scala 76:47:@1259.4]
  assign _T_211 = btb_pc_54 == if_pc_0; // @[BTB.scala 76:47:@1260.4]
  assign _T_212 = btb_pc_55 == if_pc_0; // @[BTB.scala 76:47:@1261.4]
  assign _T_213 = btb_pc_56 == if_pc_0; // @[BTB.scala 76:47:@1262.4]
  assign _T_214 = btb_pc_57 == if_pc_0; // @[BTB.scala 76:47:@1263.4]
  assign _T_215 = btb_pc_58 == if_pc_0; // @[BTB.scala 76:47:@1264.4]
  assign _T_216 = btb_pc_59 == if_pc_0; // @[BTB.scala 76:47:@1265.4]
  assign _T_217 = btb_pc_60 == if_pc_0; // @[BTB.scala 76:47:@1266.4]
  assign _T_218 = btb_pc_61 == if_pc_0; // @[BTB.scala 76:47:@1267.4]
  assign _T_219 = btb_pc_62 == if_pc_0; // @[BTB.scala 76:47:@1268.4]
  assign _T_220 = btb_pc_63 == if_pc_0; // @[BTB.scala 76:47:@1269.4]
  assign _T_297 = {_T_164,_T_163,_T_162,_T_161,_T_160,_T_159,_T_158,_T_157}; // @[BTB.scala 76:62:@1341.4]
  assign _T_305 = {_T_172,_T_171,_T_170,_T_169,_T_168,_T_167,_T_166,_T_165,_T_297}; // @[BTB.scala 76:62:@1349.4]
  assign _T_312 = {_T_180,_T_179,_T_178,_T_177,_T_176,_T_175,_T_174,_T_173}; // @[BTB.scala 76:62:@1356.4]
  assign _T_321 = {_T_188,_T_187,_T_186,_T_185,_T_184,_T_183,_T_182,_T_181,_T_312,_T_305}; // @[BTB.scala 76:62:@1365.4]
  assign _T_328 = {_T_196,_T_195,_T_194,_T_193,_T_192,_T_191,_T_190,_T_189}; // @[BTB.scala 76:62:@1372.4]
  assign _T_336 = {_T_204,_T_203,_T_202,_T_201,_T_200,_T_199,_T_198,_T_197,_T_328}; // @[BTB.scala 76:62:@1380.4]
  assign _T_343 = {_T_212,_T_211,_T_210,_T_209,_T_208,_T_207,_T_206,_T_205}; // @[BTB.scala 76:62:@1387.4]
  assign _T_352 = {_T_220,_T_219,_T_218,_T_217,_T_216,_T_215,_T_214,_T_213,_T_343,_T_336}; // @[BTB.scala 76:62:@1396.4]
  assign _T_353 = {_T_352,_T_321}; // @[BTB.scala 76:62:@1397.4]
  assign _T_355 = btb_btype_0 != 2'h0; // @[BTB.scala 52:66:@1398.4]
  assign _T_357 = btb_btype_1 != 2'h0; // @[BTB.scala 52:66:@1399.4]
  assign _T_359 = btb_btype_2 != 2'h0; // @[BTB.scala 52:66:@1400.4]
  assign _T_361 = btb_btype_3 != 2'h0; // @[BTB.scala 52:66:@1401.4]
  assign _T_363 = btb_btype_4 != 2'h0; // @[BTB.scala 52:66:@1402.4]
  assign _T_365 = btb_btype_5 != 2'h0; // @[BTB.scala 52:66:@1403.4]
  assign _T_367 = btb_btype_6 != 2'h0; // @[BTB.scala 52:66:@1404.4]
  assign _T_369 = btb_btype_7 != 2'h0; // @[BTB.scala 52:66:@1405.4]
  assign _T_371 = btb_btype_8 != 2'h0; // @[BTB.scala 52:66:@1406.4]
  assign _T_373 = btb_btype_9 != 2'h0; // @[BTB.scala 52:66:@1407.4]
  assign _T_375 = btb_btype_10 != 2'h0; // @[BTB.scala 52:66:@1408.4]
  assign _T_377 = btb_btype_11 != 2'h0; // @[BTB.scala 52:66:@1409.4]
  assign _T_379 = btb_btype_12 != 2'h0; // @[BTB.scala 52:66:@1410.4]
  assign _T_381 = btb_btype_13 != 2'h0; // @[BTB.scala 52:66:@1411.4]
  assign _T_383 = btb_btype_14 != 2'h0; // @[BTB.scala 52:66:@1412.4]
  assign _T_385 = btb_btype_15 != 2'h0; // @[BTB.scala 52:66:@1413.4]
  assign _T_387 = btb_btype_16 != 2'h0; // @[BTB.scala 52:66:@1414.4]
  assign _T_389 = btb_btype_17 != 2'h0; // @[BTB.scala 52:66:@1415.4]
  assign _T_391 = btb_btype_18 != 2'h0; // @[BTB.scala 52:66:@1416.4]
  assign _T_393 = btb_btype_19 != 2'h0; // @[BTB.scala 52:66:@1417.4]
  assign _T_395 = btb_btype_20 != 2'h0; // @[BTB.scala 52:66:@1418.4]
  assign _T_397 = btb_btype_21 != 2'h0; // @[BTB.scala 52:66:@1419.4]
  assign _T_399 = btb_btype_22 != 2'h0; // @[BTB.scala 52:66:@1420.4]
  assign _T_401 = btb_btype_23 != 2'h0; // @[BTB.scala 52:66:@1421.4]
  assign _T_403 = btb_btype_24 != 2'h0; // @[BTB.scala 52:66:@1422.4]
  assign _T_405 = btb_btype_25 != 2'h0; // @[BTB.scala 52:66:@1423.4]
  assign _T_407 = btb_btype_26 != 2'h0; // @[BTB.scala 52:66:@1424.4]
  assign _T_409 = btb_btype_27 != 2'h0; // @[BTB.scala 52:66:@1425.4]
  assign _T_411 = btb_btype_28 != 2'h0; // @[BTB.scala 52:66:@1426.4]
  assign _T_413 = btb_btype_29 != 2'h0; // @[BTB.scala 52:66:@1427.4]
  assign _T_415 = btb_btype_30 != 2'h0; // @[BTB.scala 52:66:@1428.4]
  assign _T_417 = btb_btype_31 != 2'h0; // @[BTB.scala 52:66:@1429.4]
  assign _T_419 = btb_btype_32 != 2'h0; // @[BTB.scala 52:66:@1430.4]
  assign _T_421 = btb_btype_33 != 2'h0; // @[BTB.scala 52:66:@1431.4]
  assign _T_423 = btb_btype_34 != 2'h0; // @[BTB.scala 52:66:@1432.4]
  assign _T_425 = btb_btype_35 != 2'h0; // @[BTB.scala 52:66:@1433.4]
  assign _T_427 = btb_btype_36 != 2'h0; // @[BTB.scala 52:66:@1434.4]
  assign _T_429 = btb_btype_37 != 2'h0; // @[BTB.scala 52:66:@1435.4]
  assign _T_431 = btb_btype_38 != 2'h0; // @[BTB.scala 52:66:@1436.4]
  assign _T_433 = btb_btype_39 != 2'h0; // @[BTB.scala 52:66:@1437.4]
  assign _T_435 = btb_btype_40 != 2'h0; // @[BTB.scala 52:66:@1438.4]
  assign _T_437 = btb_btype_41 != 2'h0; // @[BTB.scala 52:66:@1439.4]
  assign _T_439 = btb_btype_42 != 2'h0; // @[BTB.scala 52:66:@1440.4]
  assign _T_441 = btb_btype_43 != 2'h0; // @[BTB.scala 52:66:@1441.4]
  assign _T_443 = btb_btype_44 != 2'h0; // @[BTB.scala 52:66:@1442.4]
  assign _T_445 = btb_btype_45 != 2'h0; // @[BTB.scala 52:66:@1443.4]
  assign _T_447 = btb_btype_46 != 2'h0; // @[BTB.scala 52:66:@1444.4]
  assign _T_449 = btb_btype_47 != 2'h0; // @[BTB.scala 52:66:@1445.4]
  assign _T_451 = btb_btype_48 != 2'h0; // @[BTB.scala 52:66:@1446.4]
  assign _T_453 = btb_btype_49 != 2'h0; // @[BTB.scala 52:66:@1447.4]
  assign _T_455 = btb_btype_50 != 2'h0; // @[BTB.scala 52:66:@1448.4]
  assign _T_457 = btb_btype_51 != 2'h0; // @[BTB.scala 52:66:@1449.4]
  assign _T_459 = btb_btype_52 != 2'h0; // @[BTB.scala 52:66:@1450.4]
  assign _T_461 = btb_btype_53 != 2'h0; // @[BTB.scala 52:66:@1451.4]
  assign _T_463 = btb_btype_54 != 2'h0; // @[BTB.scala 52:66:@1452.4]
  assign _T_465 = btb_btype_55 != 2'h0; // @[BTB.scala 52:66:@1453.4]
  assign _T_467 = btb_btype_56 != 2'h0; // @[BTB.scala 52:66:@1454.4]
  assign _T_469 = btb_btype_57 != 2'h0; // @[BTB.scala 52:66:@1455.4]
  assign _T_471 = btb_btype_58 != 2'h0; // @[BTB.scala 52:66:@1456.4]
  assign _T_473 = btb_btype_59 != 2'h0; // @[BTB.scala 52:66:@1457.4]
  assign _T_475 = btb_btype_60 != 2'h0; // @[BTB.scala 52:66:@1458.4]
  assign _T_477 = btb_btype_61 != 2'h0; // @[BTB.scala 52:66:@1459.4]
  assign _T_479 = btb_btype_62 != 2'h0; // @[BTB.scala 52:66:@1460.4]
  assign _T_481 = btb_btype_63 != 2'h0; // @[BTB.scala 52:66:@1461.4]
  assign _T_558 = {_T_369,_T_367,_T_365,_T_363,_T_361,_T_359,_T_357,_T_355}; // @[BTB.scala 52:72:@1533.4]
  assign _T_566 = {_T_385,_T_383,_T_381,_T_379,_T_377,_T_375,_T_373,_T_371,_T_558}; // @[BTB.scala 52:72:@1541.4]
  assign _T_573 = {_T_401,_T_399,_T_397,_T_395,_T_393,_T_391,_T_389,_T_387}; // @[BTB.scala 52:72:@1548.4]
  assign _T_582 = {_T_417,_T_415,_T_413,_T_411,_T_409,_T_407,_T_405,_T_403,_T_573,_T_566}; // @[BTB.scala 52:72:@1557.4]
  assign _T_589 = {_T_433,_T_431,_T_429,_T_427,_T_425,_T_423,_T_421,_T_419}; // @[BTB.scala 52:72:@1564.4]
  assign _T_597 = {_T_449,_T_447,_T_445,_T_443,_T_441,_T_439,_T_437,_T_435,_T_589}; // @[BTB.scala 52:72:@1572.4]
  assign _T_604 = {_T_465,_T_463,_T_461,_T_459,_T_457,_T_455,_T_453,_T_451}; // @[BTB.scala 52:72:@1579.4]
  assign _T_613 = {_T_481,_T_479,_T_477,_T_475,_T_473,_T_471,_T_469,_T_467,_T_604,_T_597}; // @[BTB.scala 52:72:@1588.4]
  assign _T_614 = {_T_613,_T_582}; // @[BTB.scala 52:72:@1589.4]
  assign predict_0_lookup = _T_353 & _T_614; // @[BTB.scala 76:69:@1590.4]
  assign _T_616 = predict_0_lookup[0]; // @[Mux.scala 21:36:@1592.4]
  assign _T_617 = predict_0_lookup[1]; // @[Mux.scala 21:36:@1593.4]
  assign _T_618 = predict_0_lookup[2]; // @[Mux.scala 21:36:@1594.4]
  assign _T_619 = predict_0_lookup[3]; // @[Mux.scala 21:36:@1595.4]
  assign _T_620 = predict_0_lookup[4]; // @[Mux.scala 21:36:@1596.4]
  assign _T_621 = predict_0_lookup[5]; // @[Mux.scala 21:36:@1597.4]
  assign _T_622 = predict_0_lookup[6]; // @[Mux.scala 21:36:@1598.4]
  assign _T_623 = predict_0_lookup[7]; // @[Mux.scala 21:36:@1599.4]
  assign _T_624 = predict_0_lookup[8]; // @[Mux.scala 21:36:@1600.4]
  assign _T_625 = predict_0_lookup[9]; // @[Mux.scala 21:36:@1601.4]
  assign _T_626 = predict_0_lookup[10]; // @[Mux.scala 21:36:@1602.4]
  assign _T_627 = predict_0_lookup[11]; // @[Mux.scala 21:36:@1603.4]
  assign _T_628 = predict_0_lookup[12]; // @[Mux.scala 21:36:@1604.4]
  assign _T_629 = predict_0_lookup[13]; // @[Mux.scala 21:36:@1605.4]
  assign _T_630 = predict_0_lookup[14]; // @[Mux.scala 21:36:@1606.4]
  assign _T_631 = predict_0_lookup[15]; // @[Mux.scala 21:36:@1607.4]
  assign _T_632 = predict_0_lookup[16]; // @[Mux.scala 21:36:@1608.4]
  assign _T_633 = predict_0_lookup[17]; // @[Mux.scala 21:36:@1609.4]
  assign _T_634 = predict_0_lookup[18]; // @[Mux.scala 21:36:@1610.4]
  assign _T_635 = predict_0_lookup[19]; // @[Mux.scala 21:36:@1611.4]
  assign _T_636 = predict_0_lookup[20]; // @[Mux.scala 21:36:@1612.4]
  assign _T_637 = predict_0_lookup[21]; // @[Mux.scala 21:36:@1613.4]
  assign _T_638 = predict_0_lookup[22]; // @[Mux.scala 21:36:@1614.4]
  assign _T_639 = predict_0_lookup[23]; // @[Mux.scala 21:36:@1615.4]
  assign _T_640 = predict_0_lookup[24]; // @[Mux.scala 21:36:@1616.4]
  assign _T_641 = predict_0_lookup[25]; // @[Mux.scala 21:36:@1617.4]
  assign _T_642 = predict_0_lookup[26]; // @[Mux.scala 21:36:@1618.4]
  assign _T_643 = predict_0_lookup[27]; // @[Mux.scala 21:36:@1619.4]
  assign _T_644 = predict_0_lookup[28]; // @[Mux.scala 21:36:@1620.4]
  assign _T_645 = predict_0_lookup[29]; // @[Mux.scala 21:36:@1621.4]
  assign _T_646 = predict_0_lookup[30]; // @[Mux.scala 21:36:@1622.4]
  assign _T_647 = predict_0_lookup[31]; // @[Mux.scala 21:36:@1623.4]
  assign _T_648 = predict_0_lookup[32]; // @[Mux.scala 21:36:@1624.4]
  assign _T_649 = predict_0_lookup[33]; // @[Mux.scala 21:36:@1625.4]
  assign _T_650 = predict_0_lookup[34]; // @[Mux.scala 21:36:@1626.4]
  assign _T_651 = predict_0_lookup[35]; // @[Mux.scala 21:36:@1627.4]
  assign _T_652 = predict_0_lookup[36]; // @[Mux.scala 21:36:@1628.4]
  assign _T_653 = predict_0_lookup[37]; // @[Mux.scala 21:36:@1629.4]
  assign _T_654 = predict_0_lookup[38]; // @[Mux.scala 21:36:@1630.4]
  assign _T_655 = predict_0_lookup[39]; // @[Mux.scala 21:36:@1631.4]
  assign _T_656 = predict_0_lookup[40]; // @[Mux.scala 21:36:@1632.4]
  assign _T_657 = predict_0_lookup[41]; // @[Mux.scala 21:36:@1633.4]
  assign _T_658 = predict_0_lookup[42]; // @[Mux.scala 21:36:@1634.4]
  assign _T_659 = predict_0_lookup[43]; // @[Mux.scala 21:36:@1635.4]
  assign _T_660 = predict_0_lookup[44]; // @[Mux.scala 21:36:@1636.4]
  assign _T_661 = predict_0_lookup[45]; // @[Mux.scala 21:36:@1637.4]
  assign _T_662 = predict_0_lookup[46]; // @[Mux.scala 21:36:@1638.4]
  assign _T_663 = predict_0_lookup[47]; // @[Mux.scala 21:36:@1639.4]
  assign _T_664 = predict_0_lookup[48]; // @[Mux.scala 21:36:@1640.4]
  assign _T_665 = predict_0_lookup[49]; // @[Mux.scala 21:36:@1641.4]
  assign _T_666 = predict_0_lookup[50]; // @[Mux.scala 21:36:@1642.4]
  assign _T_667 = predict_0_lookup[51]; // @[Mux.scala 21:36:@1643.4]
  assign _T_668 = predict_0_lookup[52]; // @[Mux.scala 21:36:@1644.4]
  assign _T_669 = predict_0_lookup[53]; // @[Mux.scala 21:36:@1645.4]
  assign _T_670 = predict_0_lookup[54]; // @[Mux.scala 21:36:@1646.4]
  assign _T_671 = predict_0_lookup[55]; // @[Mux.scala 21:36:@1647.4]
  assign _T_672 = predict_0_lookup[56]; // @[Mux.scala 21:36:@1648.4]
  assign _T_673 = predict_0_lookup[57]; // @[Mux.scala 21:36:@1649.4]
  assign _T_674 = predict_0_lookup[58]; // @[Mux.scala 21:36:@1650.4]
  assign _T_675 = predict_0_lookup[59]; // @[Mux.scala 21:36:@1651.4]
  assign _T_676 = predict_0_lookup[60]; // @[Mux.scala 21:36:@1652.4]
  assign _T_677 = predict_0_lookup[61]; // @[Mux.scala 21:36:@1653.4]
  assign _T_678 = predict_0_lookup[62]; // @[Mux.scala 21:36:@1654.4]
  assign _T_679 = predict_0_lookup[63]; // @[Mux.scala 21:36:@1655.4]
  assign _T_682 = _T_616 ? btb_target_0 : 32'h0; // @[Mux.scala 19:72:@1656.4]
  assign _T_684 = _T_617 ? btb_target_1 : 32'h0; // @[Mux.scala 19:72:@1657.4]
  assign _T_686 = _T_618 ? btb_target_2 : 32'h0; // @[Mux.scala 19:72:@1658.4]
  assign _T_688 = _T_619 ? btb_target_3 : 32'h0; // @[Mux.scala 19:72:@1659.4]
  assign _T_690 = _T_620 ? btb_target_4 : 32'h0; // @[Mux.scala 19:72:@1660.4]
  assign _T_692 = _T_621 ? btb_target_5 : 32'h0; // @[Mux.scala 19:72:@1661.4]
  assign _T_694 = _T_622 ? btb_target_6 : 32'h0; // @[Mux.scala 19:72:@1662.4]
  assign _T_696 = _T_623 ? btb_target_7 : 32'h0; // @[Mux.scala 19:72:@1663.4]
  assign _T_698 = _T_624 ? btb_target_8 : 32'h0; // @[Mux.scala 19:72:@1664.4]
  assign _T_700 = _T_625 ? btb_target_9 : 32'h0; // @[Mux.scala 19:72:@1665.4]
  assign _T_702 = _T_626 ? btb_target_10 : 32'h0; // @[Mux.scala 19:72:@1666.4]
  assign _T_704 = _T_627 ? btb_target_11 : 32'h0; // @[Mux.scala 19:72:@1667.4]
  assign _T_706 = _T_628 ? btb_target_12 : 32'h0; // @[Mux.scala 19:72:@1668.4]
  assign _T_708 = _T_629 ? btb_target_13 : 32'h0; // @[Mux.scala 19:72:@1669.4]
  assign _T_710 = _T_630 ? btb_target_14 : 32'h0; // @[Mux.scala 19:72:@1670.4]
  assign _T_712 = _T_631 ? btb_target_15 : 32'h0; // @[Mux.scala 19:72:@1671.4]
  assign _T_714 = _T_632 ? btb_target_16 : 32'h0; // @[Mux.scala 19:72:@1672.4]
  assign _T_716 = _T_633 ? btb_target_17 : 32'h0; // @[Mux.scala 19:72:@1673.4]
  assign _T_718 = _T_634 ? btb_target_18 : 32'h0; // @[Mux.scala 19:72:@1674.4]
  assign _T_720 = _T_635 ? btb_target_19 : 32'h0; // @[Mux.scala 19:72:@1675.4]
  assign _T_722 = _T_636 ? btb_target_20 : 32'h0; // @[Mux.scala 19:72:@1676.4]
  assign _T_724 = _T_637 ? btb_target_21 : 32'h0; // @[Mux.scala 19:72:@1677.4]
  assign _T_726 = _T_638 ? btb_target_22 : 32'h0; // @[Mux.scala 19:72:@1678.4]
  assign _T_728 = _T_639 ? btb_target_23 : 32'h0; // @[Mux.scala 19:72:@1679.4]
  assign _T_730 = _T_640 ? btb_target_24 : 32'h0; // @[Mux.scala 19:72:@1680.4]
  assign _T_732 = _T_641 ? btb_target_25 : 32'h0; // @[Mux.scala 19:72:@1681.4]
  assign _T_734 = _T_642 ? btb_target_26 : 32'h0; // @[Mux.scala 19:72:@1682.4]
  assign _T_736 = _T_643 ? btb_target_27 : 32'h0; // @[Mux.scala 19:72:@1683.4]
  assign _T_738 = _T_644 ? btb_target_28 : 32'h0; // @[Mux.scala 19:72:@1684.4]
  assign _T_740 = _T_645 ? btb_target_29 : 32'h0; // @[Mux.scala 19:72:@1685.4]
  assign _T_742 = _T_646 ? btb_target_30 : 32'h0; // @[Mux.scala 19:72:@1686.4]
  assign _T_744 = _T_647 ? btb_target_31 : 32'h0; // @[Mux.scala 19:72:@1687.4]
  assign _T_746 = _T_648 ? btb_target_32 : 32'h0; // @[Mux.scala 19:72:@1688.4]
  assign _T_748 = _T_649 ? btb_target_33 : 32'h0; // @[Mux.scala 19:72:@1689.4]
  assign _T_750 = _T_650 ? btb_target_34 : 32'h0; // @[Mux.scala 19:72:@1690.4]
  assign _T_752 = _T_651 ? btb_target_35 : 32'h0; // @[Mux.scala 19:72:@1691.4]
  assign _T_754 = _T_652 ? btb_target_36 : 32'h0; // @[Mux.scala 19:72:@1692.4]
  assign _T_756 = _T_653 ? btb_target_37 : 32'h0; // @[Mux.scala 19:72:@1693.4]
  assign _T_758 = _T_654 ? btb_target_38 : 32'h0; // @[Mux.scala 19:72:@1694.4]
  assign _T_760 = _T_655 ? btb_target_39 : 32'h0; // @[Mux.scala 19:72:@1695.4]
  assign _T_762 = _T_656 ? btb_target_40 : 32'h0; // @[Mux.scala 19:72:@1696.4]
  assign _T_764 = _T_657 ? btb_target_41 : 32'h0; // @[Mux.scala 19:72:@1697.4]
  assign _T_766 = _T_658 ? btb_target_42 : 32'h0; // @[Mux.scala 19:72:@1698.4]
  assign _T_768 = _T_659 ? btb_target_43 : 32'h0; // @[Mux.scala 19:72:@1699.4]
  assign _T_770 = _T_660 ? btb_target_44 : 32'h0; // @[Mux.scala 19:72:@1700.4]
  assign _T_772 = _T_661 ? btb_target_45 : 32'h0; // @[Mux.scala 19:72:@1701.4]
  assign _T_774 = _T_662 ? btb_target_46 : 32'h0; // @[Mux.scala 19:72:@1702.4]
  assign _T_776 = _T_663 ? btb_target_47 : 32'h0; // @[Mux.scala 19:72:@1703.4]
  assign _T_778 = _T_664 ? btb_target_48 : 32'h0; // @[Mux.scala 19:72:@1704.4]
  assign _T_780 = _T_665 ? btb_target_49 : 32'h0; // @[Mux.scala 19:72:@1705.4]
  assign _T_782 = _T_666 ? btb_target_50 : 32'h0; // @[Mux.scala 19:72:@1706.4]
  assign _T_784 = _T_667 ? btb_target_51 : 32'h0; // @[Mux.scala 19:72:@1707.4]
  assign _T_786 = _T_668 ? btb_target_52 : 32'h0; // @[Mux.scala 19:72:@1708.4]
  assign _T_788 = _T_669 ? btb_target_53 : 32'h0; // @[Mux.scala 19:72:@1709.4]
  assign _T_790 = _T_670 ? btb_target_54 : 32'h0; // @[Mux.scala 19:72:@1710.4]
  assign _T_792 = _T_671 ? btb_target_55 : 32'h0; // @[Mux.scala 19:72:@1711.4]
  assign _T_794 = _T_672 ? btb_target_56 : 32'h0; // @[Mux.scala 19:72:@1712.4]
  assign _T_796 = _T_673 ? btb_target_57 : 32'h0; // @[Mux.scala 19:72:@1713.4]
  assign _T_798 = _T_674 ? btb_target_58 : 32'h0; // @[Mux.scala 19:72:@1714.4]
  assign _T_800 = _T_675 ? btb_target_59 : 32'h0; // @[Mux.scala 19:72:@1715.4]
  assign _T_802 = _T_676 ? btb_target_60 : 32'h0; // @[Mux.scala 19:72:@1716.4]
  assign _T_804 = _T_677 ? btb_target_61 : 32'h0; // @[Mux.scala 19:72:@1717.4]
  assign _T_806 = _T_678 ? btb_target_62 : 32'h0; // @[Mux.scala 19:72:@1718.4]
  assign _T_808 = _T_679 ? btb_target_63 : 32'h0; // @[Mux.scala 19:72:@1719.4]
  assign _T_809 = _T_682 | _T_684; // @[Mux.scala 19:72:@1720.4]
  assign _T_810 = _T_809 | _T_686; // @[Mux.scala 19:72:@1721.4]
  assign _T_811 = _T_810 | _T_688; // @[Mux.scala 19:72:@1722.4]
  assign _T_812 = _T_811 | _T_690; // @[Mux.scala 19:72:@1723.4]
  assign _T_813 = _T_812 | _T_692; // @[Mux.scala 19:72:@1724.4]
  assign _T_814 = _T_813 | _T_694; // @[Mux.scala 19:72:@1725.4]
  assign _T_815 = _T_814 | _T_696; // @[Mux.scala 19:72:@1726.4]
  assign _T_816 = _T_815 | _T_698; // @[Mux.scala 19:72:@1727.4]
  assign _T_817 = _T_816 | _T_700; // @[Mux.scala 19:72:@1728.4]
  assign _T_818 = _T_817 | _T_702; // @[Mux.scala 19:72:@1729.4]
  assign _T_819 = _T_818 | _T_704; // @[Mux.scala 19:72:@1730.4]
  assign _T_820 = _T_819 | _T_706; // @[Mux.scala 19:72:@1731.4]
  assign _T_821 = _T_820 | _T_708; // @[Mux.scala 19:72:@1732.4]
  assign _T_822 = _T_821 | _T_710; // @[Mux.scala 19:72:@1733.4]
  assign _T_823 = _T_822 | _T_712; // @[Mux.scala 19:72:@1734.4]
  assign _T_824 = _T_823 | _T_714; // @[Mux.scala 19:72:@1735.4]
  assign _T_825 = _T_824 | _T_716; // @[Mux.scala 19:72:@1736.4]
  assign _T_826 = _T_825 | _T_718; // @[Mux.scala 19:72:@1737.4]
  assign _T_827 = _T_826 | _T_720; // @[Mux.scala 19:72:@1738.4]
  assign _T_828 = _T_827 | _T_722; // @[Mux.scala 19:72:@1739.4]
  assign _T_829 = _T_828 | _T_724; // @[Mux.scala 19:72:@1740.4]
  assign _T_830 = _T_829 | _T_726; // @[Mux.scala 19:72:@1741.4]
  assign _T_831 = _T_830 | _T_728; // @[Mux.scala 19:72:@1742.4]
  assign _T_832 = _T_831 | _T_730; // @[Mux.scala 19:72:@1743.4]
  assign _T_833 = _T_832 | _T_732; // @[Mux.scala 19:72:@1744.4]
  assign _T_834 = _T_833 | _T_734; // @[Mux.scala 19:72:@1745.4]
  assign _T_835 = _T_834 | _T_736; // @[Mux.scala 19:72:@1746.4]
  assign _T_836 = _T_835 | _T_738; // @[Mux.scala 19:72:@1747.4]
  assign _T_837 = _T_836 | _T_740; // @[Mux.scala 19:72:@1748.4]
  assign _T_838 = _T_837 | _T_742; // @[Mux.scala 19:72:@1749.4]
  assign _T_839 = _T_838 | _T_744; // @[Mux.scala 19:72:@1750.4]
  assign _T_840 = _T_839 | _T_746; // @[Mux.scala 19:72:@1751.4]
  assign _T_841 = _T_840 | _T_748; // @[Mux.scala 19:72:@1752.4]
  assign _T_842 = _T_841 | _T_750; // @[Mux.scala 19:72:@1753.4]
  assign _T_843 = _T_842 | _T_752; // @[Mux.scala 19:72:@1754.4]
  assign _T_844 = _T_843 | _T_754; // @[Mux.scala 19:72:@1755.4]
  assign _T_845 = _T_844 | _T_756; // @[Mux.scala 19:72:@1756.4]
  assign _T_846 = _T_845 | _T_758; // @[Mux.scala 19:72:@1757.4]
  assign _T_847 = _T_846 | _T_760; // @[Mux.scala 19:72:@1758.4]
  assign _T_848 = _T_847 | _T_762; // @[Mux.scala 19:72:@1759.4]
  assign _T_849 = _T_848 | _T_764; // @[Mux.scala 19:72:@1760.4]
  assign _T_850 = _T_849 | _T_766; // @[Mux.scala 19:72:@1761.4]
  assign _T_851 = _T_850 | _T_768; // @[Mux.scala 19:72:@1762.4]
  assign _T_852 = _T_851 | _T_770; // @[Mux.scala 19:72:@1763.4]
  assign _T_853 = _T_852 | _T_772; // @[Mux.scala 19:72:@1764.4]
  assign _T_854 = _T_853 | _T_774; // @[Mux.scala 19:72:@1765.4]
  assign _T_855 = _T_854 | _T_776; // @[Mux.scala 19:72:@1766.4]
  assign _T_856 = _T_855 | _T_778; // @[Mux.scala 19:72:@1767.4]
  assign _T_857 = _T_856 | _T_780; // @[Mux.scala 19:72:@1768.4]
  assign _T_858 = _T_857 | _T_782; // @[Mux.scala 19:72:@1769.4]
  assign _T_859 = _T_858 | _T_784; // @[Mux.scala 19:72:@1770.4]
  assign _T_860 = _T_859 | _T_786; // @[Mux.scala 19:72:@1771.4]
  assign _T_861 = _T_860 | _T_788; // @[Mux.scala 19:72:@1772.4]
  assign _T_862 = _T_861 | _T_790; // @[Mux.scala 19:72:@1773.4]
  assign _T_863 = _T_862 | _T_792; // @[Mux.scala 19:72:@1774.4]
  assign _T_864 = _T_863 | _T_794; // @[Mux.scala 19:72:@1775.4]
  assign _T_865 = _T_864 | _T_796; // @[Mux.scala 19:72:@1776.4]
  assign _T_866 = _T_865 | _T_798; // @[Mux.scala 19:72:@1777.4]
  assign _T_867 = _T_866 | _T_800; // @[Mux.scala 19:72:@1778.4]
  assign _T_868 = _T_867 | _T_802; // @[Mux.scala 19:72:@1779.4]
  assign _T_869 = _T_868 | _T_804; // @[Mux.scala 19:72:@1780.4]
  assign _T_870 = _T_869 | _T_806; // @[Mux.scala 19:72:@1781.4]
  assign predict_0_jump_tgt = _T_870 | _T_808; // @[Mux.scala 19:72:@1782.4]
  assign _T_940 = _T_616 ? btb_btype_0 : 2'h0; // @[Mux.scala 19:72:@1850.4]
  assign _T_942 = _T_617 ? btb_btype_1 : 2'h0; // @[Mux.scala 19:72:@1851.4]
  assign _T_944 = _T_618 ? btb_btype_2 : 2'h0; // @[Mux.scala 19:72:@1852.4]
  assign _T_946 = _T_619 ? btb_btype_3 : 2'h0; // @[Mux.scala 19:72:@1853.4]
  assign _T_948 = _T_620 ? btb_btype_4 : 2'h0; // @[Mux.scala 19:72:@1854.4]
  assign _T_950 = _T_621 ? btb_btype_5 : 2'h0; // @[Mux.scala 19:72:@1855.4]
  assign _T_952 = _T_622 ? btb_btype_6 : 2'h0; // @[Mux.scala 19:72:@1856.4]
  assign _T_954 = _T_623 ? btb_btype_7 : 2'h0; // @[Mux.scala 19:72:@1857.4]
  assign _T_956 = _T_624 ? btb_btype_8 : 2'h0; // @[Mux.scala 19:72:@1858.4]
  assign _T_958 = _T_625 ? btb_btype_9 : 2'h0; // @[Mux.scala 19:72:@1859.4]
  assign _T_960 = _T_626 ? btb_btype_10 : 2'h0; // @[Mux.scala 19:72:@1860.4]
  assign _T_962 = _T_627 ? btb_btype_11 : 2'h0; // @[Mux.scala 19:72:@1861.4]
  assign _T_964 = _T_628 ? btb_btype_12 : 2'h0; // @[Mux.scala 19:72:@1862.4]
  assign _T_966 = _T_629 ? btb_btype_13 : 2'h0; // @[Mux.scala 19:72:@1863.4]
  assign _T_968 = _T_630 ? btb_btype_14 : 2'h0; // @[Mux.scala 19:72:@1864.4]
  assign _T_970 = _T_631 ? btb_btype_15 : 2'h0; // @[Mux.scala 19:72:@1865.4]
  assign _T_972 = _T_632 ? btb_btype_16 : 2'h0; // @[Mux.scala 19:72:@1866.4]
  assign _T_974 = _T_633 ? btb_btype_17 : 2'h0; // @[Mux.scala 19:72:@1867.4]
  assign _T_976 = _T_634 ? btb_btype_18 : 2'h0; // @[Mux.scala 19:72:@1868.4]
  assign _T_978 = _T_635 ? btb_btype_19 : 2'h0; // @[Mux.scala 19:72:@1869.4]
  assign _T_980 = _T_636 ? btb_btype_20 : 2'h0; // @[Mux.scala 19:72:@1870.4]
  assign _T_982 = _T_637 ? btb_btype_21 : 2'h0; // @[Mux.scala 19:72:@1871.4]
  assign _T_984 = _T_638 ? btb_btype_22 : 2'h0; // @[Mux.scala 19:72:@1872.4]
  assign _T_986 = _T_639 ? btb_btype_23 : 2'h0; // @[Mux.scala 19:72:@1873.4]
  assign _T_988 = _T_640 ? btb_btype_24 : 2'h0; // @[Mux.scala 19:72:@1874.4]
  assign _T_990 = _T_641 ? btb_btype_25 : 2'h0; // @[Mux.scala 19:72:@1875.4]
  assign _T_992 = _T_642 ? btb_btype_26 : 2'h0; // @[Mux.scala 19:72:@1876.4]
  assign _T_994 = _T_643 ? btb_btype_27 : 2'h0; // @[Mux.scala 19:72:@1877.4]
  assign _T_996 = _T_644 ? btb_btype_28 : 2'h0; // @[Mux.scala 19:72:@1878.4]
  assign _T_998 = _T_645 ? btb_btype_29 : 2'h0; // @[Mux.scala 19:72:@1879.4]
  assign _T_1000 = _T_646 ? btb_btype_30 : 2'h0; // @[Mux.scala 19:72:@1880.4]
  assign _T_1002 = _T_647 ? btb_btype_31 : 2'h0; // @[Mux.scala 19:72:@1881.4]
  assign _T_1004 = _T_648 ? btb_btype_32 : 2'h0; // @[Mux.scala 19:72:@1882.4]
  assign _T_1006 = _T_649 ? btb_btype_33 : 2'h0; // @[Mux.scala 19:72:@1883.4]
  assign _T_1008 = _T_650 ? btb_btype_34 : 2'h0; // @[Mux.scala 19:72:@1884.4]
  assign _T_1010 = _T_651 ? btb_btype_35 : 2'h0; // @[Mux.scala 19:72:@1885.4]
  assign _T_1012 = _T_652 ? btb_btype_36 : 2'h0; // @[Mux.scala 19:72:@1886.4]
  assign _T_1014 = _T_653 ? btb_btype_37 : 2'h0; // @[Mux.scala 19:72:@1887.4]
  assign _T_1016 = _T_654 ? btb_btype_38 : 2'h0; // @[Mux.scala 19:72:@1888.4]
  assign _T_1018 = _T_655 ? btb_btype_39 : 2'h0; // @[Mux.scala 19:72:@1889.4]
  assign _T_1020 = _T_656 ? btb_btype_40 : 2'h0; // @[Mux.scala 19:72:@1890.4]
  assign _T_1022 = _T_657 ? btb_btype_41 : 2'h0; // @[Mux.scala 19:72:@1891.4]
  assign _T_1024 = _T_658 ? btb_btype_42 : 2'h0; // @[Mux.scala 19:72:@1892.4]
  assign _T_1026 = _T_659 ? btb_btype_43 : 2'h0; // @[Mux.scala 19:72:@1893.4]
  assign _T_1028 = _T_660 ? btb_btype_44 : 2'h0; // @[Mux.scala 19:72:@1894.4]
  assign _T_1030 = _T_661 ? btb_btype_45 : 2'h0; // @[Mux.scala 19:72:@1895.4]
  assign _T_1032 = _T_662 ? btb_btype_46 : 2'h0; // @[Mux.scala 19:72:@1896.4]
  assign _T_1034 = _T_663 ? btb_btype_47 : 2'h0; // @[Mux.scala 19:72:@1897.4]
  assign _T_1036 = _T_664 ? btb_btype_48 : 2'h0; // @[Mux.scala 19:72:@1898.4]
  assign _T_1038 = _T_665 ? btb_btype_49 : 2'h0; // @[Mux.scala 19:72:@1899.4]
  assign _T_1040 = _T_666 ? btb_btype_50 : 2'h0; // @[Mux.scala 19:72:@1900.4]
  assign _T_1042 = _T_667 ? btb_btype_51 : 2'h0; // @[Mux.scala 19:72:@1901.4]
  assign _T_1044 = _T_668 ? btb_btype_52 : 2'h0; // @[Mux.scala 19:72:@1902.4]
  assign _T_1046 = _T_669 ? btb_btype_53 : 2'h0; // @[Mux.scala 19:72:@1903.4]
  assign _T_1048 = _T_670 ? btb_btype_54 : 2'h0; // @[Mux.scala 19:72:@1904.4]
  assign _T_1050 = _T_671 ? btb_btype_55 : 2'h0; // @[Mux.scala 19:72:@1905.4]
  assign _T_1052 = _T_672 ? btb_btype_56 : 2'h0; // @[Mux.scala 19:72:@1906.4]
  assign _T_1054 = _T_673 ? btb_btype_57 : 2'h0; // @[Mux.scala 19:72:@1907.4]
  assign _T_1056 = _T_674 ? btb_btype_58 : 2'h0; // @[Mux.scala 19:72:@1908.4]
  assign _T_1058 = _T_675 ? btb_btype_59 : 2'h0; // @[Mux.scala 19:72:@1909.4]
  assign _T_1060 = _T_676 ? btb_btype_60 : 2'h0; // @[Mux.scala 19:72:@1910.4]
  assign _T_1062 = _T_677 ? btb_btype_61 : 2'h0; // @[Mux.scala 19:72:@1911.4]
  assign _T_1064 = _T_678 ? btb_btype_62 : 2'h0; // @[Mux.scala 19:72:@1912.4]
  assign _T_1066 = _T_679 ? btb_btype_63 : 2'h0; // @[Mux.scala 19:72:@1913.4]
  assign _T_1067 = _T_940 | _T_942; // @[Mux.scala 19:72:@1914.4]
  assign _T_1068 = _T_1067 | _T_944; // @[Mux.scala 19:72:@1915.4]
  assign _T_1069 = _T_1068 | _T_946; // @[Mux.scala 19:72:@1916.4]
  assign _T_1070 = _T_1069 | _T_948; // @[Mux.scala 19:72:@1917.4]
  assign _T_1071 = _T_1070 | _T_950; // @[Mux.scala 19:72:@1918.4]
  assign _T_1072 = _T_1071 | _T_952; // @[Mux.scala 19:72:@1919.4]
  assign _T_1073 = _T_1072 | _T_954; // @[Mux.scala 19:72:@1920.4]
  assign _T_1074 = _T_1073 | _T_956; // @[Mux.scala 19:72:@1921.4]
  assign _T_1075 = _T_1074 | _T_958; // @[Mux.scala 19:72:@1922.4]
  assign _T_1076 = _T_1075 | _T_960; // @[Mux.scala 19:72:@1923.4]
  assign _T_1077 = _T_1076 | _T_962; // @[Mux.scala 19:72:@1924.4]
  assign _T_1078 = _T_1077 | _T_964; // @[Mux.scala 19:72:@1925.4]
  assign _T_1079 = _T_1078 | _T_966; // @[Mux.scala 19:72:@1926.4]
  assign _T_1080 = _T_1079 | _T_968; // @[Mux.scala 19:72:@1927.4]
  assign _T_1081 = _T_1080 | _T_970; // @[Mux.scala 19:72:@1928.4]
  assign _T_1082 = _T_1081 | _T_972; // @[Mux.scala 19:72:@1929.4]
  assign _T_1083 = _T_1082 | _T_974; // @[Mux.scala 19:72:@1930.4]
  assign _T_1084 = _T_1083 | _T_976; // @[Mux.scala 19:72:@1931.4]
  assign _T_1085 = _T_1084 | _T_978; // @[Mux.scala 19:72:@1932.4]
  assign _T_1086 = _T_1085 | _T_980; // @[Mux.scala 19:72:@1933.4]
  assign _T_1087 = _T_1086 | _T_982; // @[Mux.scala 19:72:@1934.4]
  assign _T_1088 = _T_1087 | _T_984; // @[Mux.scala 19:72:@1935.4]
  assign _T_1089 = _T_1088 | _T_986; // @[Mux.scala 19:72:@1936.4]
  assign _T_1090 = _T_1089 | _T_988; // @[Mux.scala 19:72:@1937.4]
  assign _T_1091 = _T_1090 | _T_990; // @[Mux.scala 19:72:@1938.4]
  assign _T_1092 = _T_1091 | _T_992; // @[Mux.scala 19:72:@1939.4]
  assign _T_1093 = _T_1092 | _T_994; // @[Mux.scala 19:72:@1940.4]
  assign _T_1094 = _T_1093 | _T_996; // @[Mux.scala 19:72:@1941.4]
  assign _T_1095 = _T_1094 | _T_998; // @[Mux.scala 19:72:@1942.4]
  assign _T_1096 = _T_1095 | _T_1000; // @[Mux.scala 19:72:@1943.4]
  assign _T_1097 = _T_1096 | _T_1002; // @[Mux.scala 19:72:@1944.4]
  assign _T_1098 = _T_1097 | _T_1004; // @[Mux.scala 19:72:@1945.4]
  assign _T_1099 = _T_1098 | _T_1006; // @[Mux.scala 19:72:@1946.4]
  assign _T_1100 = _T_1099 | _T_1008; // @[Mux.scala 19:72:@1947.4]
  assign _T_1101 = _T_1100 | _T_1010; // @[Mux.scala 19:72:@1948.4]
  assign _T_1102 = _T_1101 | _T_1012; // @[Mux.scala 19:72:@1949.4]
  assign _T_1103 = _T_1102 | _T_1014; // @[Mux.scala 19:72:@1950.4]
  assign _T_1104 = _T_1103 | _T_1016; // @[Mux.scala 19:72:@1951.4]
  assign _T_1105 = _T_1104 | _T_1018; // @[Mux.scala 19:72:@1952.4]
  assign _T_1106 = _T_1105 | _T_1020; // @[Mux.scala 19:72:@1953.4]
  assign _T_1107 = _T_1106 | _T_1022; // @[Mux.scala 19:72:@1954.4]
  assign _T_1108 = _T_1107 | _T_1024; // @[Mux.scala 19:72:@1955.4]
  assign _T_1109 = _T_1108 | _T_1026; // @[Mux.scala 19:72:@1956.4]
  assign _T_1110 = _T_1109 | _T_1028; // @[Mux.scala 19:72:@1957.4]
  assign _T_1111 = _T_1110 | _T_1030; // @[Mux.scala 19:72:@1958.4]
  assign _T_1112 = _T_1111 | _T_1032; // @[Mux.scala 19:72:@1959.4]
  assign _T_1113 = _T_1112 | _T_1034; // @[Mux.scala 19:72:@1960.4]
  assign _T_1114 = _T_1113 | _T_1036; // @[Mux.scala 19:72:@1961.4]
  assign _T_1115 = _T_1114 | _T_1038; // @[Mux.scala 19:72:@1962.4]
  assign _T_1116 = _T_1115 | _T_1040; // @[Mux.scala 19:72:@1963.4]
  assign _T_1117 = _T_1116 | _T_1042; // @[Mux.scala 19:72:@1964.4]
  assign _T_1118 = _T_1117 | _T_1044; // @[Mux.scala 19:72:@1965.4]
  assign _T_1119 = _T_1118 | _T_1046; // @[Mux.scala 19:72:@1966.4]
  assign _T_1120 = _T_1119 | _T_1048; // @[Mux.scala 19:72:@1967.4]
  assign _T_1121 = _T_1120 | _T_1050; // @[Mux.scala 19:72:@1968.4]
  assign _T_1122 = _T_1121 | _T_1052; // @[Mux.scala 19:72:@1969.4]
  assign _T_1123 = _T_1122 | _T_1054; // @[Mux.scala 19:72:@1970.4]
  assign _T_1124 = _T_1123 | _T_1056; // @[Mux.scala 19:72:@1971.4]
  assign _T_1125 = _T_1124 | _T_1058; // @[Mux.scala 19:72:@1972.4]
  assign _T_1126 = _T_1125 | _T_1060; // @[Mux.scala 19:72:@1973.4]
  assign _T_1127 = _T_1126 | _T_1062; // @[Mux.scala 19:72:@1974.4]
  assign _T_1128 = _T_1127 | _T_1064; // @[Mux.scala 19:72:@1975.4]
  assign predict_0_btype = _T_1128 | _T_1066; // @[Mux.scala 19:72:@1976.4]
  assign _T_1198 = _T_616 ? btb_hcount_0 : 2'h0; // @[Mux.scala 19:72:@2044.4]
  assign _T_1200 = _T_617 ? btb_hcount_1 : 2'h0; // @[Mux.scala 19:72:@2045.4]
  assign _T_1202 = _T_618 ? btb_hcount_2 : 2'h0; // @[Mux.scala 19:72:@2046.4]
  assign _T_1204 = _T_619 ? btb_hcount_3 : 2'h0; // @[Mux.scala 19:72:@2047.4]
  assign _T_1206 = _T_620 ? btb_hcount_4 : 2'h0; // @[Mux.scala 19:72:@2048.4]
  assign _T_1208 = _T_621 ? btb_hcount_5 : 2'h0; // @[Mux.scala 19:72:@2049.4]
  assign _T_1210 = _T_622 ? btb_hcount_6 : 2'h0; // @[Mux.scala 19:72:@2050.4]
  assign _T_1212 = _T_623 ? btb_hcount_7 : 2'h0; // @[Mux.scala 19:72:@2051.4]
  assign _T_1214 = _T_624 ? btb_hcount_8 : 2'h0; // @[Mux.scala 19:72:@2052.4]
  assign _T_1216 = _T_625 ? btb_hcount_9 : 2'h0; // @[Mux.scala 19:72:@2053.4]
  assign _T_1218 = _T_626 ? btb_hcount_10 : 2'h0; // @[Mux.scala 19:72:@2054.4]
  assign _T_1220 = _T_627 ? btb_hcount_11 : 2'h0; // @[Mux.scala 19:72:@2055.4]
  assign _T_1222 = _T_628 ? btb_hcount_12 : 2'h0; // @[Mux.scala 19:72:@2056.4]
  assign _T_1224 = _T_629 ? btb_hcount_13 : 2'h0; // @[Mux.scala 19:72:@2057.4]
  assign _T_1226 = _T_630 ? btb_hcount_14 : 2'h0; // @[Mux.scala 19:72:@2058.4]
  assign _T_1228 = _T_631 ? btb_hcount_15 : 2'h0; // @[Mux.scala 19:72:@2059.4]
  assign _T_1230 = _T_632 ? btb_hcount_16 : 2'h0; // @[Mux.scala 19:72:@2060.4]
  assign _T_1232 = _T_633 ? btb_hcount_17 : 2'h0; // @[Mux.scala 19:72:@2061.4]
  assign _T_1234 = _T_634 ? btb_hcount_18 : 2'h0; // @[Mux.scala 19:72:@2062.4]
  assign _T_1236 = _T_635 ? btb_hcount_19 : 2'h0; // @[Mux.scala 19:72:@2063.4]
  assign _T_1238 = _T_636 ? btb_hcount_20 : 2'h0; // @[Mux.scala 19:72:@2064.4]
  assign _T_1240 = _T_637 ? btb_hcount_21 : 2'h0; // @[Mux.scala 19:72:@2065.4]
  assign _T_1242 = _T_638 ? btb_hcount_22 : 2'h0; // @[Mux.scala 19:72:@2066.4]
  assign _T_1244 = _T_639 ? btb_hcount_23 : 2'h0; // @[Mux.scala 19:72:@2067.4]
  assign _T_1246 = _T_640 ? btb_hcount_24 : 2'h0; // @[Mux.scala 19:72:@2068.4]
  assign _T_1248 = _T_641 ? btb_hcount_25 : 2'h0; // @[Mux.scala 19:72:@2069.4]
  assign _T_1250 = _T_642 ? btb_hcount_26 : 2'h0; // @[Mux.scala 19:72:@2070.4]
  assign _T_1252 = _T_643 ? btb_hcount_27 : 2'h0; // @[Mux.scala 19:72:@2071.4]
  assign _T_1254 = _T_644 ? btb_hcount_28 : 2'h0; // @[Mux.scala 19:72:@2072.4]
  assign _T_1256 = _T_645 ? btb_hcount_29 : 2'h0; // @[Mux.scala 19:72:@2073.4]
  assign _T_1258 = _T_646 ? btb_hcount_30 : 2'h0; // @[Mux.scala 19:72:@2074.4]
  assign _T_1260 = _T_647 ? btb_hcount_31 : 2'h0; // @[Mux.scala 19:72:@2075.4]
  assign _T_1262 = _T_648 ? btb_hcount_32 : 2'h0; // @[Mux.scala 19:72:@2076.4]
  assign _T_1264 = _T_649 ? btb_hcount_33 : 2'h0; // @[Mux.scala 19:72:@2077.4]
  assign _T_1266 = _T_650 ? btb_hcount_34 : 2'h0; // @[Mux.scala 19:72:@2078.4]
  assign _T_1268 = _T_651 ? btb_hcount_35 : 2'h0; // @[Mux.scala 19:72:@2079.4]
  assign _T_1270 = _T_652 ? btb_hcount_36 : 2'h0; // @[Mux.scala 19:72:@2080.4]
  assign _T_1272 = _T_653 ? btb_hcount_37 : 2'h0; // @[Mux.scala 19:72:@2081.4]
  assign _T_1274 = _T_654 ? btb_hcount_38 : 2'h0; // @[Mux.scala 19:72:@2082.4]
  assign _T_1276 = _T_655 ? btb_hcount_39 : 2'h0; // @[Mux.scala 19:72:@2083.4]
  assign _T_1278 = _T_656 ? btb_hcount_40 : 2'h0; // @[Mux.scala 19:72:@2084.4]
  assign _T_1280 = _T_657 ? btb_hcount_41 : 2'h0; // @[Mux.scala 19:72:@2085.4]
  assign _T_1282 = _T_658 ? btb_hcount_42 : 2'h0; // @[Mux.scala 19:72:@2086.4]
  assign _T_1284 = _T_659 ? btb_hcount_43 : 2'h0; // @[Mux.scala 19:72:@2087.4]
  assign _T_1286 = _T_660 ? btb_hcount_44 : 2'h0; // @[Mux.scala 19:72:@2088.4]
  assign _T_1288 = _T_661 ? btb_hcount_45 : 2'h0; // @[Mux.scala 19:72:@2089.4]
  assign _T_1290 = _T_662 ? btb_hcount_46 : 2'h0; // @[Mux.scala 19:72:@2090.4]
  assign _T_1292 = _T_663 ? btb_hcount_47 : 2'h0; // @[Mux.scala 19:72:@2091.4]
  assign _T_1294 = _T_664 ? btb_hcount_48 : 2'h0; // @[Mux.scala 19:72:@2092.4]
  assign _T_1296 = _T_665 ? btb_hcount_49 : 2'h0; // @[Mux.scala 19:72:@2093.4]
  assign _T_1298 = _T_666 ? btb_hcount_50 : 2'h0; // @[Mux.scala 19:72:@2094.4]
  assign _T_1300 = _T_667 ? btb_hcount_51 : 2'h0; // @[Mux.scala 19:72:@2095.4]
  assign _T_1302 = _T_668 ? btb_hcount_52 : 2'h0; // @[Mux.scala 19:72:@2096.4]
  assign _T_1304 = _T_669 ? btb_hcount_53 : 2'h0; // @[Mux.scala 19:72:@2097.4]
  assign _T_1306 = _T_670 ? btb_hcount_54 : 2'h0; // @[Mux.scala 19:72:@2098.4]
  assign _T_1308 = _T_671 ? btb_hcount_55 : 2'h0; // @[Mux.scala 19:72:@2099.4]
  assign _T_1310 = _T_672 ? btb_hcount_56 : 2'h0; // @[Mux.scala 19:72:@2100.4]
  assign _T_1312 = _T_673 ? btb_hcount_57 : 2'h0; // @[Mux.scala 19:72:@2101.4]
  assign _T_1314 = _T_674 ? btb_hcount_58 : 2'h0; // @[Mux.scala 19:72:@2102.4]
  assign _T_1316 = _T_675 ? btb_hcount_59 : 2'h0; // @[Mux.scala 19:72:@2103.4]
  assign _T_1318 = _T_676 ? btb_hcount_60 : 2'h0; // @[Mux.scala 19:72:@2104.4]
  assign _T_1320 = _T_677 ? btb_hcount_61 : 2'h0; // @[Mux.scala 19:72:@2105.4]
  assign _T_1322 = _T_678 ? btb_hcount_62 : 2'h0; // @[Mux.scala 19:72:@2106.4]
  assign _T_1324 = _T_679 ? btb_hcount_63 : 2'h0; // @[Mux.scala 19:72:@2107.4]
  assign _T_1325 = _T_1198 | _T_1200; // @[Mux.scala 19:72:@2108.4]
  assign _T_1326 = _T_1325 | _T_1202; // @[Mux.scala 19:72:@2109.4]
  assign _T_1327 = _T_1326 | _T_1204; // @[Mux.scala 19:72:@2110.4]
  assign _T_1328 = _T_1327 | _T_1206; // @[Mux.scala 19:72:@2111.4]
  assign _T_1329 = _T_1328 | _T_1208; // @[Mux.scala 19:72:@2112.4]
  assign _T_1330 = _T_1329 | _T_1210; // @[Mux.scala 19:72:@2113.4]
  assign _T_1331 = _T_1330 | _T_1212; // @[Mux.scala 19:72:@2114.4]
  assign _T_1332 = _T_1331 | _T_1214; // @[Mux.scala 19:72:@2115.4]
  assign _T_1333 = _T_1332 | _T_1216; // @[Mux.scala 19:72:@2116.4]
  assign _T_1334 = _T_1333 | _T_1218; // @[Mux.scala 19:72:@2117.4]
  assign _T_1335 = _T_1334 | _T_1220; // @[Mux.scala 19:72:@2118.4]
  assign _T_1336 = _T_1335 | _T_1222; // @[Mux.scala 19:72:@2119.4]
  assign _T_1337 = _T_1336 | _T_1224; // @[Mux.scala 19:72:@2120.4]
  assign _T_1338 = _T_1337 | _T_1226; // @[Mux.scala 19:72:@2121.4]
  assign _T_1339 = _T_1338 | _T_1228; // @[Mux.scala 19:72:@2122.4]
  assign _T_1340 = _T_1339 | _T_1230; // @[Mux.scala 19:72:@2123.4]
  assign _T_1341 = _T_1340 | _T_1232; // @[Mux.scala 19:72:@2124.4]
  assign _T_1342 = _T_1341 | _T_1234; // @[Mux.scala 19:72:@2125.4]
  assign _T_1343 = _T_1342 | _T_1236; // @[Mux.scala 19:72:@2126.4]
  assign _T_1344 = _T_1343 | _T_1238; // @[Mux.scala 19:72:@2127.4]
  assign _T_1345 = _T_1344 | _T_1240; // @[Mux.scala 19:72:@2128.4]
  assign _T_1346 = _T_1345 | _T_1242; // @[Mux.scala 19:72:@2129.4]
  assign _T_1347 = _T_1346 | _T_1244; // @[Mux.scala 19:72:@2130.4]
  assign _T_1348 = _T_1347 | _T_1246; // @[Mux.scala 19:72:@2131.4]
  assign _T_1349 = _T_1348 | _T_1248; // @[Mux.scala 19:72:@2132.4]
  assign _T_1350 = _T_1349 | _T_1250; // @[Mux.scala 19:72:@2133.4]
  assign _T_1351 = _T_1350 | _T_1252; // @[Mux.scala 19:72:@2134.4]
  assign _T_1352 = _T_1351 | _T_1254; // @[Mux.scala 19:72:@2135.4]
  assign _T_1353 = _T_1352 | _T_1256; // @[Mux.scala 19:72:@2136.4]
  assign _T_1354 = _T_1353 | _T_1258; // @[Mux.scala 19:72:@2137.4]
  assign _T_1355 = _T_1354 | _T_1260; // @[Mux.scala 19:72:@2138.4]
  assign _T_1356 = _T_1355 | _T_1262; // @[Mux.scala 19:72:@2139.4]
  assign _T_1357 = _T_1356 | _T_1264; // @[Mux.scala 19:72:@2140.4]
  assign _T_1358 = _T_1357 | _T_1266; // @[Mux.scala 19:72:@2141.4]
  assign _T_1359 = _T_1358 | _T_1268; // @[Mux.scala 19:72:@2142.4]
  assign _T_1360 = _T_1359 | _T_1270; // @[Mux.scala 19:72:@2143.4]
  assign _T_1361 = _T_1360 | _T_1272; // @[Mux.scala 19:72:@2144.4]
  assign _T_1362 = _T_1361 | _T_1274; // @[Mux.scala 19:72:@2145.4]
  assign _T_1363 = _T_1362 | _T_1276; // @[Mux.scala 19:72:@2146.4]
  assign _T_1364 = _T_1363 | _T_1278; // @[Mux.scala 19:72:@2147.4]
  assign _T_1365 = _T_1364 | _T_1280; // @[Mux.scala 19:72:@2148.4]
  assign _T_1366 = _T_1365 | _T_1282; // @[Mux.scala 19:72:@2149.4]
  assign _T_1367 = _T_1366 | _T_1284; // @[Mux.scala 19:72:@2150.4]
  assign _T_1368 = _T_1367 | _T_1286; // @[Mux.scala 19:72:@2151.4]
  assign _T_1369 = _T_1368 | _T_1288; // @[Mux.scala 19:72:@2152.4]
  assign _T_1370 = _T_1369 | _T_1290; // @[Mux.scala 19:72:@2153.4]
  assign _T_1371 = _T_1370 | _T_1292; // @[Mux.scala 19:72:@2154.4]
  assign _T_1372 = _T_1371 | _T_1294; // @[Mux.scala 19:72:@2155.4]
  assign _T_1373 = _T_1372 | _T_1296; // @[Mux.scala 19:72:@2156.4]
  assign _T_1374 = _T_1373 | _T_1298; // @[Mux.scala 19:72:@2157.4]
  assign _T_1375 = _T_1374 | _T_1300; // @[Mux.scala 19:72:@2158.4]
  assign _T_1376 = _T_1375 | _T_1302; // @[Mux.scala 19:72:@2159.4]
  assign _T_1377 = _T_1376 | _T_1304; // @[Mux.scala 19:72:@2160.4]
  assign _T_1378 = _T_1377 | _T_1306; // @[Mux.scala 19:72:@2161.4]
  assign _T_1379 = _T_1378 | _T_1308; // @[Mux.scala 19:72:@2162.4]
  assign _T_1380 = _T_1379 | _T_1310; // @[Mux.scala 19:72:@2163.4]
  assign _T_1381 = _T_1380 | _T_1312; // @[Mux.scala 19:72:@2164.4]
  assign _T_1382 = _T_1381 | _T_1314; // @[Mux.scala 19:72:@2165.4]
  assign _T_1383 = _T_1382 | _T_1316; // @[Mux.scala 19:72:@2166.4]
  assign _T_1384 = _T_1383 | _T_1318; // @[Mux.scala 19:72:@2167.4]
  assign _T_1385 = _T_1384 | _T_1320; // @[Mux.scala 19:72:@2168.4]
  assign _T_1386 = _T_1385 | _T_1322; // @[Mux.scala 19:72:@2169.4]
  assign predict_0_hcount = _T_1386 | _T_1324; // @[Mux.scala 19:72:@2170.4]
  assign _T_1391 = predict_0_btype == 2'h1; // @[BTB.scala 80:44:@2174.4]
  assign _T_1393 = predict_0_btype == 2'h2; // @[BTB.scala 69:34:@2175.4]
  assign _T_1394 = predict_0_hcount[1]; // @[BTB.scala 69:65:@2176.4]
  assign _T_1396 = _T_1394 == 1'h0; // @[BTB.scala 69:58:@2177.4]
  assign _T_1397 = _T_1393 & _T_1396; // @[BTB.scala 69:55:@2178.4]
  assign _T_1399 = _T_1397 == 1'h0; // @[BTB.scala 69:26:@2179.4]
  assign _T_1401 = predict_0_lookup != 64'h0; // @[BTB.scala 69:80:@2180.4]
  assign _T_1402 = _T_1399 & _T_1401; // @[BTB.scala 69:70:@2181.4]
  assign if_pc_1 = {_T_152,1'h1,2'h0}; // @[Cat.scala 30:58:@2187.4]
  assign _T_1403 = _T_1402 ? predict_0_jump_tgt : if_pc_1; // @[BTB.scala 70:27:@2182.4]
  assign _T_1410 = btb_pc_0 == if_pc_1; // @[BTB.scala 76:47:@2189.4]
  assign _T_1411 = btb_pc_1 == if_pc_1; // @[BTB.scala 76:47:@2190.4]
  assign _T_1412 = btb_pc_2 == if_pc_1; // @[BTB.scala 76:47:@2191.4]
  assign _T_1413 = btb_pc_3 == if_pc_1; // @[BTB.scala 76:47:@2192.4]
  assign _T_1414 = btb_pc_4 == if_pc_1; // @[BTB.scala 76:47:@2193.4]
  assign _T_1415 = btb_pc_5 == if_pc_1; // @[BTB.scala 76:47:@2194.4]
  assign _T_1416 = btb_pc_6 == if_pc_1; // @[BTB.scala 76:47:@2195.4]
  assign _T_1417 = btb_pc_7 == if_pc_1; // @[BTB.scala 76:47:@2196.4]
  assign _T_1418 = btb_pc_8 == if_pc_1; // @[BTB.scala 76:47:@2197.4]
  assign _T_1419 = btb_pc_9 == if_pc_1; // @[BTB.scala 76:47:@2198.4]
  assign _T_1420 = btb_pc_10 == if_pc_1; // @[BTB.scala 76:47:@2199.4]
  assign _T_1421 = btb_pc_11 == if_pc_1; // @[BTB.scala 76:47:@2200.4]
  assign _T_1422 = btb_pc_12 == if_pc_1; // @[BTB.scala 76:47:@2201.4]
  assign _T_1423 = btb_pc_13 == if_pc_1; // @[BTB.scala 76:47:@2202.4]
  assign _T_1424 = btb_pc_14 == if_pc_1; // @[BTB.scala 76:47:@2203.4]
  assign _T_1425 = btb_pc_15 == if_pc_1; // @[BTB.scala 76:47:@2204.4]
  assign _T_1426 = btb_pc_16 == if_pc_1; // @[BTB.scala 76:47:@2205.4]
  assign _T_1427 = btb_pc_17 == if_pc_1; // @[BTB.scala 76:47:@2206.4]
  assign _T_1428 = btb_pc_18 == if_pc_1; // @[BTB.scala 76:47:@2207.4]
  assign _T_1429 = btb_pc_19 == if_pc_1; // @[BTB.scala 76:47:@2208.4]
  assign _T_1430 = btb_pc_20 == if_pc_1; // @[BTB.scala 76:47:@2209.4]
  assign _T_1431 = btb_pc_21 == if_pc_1; // @[BTB.scala 76:47:@2210.4]
  assign _T_1432 = btb_pc_22 == if_pc_1; // @[BTB.scala 76:47:@2211.4]
  assign _T_1433 = btb_pc_23 == if_pc_1; // @[BTB.scala 76:47:@2212.4]
  assign _T_1434 = btb_pc_24 == if_pc_1; // @[BTB.scala 76:47:@2213.4]
  assign _T_1435 = btb_pc_25 == if_pc_1; // @[BTB.scala 76:47:@2214.4]
  assign _T_1436 = btb_pc_26 == if_pc_1; // @[BTB.scala 76:47:@2215.4]
  assign _T_1437 = btb_pc_27 == if_pc_1; // @[BTB.scala 76:47:@2216.4]
  assign _T_1438 = btb_pc_28 == if_pc_1; // @[BTB.scala 76:47:@2217.4]
  assign _T_1439 = btb_pc_29 == if_pc_1; // @[BTB.scala 76:47:@2218.4]
  assign _T_1440 = btb_pc_30 == if_pc_1; // @[BTB.scala 76:47:@2219.4]
  assign _T_1441 = btb_pc_31 == if_pc_1; // @[BTB.scala 76:47:@2220.4]
  assign _T_1442 = btb_pc_32 == if_pc_1; // @[BTB.scala 76:47:@2221.4]
  assign _T_1443 = btb_pc_33 == if_pc_1; // @[BTB.scala 76:47:@2222.4]
  assign _T_1444 = btb_pc_34 == if_pc_1; // @[BTB.scala 76:47:@2223.4]
  assign _T_1445 = btb_pc_35 == if_pc_1; // @[BTB.scala 76:47:@2224.4]
  assign _T_1446 = btb_pc_36 == if_pc_1; // @[BTB.scala 76:47:@2225.4]
  assign _T_1447 = btb_pc_37 == if_pc_1; // @[BTB.scala 76:47:@2226.4]
  assign _T_1448 = btb_pc_38 == if_pc_1; // @[BTB.scala 76:47:@2227.4]
  assign _T_1449 = btb_pc_39 == if_pc_1; // @[BTB.scala 76:47:@2228.4]
  assign _T_1450 = btb_pc_40 == if_pc_1; // @[BTB.scala 76:47:@2229.4]
  assign _T_1451 = btb_pc_41 == if_pc_1; // @[BTB.scala 76:47:@2230.4]
  assign _T_1452 = btb_pc_42 == if_pc_1; // @[BTB.scala 76:47:@2231.4]
  assign _T_1453 = btb_pc_43 == if_pc_1; // @[BTB.scala 76:47:@2232.4]
  assign _T_1454 = btb_pc_44 == if_pc_1; // @[BTB.scala 76:47:@2233.4]
  assign _T_1455 = btb_pc_45 == if_pc_1; // @[BTB.scala 76:47:@2234.4]
  assign _T_1456 = btb_pc_46 == if_pc_1; // @[BTB.scala 76:47:@2235.4]
  assign _T_1457 = btb_pc_47 == if_pc_1; // @[BTB.scala 76:47:@2236.4]
  assign _T_1458 = btb_pc_48 == if_pc_1; // @[BTB.scala 76:47:@2237.4]
  assign _T_1459 = btb_pc_49 == if_pc_1; // @[BTB.scala 76:47:@2238.4]
  assign _T_1460 = btb_pc_50 == if_pc_1; // @[BTB.scala 76:47:@2239.4]
  assign _T_1461 = btb_pc_51 == if_pc_1; // @[BTB.scala 76:47:@2240.4]
  assign _T_1462 = btb_pc_52 == if_pc_1; // @[BTB.scala 76:47:@2241.4]
  assign _T_1463 = btb_pc_53 == if_pc_1; // @[BTB.scala 76:47:@2242.4]
  assign _T_1464 = btb_pc_54 == if_pc_1; // @[BTB.scala 76:47:@2243.4]
  assign _T_1465 = btb_pc_55 == if_pc_1; // @[BTB.scala 76:47:@2244.4]
  assign _T_1466 = btb_pc_56 == if_pc_1; // @[BTB.scala 76:47:@2245.4]
  assign _T_1467 = btb_pc_57 == if_pc_1; // @[BTB.scala 76:47:@2246.4]
  assign _T_1468 = btb_pc_58 == if_pc_1; // @[BTB.scala 76:47:@2247.4]
  assign _T_1469 = btb_pc_59 == if_pc_1; // @[BTB.scala 76:47:@2248.4]
  assign _T_1470 = btb_pc_60 == if_pc_1; // @[BTB.scala 76:47:@2249.4]
  assign _T_1471 = btb_pc_61 == if_pc_1; // @[BTB.scala 76:47:@2250.4]
  assign _T_1472 = btb_pc_62 == if_pc_1; // @[BTB.scala 76:47:@2251.4]
  assign _T_1473 = btb_pc_63 == if_pc_1; // @[BTB.scala 76:47:@2252.4]
  assign _T_1550 = {_T_1417,_T_1416,_T_1415,_T_1414,_T_1413,_T_1412,_T_1411,_T_1410}; // @[BTB.scala 76:62:@2324.4]
  assign _T_1558 = {_T_1425,_T_1424,_T_1423,_T_1422,_T_1421,_T_1420,_T_1419,_T_1418,_T_1550}; // @[BTB.scala 76:62:@2332.4]
  assign _T_1565 = {_T_1433,_T_1432,_T_1431,_T_1430,_T_1429,_T_1428,_T_1427,_T_1426}; // @[BTB.scala 76:62:@2339.4]
  assign _T_1574 = {_T_1441,_T_1440,_T_1439,_T_1438,_T_1437,_T_1436,_T_1435,_T_1434,_T_1565,_T_1558}; // @[BTB.scala 76:62:@2348.4]
  assign _T_1581 = {_T_1449,_T_1448,_T_1447,_T_1446,_T_1445,_T_1444,_T_1443,_T_1442}; // @[BTB.scala 76:62:@2355.4]
  assign _T_1589 = {_T_1457,_T_1456,_T_1455,_T_1454,_T_1453,_T_1452,_T_1451,_T_1450,_T_1581}; // @[BTB.scala 76:62:@2363.4]
  assign _T_1596 = {_T_1465,_T_1464,_T_1463,_T_1462,_T_1461,_T_1460,_T_1459,_T_1458}; // @[BTB.scala 76:62:@2370.4]
  assign _T_1605 = {_T_1473,_T_1472,_T_1471,_T_1470,_T_1469,_T_1468,_T_1467,_T_1466,_T_1596,_T_1589}; // @[BTB.scala 76:62:@2379.4]
  assign _T_1606 = {_T_1605,_T_1574}; // @[BTB.scala 76:62:@2380.4]
  assign predict_1_lookup = _T_1606 & _T_614; // @[BTB.scala 76:69:@2573.4]
  assign _T_1869 = predict_1_lookup[0]; // @[Mux.scala 21:36:@2575.4]
  assign _T_1870 = predict_1_lookup[1]; // @[Mux.scala 21:36:@2576.4]
  assign _T_1871 = predict_1_lookup[2]; // @[Mux.scala 21:36:@2577.4]
  assign _T_1872 = predict_1_lookup[3]; // @[Mux.scala 21:36:@2578.4]
  assign _T_1873 = predict_1_lookup[4]; // @[Mux.scala 21:36:@2579.4]
  assign _T_1874 = predict_1_lookup[5]; // @[Mux.scala 21:36:@2580.4]
  assign _T_1875 = predict_1_lookup[6]; // @[Mux.scala 21:36:@2581.4]
  assign _T_1876 = predict_1_lookup[7]; // @[Mux.scala 21:36:@2582.4]
  assign _T_1877 = predict_1_lookup[8]; // @[Mux.scala 21:36:@2583.4]
  assign _T_1878 = predict_1_lookup[9]; // @[Mux.scala 21:36:@2584.4]
  assign _T_1879 = predict_1_lookup[10]; // @[Mux.scala 21:36:@2585.4]
  assign _T_1880 = predict_1_lookup[11]; // @[Mux.scala 21:36:@2586.4]
  assign _T_1881 = predict_1_lookup[12]; // @[Mux.scala 21:36:@2587.4]
  assign _T_1882 = predict_1_lookup[13]; // @[Mux.scala 21:36:@2588.4]
  assign _T_1883 = predict_1_lookup[14]; // @[Mux.scala 21:36:@2589.4]
  assign _T_1884 = predict_1_lookup[15]; // @[Mux.scala 21:36:@2590.4]
  assign _T_1885 = predict_1_lookup[16]; // @[Mux.scala 21:36:@2591.4]
  assign _T_1886 = predict_1_lookup[17]; // @[Mux.scala 21:36:@2592.4]
  assign _T_1887 = predict_1_lookup[18]; // @[Mux.scala 21:36:@2593.4]
  assign _T_1888 = predict_1_lookup[19]; // @[Mux.scala 21:36:@2594.4]
  assign _T_1889 = predict_1_lookup[20]; // @[Mux.scala 21:36:@2595.4]
  assign _T_1890 = predict_1_lookup[21]; // @[Mux.scala 21:36:@2596.4]
  assign _T_1891 = predict_1_lookup[22]; // @[Mux.scala 21:36:@2597.4]
  assign _T_1892 = predict_1_lookup[23]; // @[Mux.scala 21:36:@2598.4]
  assign _T_1893 = predict_1_lookup[24]; // @[Mux.scala 21:36:@2599.4]
  assign _T_1894 = predict_1_lookup[25]; // @[Mux.scala 21:36:@2600.4]
  assign _T_1895 = predict_1_lookup[26]; // @[Mux.scala 21:36:@2601.4]
  assign _T_1896 = predict_1_lookup[27]; // @[Mux.scala 21:36:@2602.4]
  assign _T_1897 = predict_1_lookup[28]; // @[Mux.scala 21:36:@2603.4]
  assign _T_1898 = predict_1_lookup[29]; // @[Mux.scala 21:36:@2604.4]
  assign _T_1899 = predict_1_lookup[30]; // @[Mux.scala 21:36:@2605.4]
  assign _T_1900 = predict_1_lookup[31]; // @[Mux.scala 21:36:@2606.4]
  assign _T_1901 = predict_1_lookup[32]; // @[Mux.scala 21:36:@2607.4]
  assign _T_1902 = predict_1_lookup[33]; // @[Mux.scala 21:36:@2608.4]
  assign _T_1903 = predict_1_lookup[34]; // @[Mux.scala 21:36:@2609.4]
  assign _T_1904 = predict_1_lookup[35]; // @[Mux.scala 21:36:@2610.4]
  assign _T_1905 = predict_1_lookup[36]; // @[Mux.scala 21:36:@2611.4]
  assign _T_1906 = predict_1_lookup[37]; // @[Mux.scala 21:36:@2612.4]
  assign _T_1907 = predict_1_lookup[38]; // @[Mux.scala 21:36:@2613.4]
  assign _T_1908 = predict_1_lookup[39]; // @[Mux.scala 21:36:@2614.4]
  assign _T_1909 = predict_1_lookup[40]; // @[Mux.scala 21:36:@2615.4]
  assign _T_1910 = predict_1_lookup[41]; // @[Mux.scala 21:36:@2616.4]
  assign _T_1911 = predict_1_lookup[42]; // @[Mux.scala 21:36:@2617.4]
  assign _T_1912 = predict_1_lookup[43]; // @[Mux.scala 21:36:@2618.4]
  assign _T_1913 = predict_1_lookup[44]; // @[Mux.scala 21:36:@2619.4]
  assign _T_1914 = predict_1_lookup[45]; // @[Mux.scala 21:36:@2620.4]
  assign _T_1915 = predict_1_lookup[46]; // @[Mux.scala 21:36:@2621.4]
  assign _T_1916 = predict_1_lookup[47]; // @[Mux.scala 21:36:@2622.4]
  assign _T_1917 = predict_1_lookup[48]; // @[Mux.scala 21:36:@2623.4]
  assign _T_1918 = predict_1_lookup[49]; // @[Mux.scala 21:36:@2624.4]
  assign _T_1919 = predict_1_lookup[50]; // @[Mux.scala 21:36:@2625.4]
  assign _T_1920 = predict_1_lookup[51]; // @[Mux.scala 21:36:@2626.4]
  assign _T_1921 = predict_1_lookup[52]; // @[Mux.scala 21:36:@2627.4]
  assign _T_1922 = predict_1_lookup[53]; // @[Mux.scala 21:36:@2628.4]
  assign _T_1923 = predict_1_lookup[54]; // @[Mux.scala 21:36:@2629.4]
  assign _T_1924 = predict_1_lookup[55]; // @[Mux.scala 21:36:@2630.4]
  assign _T_1925 = predict_1_lookup[56]; // @[Mux.scala 21:36:@2631.4]
  assign _T_1926 = predict_1_lookup[57]; // @[Mux.scala 21:36:@2632.4]
  assign _T_1927 = predict_1_lookup[58]; // @[Mux.scala 21:36:@2633.4]
  assign _T_1928 = predict_1_lookup[59]; // @[Mux.scala 21:36:@2634.4]
  assign _T_1929 = predict_1_lookup[60]; // @[Mux.scala 21:36:@2635.4]
  assign _T_1930 = predict_1_lookup[61]; // @[Mux.scala 21:36:@2636.4]
  assign _T_1931 = predict_1_lookup[62]; // @[Mux.scala 21:36:@2637.4]
  assign _T_1932 = predict_1_lookup[63]; // @[Mux.scala 21:36:@2638.4]
  assign _T_1935 = _T_1869 ? btb_target_0 : 32'h0; // @[Mux.scala 19:72:@2639.4]
  assign _T_1937 = _T_1870 ? btb_target_1 : 32'h0; // @[Mux.scala 19:72:@2640.4]
  assign _T_1939 = _T_1871 ? btb_target_2 : 32'h0; // @[Mux.scala 19:72:@2641.4]
  assign _T_1941 = _T_1872 ? btb_target_3 : 32'h0; // @[Mux.scala 19:72:@2642.4]
  assign _T_1943 = _T_1873 ? btb_target_4 : 32'h0; // @[Mux.scala 19:72:@2643.4]
  assign _T_1945 = _T_1874 ? btb_target_5 : 32'h0; // @[Mux.scala 19:72:@2644.4]
  assign _T_1947 = _T_1875 ? btb_target_6 : 32'h0; // @[Mux.scala 19:72:@2645.4]
  assign _T_1949 = _T_1876 ? btb_target_7 : 32'h0; // @[Mux.scala 19:72:@2646.4]
  assign _T_1951 = _T_1877 ? btb_target_8 : 32'h0; // @[Mux.scala 19:72:@2647.4]
  assign _T_1953 = _T_1878 ? btb_target_9 : 32'h0; // @[Mux.scala 19:72:@2648.4]
  assign _T_1955 = _T_1879 ? btb_target_10 : 32'h0; // @[Mux.scala 19:72:@2649.4]
  assign _T_1957 = _T_1880 ? btb_target_11 : 32'h0; // @[Mux.scala 19:72:@2650.4]
  assign _T_1959 = _T_1881 ? btb_target_12 : 32'h0; // @[Mux.scala 19:72:@2651.4]
  assign _T_1961 = _T_1882 ? btb_target_13 : 32'h0; // @[Mux.scala 19:72:@2652.4]
  assign _T_1963 = _T_1883 ? btb_target_14 : 32'h0; // @[Mux.scala 19:72:@2653.4]
  assign _T_1965 = _T_1884 ? btb_target_15 : 32'h0; // @[Mux.scala 19:72:@2654.4]
  assign _T_1967 = _T_1885 ? btb_target_16 : 32'h0; // @[Mux.scala 19:72:@2655.4]
  assign _T_1969 = _T_1886 ? btb_target_17 : 32'h0; // @[Mux.scala 19:72:@2656.4]
  assign _T_1971 = _T_1887 ? btb_target_18 : 32'h0; // @[Mux.scala 19:72:@2657.4]
  assign _T_1973 = _T_1888 ? btb_target_19 : 32'h0; // @[Mux.scala 19:72:@2658.4]
  assign _T_1975 = _T_1889 ? btb_target_20 : 32'h0; // @[Mux.scala 19:72:@2659.4]
  assign _T_1977 = _T_1890 ? btb_target_21 : 32'h0; // @[Mux.scala 19:72:@2660.4]
  assign _T_1979 = _T_1891 ? btb_target_22 : 32'h0; // @[Mux.scala 19:72:@2661.4]
  assign _T_1981 = _T_1892 ? btb_target_23 : 32'h0; // @[Mux.scala 19:72:@2662.4]
  assign _T_1983 = _T_1893 ? btb_target_24 : 32'h0; // @[Mux.scala 19:72:@2663.4]
  assign _T_1985 = _T_1894 ? btb_target_25 : 32'h0; // @[Mux.scala 19:72:@2664.4]
  assign _T_1987 = _T_1895 ? btb_target_26 : 32'h0; // @[Mux.scala 19:72:@2665.4]
  assign _T_1989 = _T_1896 ? btb_target_27 : 32'h0; // @[Mux.scala 19:72:@2666.4]
  assign _T_1991 = _T_1897 ? btb_target_28 : 32'h0; // @[Mux.scala 19:72:@2667.4]
  assign _T_1993 = _T_1898 ? btb_target_29 : 32'h0; // @[Mux.scala 19:72:@2668.4]
  assign _T_1995 = _T_1899 ? btb_target_30 : 32'h0; // @[Mux.scala 19:72:@2669.4]
  assign _T_1997 = _T_1900 ? btb_target_31 : 32'h0; // @[Mux.scala 19:72:@2670.4]
  assign _T_1999 = _T_1901 ? btb_target_32 : 32'h0; // @[Mux.scala 19:72:@2671.4]
  assign _T_2001 = _T_1902 ? btb_target_33 : 32'h0; // @[Mux.scala 19:72:@2672.4]
  assign _T_2003 = _T_1903 ? btb_target_34 : 32'h0; // @[Mux.scala 19:72:@2673.4]
  assign _T_2005 = _T_1904 ? btb_target_35 : 32'h0; // @[Mux.scala 19:72:@2674.4]
  assign _T_2007 = _T_1905 ? btb_target_36 : 32'h0; // @[Mux.scala 19:72:@2675.4]
  assign _T_2009 = _T_1906 ? btb_target_37 : 32'h0; // @[Mux.scala 19:72:@2676.4]
  assign _T_2011 = _T_1907 ? btb_target_38 : 32'h0; // @[Mux.scala 19:72:@2677.4]
  assign _T_2013 = _T_1908 ? btb_target_39 : 32'h0; // @[Mux.scala 19:72:@2678.4]
  assign _T_2015 = _T_1909 ? btb_target_40 : 32'h0; // @[Mux.scala 19:72:@2679.4]
  assign _T_2017 = _T_1910 ? btb_target_41 : 32'h0; // @[Mux.scala 19:72:@2680.4]
  assign _T_2019 = _T_1911 ? btb_target_42 : 32'h0; // @[Mux.scala 19:72:@2681.4]
  assign _T_2021 = _T_1912 ? btb_target_43 : 32'h0; // @[Mux.scala 19:72:@2682.4]
  assign _T_2023 = _T_1913 ? btb_target_44 : 32'h0; // @[Mux.scala 19:72:@2683.4]
  assign _T_2025 = _T_1914 ? btb_target_45 : 32'h0; // @[Mux.scala 19:72:@2684.4]
  assign _T_2027 = _T_1915 ? btb_target_46 : 32'h0; // @[Mux.scala 19:72:@2685.4]
  assign _T_2029 = _T_1916 ? btb_target_47 : 32'h0; // @[Mux.scala 19:72:@2686.4]
  assign _T_2031 = _T_1917 ? btb_target_48 : 32'h0; // @[Mux.scala 19:72:@2687.4]
  assign _T_2033 = _T_1918 ? btb_target_49 : 32'h0; // @[Mux.scala 19:72:@2688.4]
  assign _T_2035 = _T_1919 ? btb_target_50 : 32'h0; // @[Mux.scala 19:72:@2689.4]
  assign _T_2037 = _T_1920 ? btb_target_51 : 32'h0; // @[Mux.scala 19:72:@2690.4]
  assign _T_2039 = _T_1921 ? btb_target_52 : 32'h0; // @[Mux.scala 19:72:@2691.4]
  assign _T_2041 = _T_1922 ? btb_target_53 : 32'h0; // @[Mux.scala 19:72:@2692.4]
  assign _T_2043 = _T_1923 ? btb_target_54 : 32'h0; // @[Mux.scala 19:72:@2693.4]
  assign _T_2045 = _T_1924 ? btb_target_55 : 32'h0; // @[Mux.scala 19:72:@2694.4]
  assign _T_2047 = _T_1925 ? btb_target_56 : 32'h0; // @[Mux.scala 19:72:@2695.4]
  assign _T_2049 = _T_1926 ? btb_target_57 : 32'h0; // @[Mux.scala 19:72:@2696.4]
  assign _T_2051 = _T_1927 ? btb_target_58 : 32'h0; // @[Mux.scala 19:72:@2697.4]
  assign _T_2053 = _T_1928 ? btb_target_59 : 32'h0; // @[Mux.scala 19:72:@2698.4]
  assign _T_2055 = _T_1929 ? btb_target_60 : 32'h0; // @[Mux.scala 19:72:@2699.4]
  assign _T_2057 = _T_1930 ? btb_target_61 : 32'h0; // @[Mux.scala 19:72:@2700.4]
  assign _T_2059 = _T_1931 ? btb_target_62 : 32'h0; // @[Mux.scala 19:72:@2701.4]
  assign _T_2061 = _T_1932 ? btb_target_63 : 32'h0; // @[Mux.scala 19:72:@2702.4]
  assign _T_2062 = _T_1935 | _T_1937; // @[Mux.scala 19:72:@2703.4]
  assign _T_2063 = _T_2062 | _T_1939; // @[Mux.scala 19:72:@2704.4]
  assign _T_2064 = _T_2063 | _T_1941; // @[Mux.scala 19:72:@2705.4]
  assign _T_2065 = _T_2064 | _T_1943; // @[Mux.scala 19:72:@2706.4]
  assign _T_2066 = _T_2065 | _T_1945; // @[Mux.scala 19:72:@2707.4]
  assign _T_2067 = _T_2066 | _T_1947; // @[Mux.scala 19:72:@2708.4]
  assign _T_2068 = _T_2067 | _T_1949; // @[Mux.scala 19:72:@2709.4]
  assign _T_2069 = _T_2068 | _T_1951; // @[Mux.scala 19:72:@2710.4]
  assign _T_2070 = _T_2069 | _T_1953; // @[Mux.scala 19:72:@2711.4]
  assign _T_2071 = _T_2070 | _T_1955; // @[Mux.scala 19:72:@2712.4]
  assign _T_2072 = _T_2071 | _T_1957; // @[Mux.scala 19:72:@2713.4]
  assign _T_2073 = _T_2072 | _T_1959; // @[Mux.scala 19:72:@2714.4]
  assign _T_2074 = _T_2073 | _T_1961; // @[Mux.scala 19:72:@2715.4]
  assign _T_2075 = _T_2074 | _T_1963; // @[Mux.scala 19:72:@2716.4]
  assign _T_2076 = _T_2075 | _T_1965; // @[Mux.scala 19:72:@2717.4]
  assign _T_2077 = _T_2076 | _T_1967; // @[Mux.scala 19:72:@2718.4]
  assign _T_2078 = _T_2077 | _T_1969; // @[Mux.scala 19:72:@2719.4]
  assign _T_2079 = _T_2078 | _T_1971; // @[Mux.scala 19:72:@2720.4]
  assign _T_2080 = _T_2079 | _T_1973; // @[Mux.scala 19:72:@2721.4]
  assign _T_2081 = _T_2080 | _T_1975; // @[Mux.scala 19:72:@2722.4]
  assign _T_2082 = _T_2081 | _T_1977; // @[Mux.scala 19:72:@2723.4]
  assign _T_2083 = _T_2082 | _T_1979; // @[Mux.scala 19:72:@2724.4]
  assign _T_2084 = _T_2083 | _T_1981; // @[Mux.scala 19:72:@2725.4]
  assign _T_2085 = _T_2084 | _T_1983; // @[Mux.scala 19:72:@2726.4]
  assign _T_2086 = _T_2085 | _T_1985; // @[Mux.scala 19:72:@2727.4]
  assign _T_2087 = _T_2086 | _T_1987; // @[Mux.scala 19:72:@2728.4]
  assign _T_2088 = _T_2087 | _T_1989; // @[Mux.scala 19:72:@2729.4]
  assign _T_2089 = _T_2088 | _T_1991; // @[Mux.scala 19:72:@2730.4]
  assign _T_2090 = _T_2089 | _T_1993; // @[Mux.scala 19:72:@2731.4]
  assign _T_2091 = _T_2090 | _T_1995; // @[Mux.scala 19:72:@2732.4]
  assign _T_2092 = _T_2091 | _T_1997; // @[Mux.scala 19:72:@2733.4]
  assign _T_2093 = _T_2092 | _T_1999; // @[Mux.scala 19:72:@2734.4]
  assign _T_2094 = _T_2093 | _T_2001; // @[Mux.scala 19:72:@2735.4]
  assign _T_2095 = _T_2094 | _T_2003; // @[Mux.scala 19:72:@2736.4]
  assign _T_2096 = _T_2095 | _T_2005; // @[Mux.scala 19:72:@2737.4]
  assign _T_2097 = _T_2096 | _T_2007; // @[Mux.scala 19:72:@2738.4]
  assign _T_2098 = _T_2097 | _T_2009; // @[Mux.scala 19:72:@2739.4]
  assign _T_2099 = _T_2098 | _T_2011; // @[Mux.scala 19:72:@2740.4]
  assign _T_2100 = _T_2099 | _T_2013; // @[Mux.scala 19:72:@2741.4]
  assign _T_2101 = _T_2100 | _T_2015; // @[Mux.scala 19:72:@2742.4]
  assign _T_2102 = _T_2101 | _T_2017; // @[Mux.scala 19:72:@2743.4]
  assign _T_2103 = _T_2102 | _T_2019; // @[Mux.scala 19:72:@2744.4]
  assign _T_2104 = _T_2103 | _T_2021; // @[Mux.scala 19:72:@2745.4]
  assign _T_2105 = _T_2104 | _T_2023; // @[Mux.scala 19:72:@2746.4]
  assign _T_2106 = _T_2105 | _T_2025; // @[Mux.scala 19:72:@2747.4]
  assign _T_2107 = _T_2106 | _T_2027; // @[Mux.scala 19:72:@2748.4]
  assign _T_2108 = _T_2107 | _T_2029; // @[Mux.scala 19:72:@2749.4]
  assign _T_2109 = _T_2108 | _T_2031; // @[Mux.scala 19:72:@2750.4]
  assign _T_2110 = _T_2109 | _T_2033; // @[Mux.scala 19:72:@2751.4]
  assign _T_2111 = _T_2110 | _T_2035; // @[Mux.scala 19:72:@2752.4]
  assign _T_2112 = _T_2111 | _T_2037; // @[Mux.scala 19:72:@2753.4]
  assign _T_2113 = _T_2112 | _T_2039; // @[Mux.scala 19:72:@2754.4]
  assign _T_2114 = _T_2113 | _T_2041; // @[Mux.scala 19:72:@2755.4]
  assign _T_2115 = _T_2114 | _T_2043; // @[Mux.scala 19:72:@2756.4]
  assign _T_2116 = _T_2115 | _T_2045; // @[Mux.scala 19:72:@2757.4]
  assign _T_2117 = _T_2116 | _T_2047; // @[Mux.scala 19:72:@2758.4]
  assign _T_2118 = _T_2117 | _T_2049; // @[Mux.scala 19:72:@2759.4]
  assign _T_2119 = _T_2118 | _T_2051; // @[Mux.scala 19:72:@2760.4]
  assign _T_2120 = _T_2119 | _T_2053; // @[Mux.scala 19:72:@2761.4]
  assign _T_2121 = _T_2120 | _T_2055; // @[Mux.scala 19:72:@2762.4]
  assign _T_2122 = _T_2121 | _T_2057; // @[Mux.scala 19:72:@2763.4]
  assign _T_2123 = _T_2122 | _T_2059; // @[Mux.scala 19:72:@2764.4]
  assign predict_1_jump_tgt = _T_2123 | _T_2061; // @[Mux.scala 19:72:@2765.4]
  assign _T_2193 = _T_1869 ? btb_btype_0 : 2'h0; // @[Mux.scala 19:72:@2833.4]
  assign _T_2195 = _T_1870 ? btb_btype_1 : 2'h0; // @[Mux.scala 19:72:@2834.4]
  assign _T_2197 = _T_1871 ? btb_btype_2 : 2'h0; // @[Mux.scala 19:72:@2835.4]
  assign _T_2199 = _T_1872 ? btb_btype_3 : 2'h0; // @[Mux.scala 19:72:@2836.4]
  assign _T_2201 = _T_1873 ? btb_btype_4 : 2'h0; // @[Mux.scala 19:72:@2837.4]
  assign _T_2203 = _T_1874 ? btb_btype_5 : 2'h0; // @[Mux.scala 19:72:@2838.4]
  assign _T_2205 = _T_1875 ? btb_btype_6 : 2'h0; // @[Mux.scala 19:72:@2839.4]
  assign _T_2207 = _T_1876 ? btb_btype_7 : 2'h0; // @[Mux.scala 19:72:@2840.4]
  assign _T_2209 = _T_1877 ? btb_btype_8 : 2'h0; // @[Mux.scala 19:72:@2841.4]
  assign _T_2211 = _T_1878 ? btb_btype_9 : 2'h0; // @[Mux.scala 19:72:@2842.4]
  assign _T_2213 = _T_1879 ? btb_btype_10 : 2'h0; // @[Mux.scala 19:72:@2843.4]
  assign _T_2215 = _T_1880 ? btb_btype_11 : 2'h0; // @[Mux.scala 19:72:@2844.4]
  assign _T_2217 = _T_1881 ? btb_btype_12 : 2'h0; // @[Mux.scala 19:72:@2845.4]
  assign _T_2219 = _T_1882 ? btb_btype_13 : 2'h0; // @[Mux.scala 19:72:@2846.4]
  assign _T_2221 = _T_1883 ? btb_btype_14 : 2'h0; // @[Mux.scala 19:72:@2847.4]
  assign _T_2223 = _T_1884 ? btb_btype_15 : 2'h0; // @[Mux.scala 19:72:@2848.4]
  assign _T_2225 = _T_1885 ? btb_btype_16 : 2'h0; // @[Mux.scala 19:72:@2849.4]
  assign _T_2227 = _T_1886 ? btb_btype_17 : 2'h0; // @[Mux.scala 19:72:@2850.4]
  assign _T_2229 = _T_1887 ? btb_btype_18 : 2'h0; // @[Mux.scala 19:72:@2851.4]
  assign _T_2231 = _T_1888 ? btb_btype_19 : 2'h0; // @[Mux.scala 19:72:@2852.4]
  assign _T_2233 = _T_1889 ? btb_btype_20 : 2'h0; // @[Mux.scala 19:72:@2853.4]
  assign _T_2235 = _T_1890 ? btb_btype_21 : 2'h0; // @[Mux.scala 19:72:@2854.4]
  assign _T_2237 = _T_1891 ? btb_btype_22 : 2'h0; // @[Mux.scala 19:72:@2855.4]
  assign _T_2239 = _T_1892 ? btb_btype_23 : 2'h0; // @[Mux.scala 19:72:@2856.4]
  assign _T_2241 = _T_1893 ? btb_btype_24 : 2'h0; // @[Mux.scala 19:72:@2857.4]
  assign _T_2243 = _T_1894 ? btb_btype_25 : 2'h0; // @[Mux.scala 19:72:@2858.4]
  assign _T_2245 = _T_1895 ? btb_btype_26 : 2'h0; // @[Mux.scala 19:72:@2859.4]
  assign _T_2247 = _T_1896 ? btb_btype_27 : 2'h0; // @[Mux.scala 19:72:@2860.4]
  assign _T_2249 = _T_1897 ? btb_btype_28 : 2'h0; // @[Mux.scala 19:72:@2861.4]
  assign _T_2251 = _T_1898 ? btb_btype_29 : 2'h0; // @[Mux.scala 19:72:@2862.4]
  assign _T_2253 = _T_1899 ? btb_btype_30 : 2'h0; // @[Mux.scala 19:72:@2863.4]
  assign _T_2255 = _T_1900 ? btb_btype_31 : 2'h0; // @[Mux.scala 19:72:@2864.4]
  assign _T_2257 = _T_1901 ? btb_btype_32 : 2'h0; // @[Mux.scala 19:72:@2865.4]
  assign _T_2259 = _T_1902 ? btb_btype_33 : 2'h0; // @[Mux.scala 19:72:@2866.4]
  assign _T_2261 = _T_1903 ? btb_btype_34 : 2'h0; // @[Mux.scala 19:72:@2867.4]
  assign _T_2263 = _T_1904 ? btb_btype_35 : 2'h0; // @[Mux.scala 19:72:@2868.4]
  assign _T_2265 = _T_1905 ? btb_btype_36 : 2'h0; // @[Mux.scala 19:72:@2869.4]
  assign _T_2267 = _T_1906 ? btb_btype_37 : 2'h0; // @[Mux.scala 19:72:@2870.4]
  assign _T_2269 = _T_1907 ? btb_btype_38 : 2'h0; // @[Mux.scala 19:72:@2871.4]
  assign _T_2271 = _T_1908 ? btb_btype_39 : 2'h0; // @[Mux.scala 19:72:@2872.4]
  assign _T_2273 = _T_1909 ? btb_btype_40 : 2'h0; // @[Mux.scala 19:72:@2873.4]
  assign _T_2275 = _T_1910 ? btb_btype_41 : 2'h0; // @[Mux.scala 19:72:@2874.4]
  assign _T_2277 = _T_1911 ? btb_btype_42 : 2'h0; // @[Mux.scala 19:72:@2875.4]
  assign _T_2279 = _T_1912 ? btb_btype_43 : 2'h0; // @[Mux.scala 19:72:@2876.4]
  assign _T_2281 = _T_1913 ? btb_btype_44 : 2'h0; // @[Mux.scala 19:72:@2877.4]
  assign _T_2283 = _T_1914 ? btb_btype_45 : 2'h0; // @[Mux.scala 19:72:@2878.4]
  assign _T_2285 = _T_1915 ? btb_btype_46 : 2'h0; // @[Mux.scala 19:72:@2879.4]
  assign _T_2287 = _T_1916 ? btb_btype_47 : 2'h0; // @[Mux.scala 19:72:@2880.4]
  assign _T_2289 = _T_1917 ? btb_btype_48 : 2'h0; // @[Mux.scala 19:72:@2881.4]
  assign _T_2291 = _T_1918 ? btb_btype_49 : 2'h0; // @[Mux.scala 19:72:@2882.4]
  assign _T_2293 = _T_1919 ? btb_btype_50 : 2'h0; // @[Mux.scala 19:72:@2883.4]
  assign _T_2295 = _T_1920 ? btb_btype_51 : 2'h0; // @[Mux.scala 19:72:@2884.4]
  assign _T_2297 = _T_1921 ? btb_btype_52 : 2'h0; // @[Mux.scala 19:72:@2885.4]
  assign _T_2299 = _T_1922 ? btb_btype_53 : 2'h0; // @[Mux.scala 19:72:@2886.4]
  assign _T_2301 = _T_1923 ? btb_btype_54 : 2'h0; // @[Mux.scala 19:72:@2887.4]
  assign _T_2303 = _T_1924 ? btb_btype_55 : 2'h0; // @[Mux.scala 19:72:@2888.4]
  assign _T_2305 = _T_1925 ? btb_btype_56 : 2'h0; // @[Mux.scala 19:72:@2889.4]
  assign _T_2307 = _T_1926 ? btb_btype_57 : 2'h0; // @[Mux.scala 19:72:@2890.4]
  assign _T_2309 = _T_1927 ? btb_btype_58 : 2'h0; // @[Mux.scala 19:72:@2891.4]
  assign _T_2311 = _T_1928 ? btb_btype_59 : 2'h0; // @[Mux.scala 19:72:@2892.4]
  assign _T_2313 = _T_1929 ? btb_btype_60 : 2'h0; // @[Mux.scala 19:72:@2893.4]
  assign _T_2315 = _T_1930 ? btb_btype_61 : 2'h0; // @[Mux.scala 19:72:@2894.4]
  assign _T_2317 = _T_1931 ? btb_btype_62 : 2'h0; // @[Mux.scala 19:72:@2895.4]
  assign _T_2319 = _T_1932 ? btb_btype_63 : 2'h0; // @[Mux.scala 19:72:@2896.4]
  assign _T_2320 = _T_2193 | _T_2195; // @[Mux.scala 19:72:@2897.4]
  assign _T_2321 = _T_2320 | _T_2197; // @[Mux.scala 19:72:@2898.4]
  assign _T_2322 = _T_2321 | _T_2199; // @[Mux.scala 19:72:@2899.4]
  assign _T_2323 = _T_2322 | _T_2201; // @[Mux.scala 19:72:@2900.4]
  assign _T_2324 = _T_2323 | _T_2203; // @[Mux.scala 19:72:@2901.4]
  assign _T_2325 = _T_2324 | _T_2205; // @[Mux.scala 19:72:@2902.4]
  assign _T_2326 = _T_2325 | _T_2207; // @[Mux.scala 19:72:@2903.4]
  assign _T_2327 = _T_2326 | _T_2209; // @[Mux.scala 19:72:@2904.4]
  assign _T_2328 = _T_2327 | _T_2211; // @[Mux.scala 19:72:@2905.4]
  assign _T_2329 = _T_2328 | _T_2213; // @[Mux.scala 19:72:@2906.4]
  assign _T_2330 = _T_2329 | _T_2215; // @[Mux.scala 19:72:@2907.4]
  assign _T_2331 = _T_2330 | _T_2217; // @[Mux.scala 19:72:@2908.4]
  assign _T_2332 = _T_2331 | _T_2219; // @[Mux.scala 19:72:@2909.4]
  assign _T_2333 = _T_2332 | _T_2221; // @[Mux.scala 19:72:@2910.4]
  assign _T_2334 = _T_2333 | _T_2223; // @[Mux.scala 19:72:@2911.4]
  assign _T_2335 = _T_2334 | _T_2225; // @[Mux.scala 19:72:@2912.4]
  assign _T_2336 = _T_2335 | _T_2227; // @[Mux.scala 19:72:@2913.4]
  assign _T_2337 = _T_2336 | _T_2229; // @[Mux.scala 19:72:@2914.4]
  assign _T_2338 = _T_2337 | _T_2231; // @[Mux.scala 19:72:@2915.4]
  assign _T_2339 = _T_2338 | _T_2233; // @[Mux.scala 19:72:@2916.4]
  assign _T_2340 = _T_2339 | _T_2235; // @[Mux.scala 19:72:@2917.4]
  assign _T_2341 = _T_2340 | _T_2237; // @[Mux.scala 19:72:@2918.4]
  assign _T_2342 = _T_2341 | _T_2239; // @[Mux.scala 19:72:@2919.4]
  assign _T_2343 = _T_2342 | _T_2241; // @[Mux.scala 19:72:@2920.4]
  assign _T_2344 = _T_2343 | _T_2243; // @[Mux.scala 19:72:@2921.4]
  assign _T_2345 = _T_2344 | _T_2245; // @[Mux.scala 19:72:@2922.4]
  assign _T_2346 = _T_2345 | _T_2247; // @[Mux.scala 19:72:@2923.4]
  assign _T_2347 = _T_2346 | _T_2249; // @[Mux.scala 19:72:@2924.4]
  assign _T_2348 = _T_2347 | _T_2251; // @[Mux.scala 19:72:@2925.4]
  assign _T_2349 = _T_2348 | _T_2253; // @[Mux.scala 19:72:@2926.4]
  assign _T_2350 = _T_2349 | _T_2255; // @[Mux.scala 19:72:@2927.4]
  assign _T_2351 = _T_2350 | _T_2257; // @[Mux.scala 19:72:@2928.4]
  assign _T_2352 = _T_2351 | _T_2259; // @[Mux.scala 19:72:@2929.4]
  assign _T_2353 = _T_2352 | _T_2261; // @[Mux.scala 19:72:@2930.4]
  assign _T_2354 = _T_2353 | _T_2263; // @[Mux.scala 19:72:@2931.4]
  assign _T_2355 = _T_2354 | _T_2265; // @[Mux.scala 19:72:@2932.4]
  assign _T_2356 = _T_2355 | _T_2267; // @[Mux.scala 19:72:@2933.4]
  assign _T_2357 = _T_2356 | _T_2269; // @[Mux.scala 19:72:@2934.4]
  assign _T_2358 = _T_2357 | _T_2271; // @[Mux.scala 19:72:@2935.4]
  assign _T_2359 = _T_2358 | _T_2273; // @[Mux.scala 19:72:@2936.4]
  assign _T_2360 = _T_2359 | _T_2275; // @[Mux.scala 19:72:@2937.4]
  assign _T_2361 = _T_2360 | _T_2277; // @[Mux.scala 19:72:@2938.4]
  assign _T_2362 = _T_2361 | _T_2279; // @[Mux.scala 19:72:@2939.4]
  assign _T_2363 = _T_2362 | _T_2281; // @[Mux.scala 19:72:@2940.4]
  assign _T_2364 = _T_2363 | _T_2283; // @[Mux.scala 19:72:@2941.4]
  assign _T_2365 = _T_2364 | _T_2285; // @[Mux.scala 19:72:@2942.4]
  assign _T_2366 = _T_2365 | _T_2287; // @[Mux.scala 19:72:@2943.4]
  assign _T_2367 = _T_2366 | _T_2289; // @[Mux.scala 19:72:@2944.4]
  assign _T_2368 = _T_2367 | _T_2291; // @[Mux.scala 19:72:@2945.4]
  assign _T_2369 = _T_2368 | _T_2293; // @[Mux.scala 19:72:@2946.4]
  assign _T_2370 = _T_2369 | _T_2295; // @[Mux.scala 19:72:@2947.4]
  assign _T_2371 = _T_2370 | _T_2297; // @[Mux.scala 19:72:@2948.4]
  assign _T_2372 = _T_2371 | _T_2299; // @[Mux.scala 19:72:@2949.4]
  assign _T_2373 = _T_2372 | _T_2301; // @[Mux.scala 19:72:@2950.4]
  assign _T_2374 = _T_2373 | _T_2303; // @[Mux.scala 19:72:@2951.4]
  assign _T_2375 = _T_2374 | _T_2305; // @[Mux.scala 19:72:@2952.4]
  assign _T_2376 = _T_2375 | _T_2307; // @[Mux.scala 19:72:@2953.4]
  assign _T_2377 = _T_2376 | _T_2309; // @[Mux.scala 19:72:@2954.4]
  assign _T_2378 = _T_2377 | _T_2311; // @[Mux.scala 19:72:@2955.4]
  assign _T_2379 = _T_2378 | _T_2313; // @[Mux.scala 19:72:@2956.4]
  assign _T_2380 = _T_2379 | _T_2315; // @[Mux.scala 19:72:@2957.4]
  assign _T_2381 = _T_2380 | _T_2317; // @[Mux.scala 19:72:@2958.4]
  assign predict_1_btype = _T_2381 | _T_2319; // @[Mux.scala 19:72:@2959.4]
  assign _T_2451 = _T_1869 ? btb_hcount_0 : 2'h0; // @[Mux.scala 19:72:@3027.4]
  assign _T_2453 = _T_1870 ? btb_hcount_1 : 2'h0; // @[Mux.scala 19:72:@3028.4]
  assign _T_2455 = _T_1871 ? btb_hcount_2 : 2'h0; // @[Mux.scala 19:72:@3029.4]
  assign _T_2457 = _T_1872 ? btb_hcount_3 : 2'h0; // @[Mux.scala 19:72:@3030.4]
  assign _T_2459 = _T_1873 ? btb_hcount_4 : 2'h0; // @[Mux.scala 19:72:@3031.4]
  assign _T_2461 = _T_1874 ? btb_hcount_5 : 2'h0; // @[Mux.scala 19:72:@3032.4]
  assign _T_2463 = _T_1875 ? btb_hcount_6 : 2'h0; // @[Mux.scala 19:72:@3033.4]
  assign _T_2465 = _T_1876 ? btb_hcount_7 : 2'h0; // @[Mux.scala 19:72:@3034.4]
  assign _T_2467 = _T_1877 ? btb_hcount_8 : 2'h0; // @[Mux.scala 19:72:@3035.4]
  assign _T_2469 = _T_1878 ? btb_hcount_9 : 2'h0; // @[Mux.scala 19:72:@3036.4]
  assign _T_2471 = _T_1879 ? btb_hcount_10 : 2'h0; // @[Mux.scala 19:72:@3037.4]
  assign _T_2473 = _T_1880 ? btb_hcount_11 : 2'h0; // @[Mux.scala 19:72:@3038.4]
  assign _T_2475 = _T_1881 ? btb_hcount_12 : 2'h0; // @[Mux.scala 19:72:@3039.4]
  assign _T_2477 = _T_1882 ? btb_hcount_13 : 2'h0; // @[Mux.scala 19:72:@3040.4]
  assign _T_2479 = _T_1883 ? btb_hcount_14 : 2'h0; // @[Mux.scala 19:72:@3041.4]
  assign _T_2481 = _T_1884 ? btb_hcount_15 : 2'h0; // @[Mux.scala 19:72:@3042.4]
  assign _T_2483 = _T_1885 ? btb_hcount_16 : 2'h0; // @[Mux.scala 19:72:@3043.4]
  assign _T_2485 = _T_1886 ? btb_hcount_17 : 2'h0; // @[Mux.scala 19:72:@3044.4]
  assign _T_2487 = _T_1887 ? btb_hcount_18 : 2'h0; // @[Mux.scala 19:72:@3045.4]
  assign _T_2489 = _T_1888 ? btb_hcount_19 : 2'h0; // @[Mux.scala 19:72:@3046.4]
  assign _T_2491 = _T_1889 ? btb_hcount_20 : 2'h0; // @[Mux.scala 19:72:@3047.4]
  assign _T_2493 = _T_1890 ? btb_hcount_21 : 2'h0; // @[Mux.scala 19:72:@3048.4]
  assign _T_2495 = _T_1891 ? btb_hcount_22 : 2'h0; // @[Mux.scala 19:72:@3049.4]
  assign _T_2497 = _T_1892 ? btb_hcount_23 : 2'h0; // @[Mux.scala 19:72:@3050.4]
  assign _T_2499 = _T_1893 ? btb_hcount_24 : 2'h0; // @[Mux.scala 19:72:@3051.4]
  assign _T_2501 = _T_1894 ? btb_hcount_25 : 2'h0; // @[Mux.scala 19:72:@3052.4]
  assign _T_2503 = _T_1895 ? btb_hcount_26 : 2'h0; // @[Mux.scala 19:72:@3053.4]
  assign _T_2505 = _T_1896 ? btb_hcount_27 : 2'h0; // @[Mux.scala 19:72:@3054.4]
  assign _T_2507 = _T_1897 ? btb_hcount_28 : 2'h0; // @[Mux.scala 19:72:@3055.4]
  assign _T_2509 = _T_1898 ? btb_hcount_29 : 2'h0; // @[Mux.scala 19:72:@3056.4]
  assign _T_2511 = _T_1899 ? btb_hcount_30 : 2'h0; // @[Mux.scala 19:72:@3057.4]
  assign _T_2513 = _T_1900 ? btb_hcount_31 : 2'h0; // @[Mux.scala 19:72:@3058.4]
  assign _T_2515 = _T_1901 ? btb_hcount_32 : 2'h0; // @[Mux.scala 19:72:@3059.4]
  assign _T_2517 = _T_1902 ? btb_hcount_33 : 2'h0; // @[Mux.scala 19:72:@3060.4]
  assign _T_2519 = _T_1903 ? btb_hcount_34 : 2'h0; // @[Mux.scala 19:72:@3061.4]
  assign _T_2521 = _T_1904 ? btb_hcount_35 : 2'h0; // @[Mux.scala 19:72:@3062.4]
  assign _T_2523 = _T_1905 ? btb_hcount_36 : 2'h0; // @[Mux.scala 19:72:@3063.4]
  assign _T_2525 = _T_1906 ? btb_hcount_37 : 2'h0; // @[Mux.scala 19:72:@3064.4]
  assign _T_2527 = _T_1907 ? btb_hcount_38 : 2'h0; // @[Mux.scala 19:72:@3065.4]
  assign _T_2529 = _T_1908 ? btb_hcount_39 : 2'h0; // @[Mux.scala 19:72:@3066.4]
  assign _T_2531 = _T_1909 ? btb_hcount_40 : 2'h0; // @[Mux.scala 19:72:@3067.4]
  assign _T_2533 = _T_1910 ? btb_hcount_41 : 2'h0; // @[Mux.scala 19:72:@3068.4]
  assign _T_2535 = _T_1911 ? btb_hcount_42 : 2'h0; // @[Mux.scala 19:72:@3069.4]
  assign _T_2537 = _T_1912 ? btb_hcount_43 : 2'h0; // @[Mux.scala 19:72:@3070.4]
  assign _T_2539 = _T_1913 ? btb_hcount_44 : 2'h0; // @[Mux.scala 19:72:@3071.4]
  assign _T_2541 = _T_1914 ? btb_hcount_45 : 2'h0; // @[Mux.scala 19:72:@3072.4]
  assign _T_2543 = _T_1915 ? btb_hcount_46 : 2'h0; // @[Mux.scala 19:72:@3073.4]
  assign _T_2545 = _T_1916 ? btb_hcount_47 : 2'h0; // @[Mux.scala 19:72:@3074.4]
  assign _T_2547 = _T_1917 ? btb_hcount_48 : 2'h0; // @[Mux.scala 19:72:@3075.4]
  assign _T_2549 = _T_1918 ? btb_hcount_49 : 2'h0; // @[Mux.scala 19:72:@3076.4]
  assign _T_2551 = _T_1919 ? btb_hcount_50 : 2'h0; // @[Mux.scala 19:72:@3077.4]
  assign _T_2553 = _T_1920 ? btb_hcount_51 : 2'h0; // @[Mux.scala 19:72:@3078.4]
  assign _T_2555 = _T_1921 ? btb_hcount_52 : 2'h0; // @[Mux.scala 19:72:@3079.4]
  assign _T_2557 = _T_1922 ? btb_hcount_53 : 2'h0; // @[Mux.scala 19:72:@3080.4]
  assign _T_2559 = _T_1923 ? btb_hcount_54 : 2'h0; // @[Mux.scala 19:72:@3081.4]
  assign _T_2561 = _T_1924 ? btb_hcount_55 : 2'h0; // @[Mux.scala 19:72:@3082.4]
  assign _T_2563 = _T_1925 ? btb_hcount_56 : 2'h0; // @[Mux.scala 19:72:@3083.4]
  assign _T_2565 = _T_1926 ? btb_hcount_57 : 2'h0; // @[Mux.scala 19:72:@3084.4]
  assign _T_2567 = _T_1927 ? btb_hcount_58 : 2'h0; // @[Mux.scala 19:72:@3085.4]
  assign _T_2569 = _T_1928 ? btb_hcount_59 : 2'h0; // @[Mux.scala 19:72:@3086.4]
  assign _T_2571 = _T_1929 ? btb_hcount_60 : 2'h0; // @[Mux.scala 19:72:@3087.4]
  assign _T_2573 = _T_1930 ? btb_hcount_61 : 2'h0; // @[Mux.scala 19:72:@3088.4]
  assign _T_2575 = _T_1931 ? btb_hcount_62 : 2'h0; // @[Mux.scala 19:72:@3089.4]
  assign _T_2577 = _T_1932 ? btb_hcount_63 : 2'h0; // @[Mux.scala 19:72:@3090.4]
  assign _T_2578 = _T_2451 | _T_2453; // @[Mux.scala 19:72:@3091.4]
  assign _T_2579 = _T_2578 | _T_2455; // @[Mux.scala 19:72:@3092.4]
  assign _T_2580 = _T_2579 | _T_2457; // @[Mux.scala 19:72:@3093.4]
  assign _T_2581 = _T_2580 | _T_2459; // @[Mux.scala 19:72:@3094.4]
  assign _T_2582 = _T_2581 | _T_2461; // @[Mux.scala 19:72:@3095.4]
  assign _T_2583 = _T_2582 | _T_2463; // @[Mux.scala 19:72:@3096.4]
  assign _T_2584 = _T_2583 | _T_2465; // @[Mux.scala 19:72:@3097.4]
  assign _T_2585 = _T_2584 | _T_2467; // @[Mux.scala 19:72:@3098.4]
  assign _T_2586 = _T_2585 | _T_2469; // @[Mux.scala 19:72:@3099.4]
  assign _T_2587 = _T_2586 | _T_2471; // @[Mux.scala 19:72:@3100.4]
  assign _T_2588 = _T_2587 | _T_2473; // @[Mux.scala 19:72:@3101.4]
  assign _T_2589 = _T_2588 | _T_2475; // @[Mux.scala 19:72:@3102.4]
  assign _T_2590 = _T_2589 | _T_2477; // @[Mux.scala 19:72:@3103.4]
  assign _T_2591 = _T_2590 | _T_2479; // @[Mux.scala 19:72:@3104.4]
  assign _T_2592 = _T_2591 | _T_2481; // @[Mux.scala 19:72:@3105.4]
  assign _T_2593 = _T_2592 | _T_2483; // @[Mux.scala 19:72:@3106.4]
  assign _T_2594 = _T_2593 | _T_2485; // @[Mux.scala 19:72:@3107.4]
  assign _T_2595 = _T_2594 | _T_2487; // @[Mux.scala 19:72:@3108.4]
  assign _T_2596 = _T_2595 | _T_2489; // @[Mux.scala 19:72:@3109.4]
  assign _T_2597 = _T_2596 | _T_2491; // @[Mux.scala 19:72:@3110.4]
  assign _T_2598 = _T_2597 | _T_2493; // @[Mux.scala 19:72:@3111.4]
  assign _T_2599 = _T_2598 | _T_2495; // @[Mux.scala 19:72:@3112.4]
  assign _T_2600 = _T_2599 | _T_2497; // @[Mux.scala 19:72:@3113.4]
  assign _T_2601 = _T_2600 | _T_2499; // @[Mux.scala 19:72:@3114.4]
  assign _T_2602 = _T_2601 | _T_2501; // @[Mux.scala 19:72:@3115.4]
  assign _T_2603 = _T_2602 | _T_2503; // @[Mux.scala 19:72:@3116.4]
  assign _T_2604 = _T_2603 | _T_2505; // @[Mux.scala 19:72:@3117.4]
  assign _T_2605 = _T_2604 | _T_2507; // @[Mux.scala 19:72:@3118.4]
  assign _T_2606 = _T_2605 | _T_2509; // @[Mux.scala 19:72:@3119.4]
  assign _T_2607 = _T_2606 | _T_2511; // @[Mux.scala 19:72:@3120.4]
  assign _T_2608 = _T_2607 | _T_2513; // @[Mux.scala 19:72:@3121.4]
  assign _T_2609 = _T_2608 | _T_2515; // @[Mux.scala 19:72:@3122.4]
  assign _T_2610 = _T_2609 | _T_2517; // @[Mux.scala 19:72:@3123.4]
  assign _T_2611 = _T_2610 | _T_2519; // @[Mux.scala 19:72:@3124.4]
  assign _T_2612 = _T_2611 | _T_2521; // @[Mux.scala 19:72:@3125.4]
  assign _T_2613 = _T_2612 | _T_2523; // @[Mux.scala 19:72:@3126.4]
  assign _T_2614 = _T_2613 | _T_2525; // @[Mux.scala 19:72:@3127.4]
  assign _T_2615 = _T_2614 | _T_2527; // @[Mux.scala 19:72:@3128.4]
  assign _T_2616 = _T_2615 | _T_2529; // @[Mux.scala 19:72:@3129.4]
  assign _T_2617 = _T_2616 | _T_2531; // @[Mux.scala 19:72:@3130.4]
  assign _T_2618 = _T_2617 | _T_2533; // @[Mux.scala 19:72:@3131.4]
  assign _T_2619 = _T_2618 | _T_2535; // @[Mux.scala 19:72:@3132.4]
  assign _T_2620 = _T_2619 | _T_2537; // @[Mux.scala 19:72:@3133.4]
  assign _T_2621 = _T_2620 | _T_2539; // @[Mux.scala 19:72:@3134.4]
  assign _T_2622 = _T_2621 | _T_2541; // @[Mux.scala 19:72:@3135.4]
  assign _T_2623 = _T_2622 | _T_2543; // @[Mux.scala 19:72:@3136.4]
  assign _T_2624 = _T_2623 | _T_2545; // @[Mux.scala 19:72:@3137.4]
  assign _T_2625 = _T_2624 | _T_2547; // @[Mux.scala 19:72:@3138.4]
  assign _T_2626 = _T_2625 | _T_2549; // @[Mux.scala 19:72:@3139.4]
  assign _T_2627 = _T_2626 | _T_2551; // @[Mux.scala 19:72:@3140.4]
  assign _T_2628 = _T_2627 | _T_2553; // @[Mux.scala 19:72:@3141.4]
  assign _T_2629 = _T_2628 | _T_2555; // @[Mux.scala 19:72:@3142.4]
  assign _T_2630 = _T_2629 | _T_2557; // @[Mux.scala 19:72:@3143.4]
  assign _T_2631 = _T_2630 | _T_2559; // @[Mux.scala 19:72:@3144.4]
  assign _T_2632 = _T_2631 | _T_2561; // @[Mux.scala 19:72:@3145.4]
  assign _T_2633 = _T_2632 | _T_2563; // @[Mux.scala 19:72:@3146.4]
  assign _T_2634 = _T_2633 | _T_2565; // @[Mux.scala 19:72:@3147.4]
  assign _T_2635 = _T_2634 | _T_2567; // @[Mux.scala 19:72:@3148.4]
  assign _T_2636 = _T_2635 | _T_2569; // @[Mux.scala 19:72:@3149.4]
  assign _T_2637 = _T_2636 | _T_2571; // @[Mux.scala 19:72:@3150.4]
  assign _T_2638 = _T_2637 | _T_2573; // @[Mux.scala 19:72:@3151.4]
  assign _T_2639 = _T_2638 | _T_2575; // @[Mux.scala 19:72:@3152.4]
  assign predict_1_hcount = _T_2639 | _T_2577; // @[Mux.scala 19:72:@3153.4]
  assign _T_2644 = predict_1_btype == 2'h1; // @[BTB.scala 80:44:@3157.4]
  assign _T_2646 = predict_1_btype == 2'h2; // @[BTB.scala 69:34:@3158.4]
  assign _T_2647 = predict_1_hcount[1]; // @[BTB.scala 69:65:@3159.4]
  assign _T_2649 = _T_2647 == 1'h0; // @[BTB.scala 69:58:@3160.4]
  assign _T_2650 = _T_2646 & _T_2649; // @[BTB.scala 69:55:@3161.4]
  assign _T_2652 = _T_2650 == 1'h0; // @[BTB.scala 69:26:@3162.4]
  assign _T_2654 = predict_1_lookup != 64'h0; // @[BTB.scala 69:80:@3163.4]
  assign _T_2655 = _T_2652 & _T_2654; // @[BTB.scala 69:70:@3164.4]
  assign _T_2659 = if_pc_1 + 32'h4; // @[BTB.scala 84:35:@3169.4]
  assign predict_1_cont_tgt = if_pc_1 + 32'h4; // @[BTB.scala 84:35:@3170.4]
  assign _T_2656 = _T_2655 ? predict_1_jump_tgt : predict_1_cont_tgt; // @[BTB.scala 70:27:@3165.4]
  assign _T_2672 = io_if_pc[2]; // @[BTB.scala 85:47:@3179.4]
  assign _T_2675 = _T_2672 == 1'h0; // @[BTB.scala 85:38:@3181.4]
  assign _T_2683 = fb_reg_lfsr[0]; // @[BTB.scala 99:36:@3197.4]
  assign _T_2684 = fb_reg_lfsr[1]; // @[BTB.scala 99:46:@3198.4]
  assign _T_2685 = _T_2683 ^ _T_2684; // @[BTB.scala 99:40:@3199.4]
  assign _T_2686 = fb_reg_lfsr[5:1]; // @[BTB.scala 99:55:@3200.4]
  assign _T_2687 = {_T_2685,_T_2686}; // @[Cat.scala 30:58:@3201.4]
  assign _T_2689 = btb_pc_0 == fb_reg_pc; // @[BTB.scala 123:42:@3204.4]
  assign _T_2690 = btb_pc_1 == fb_reg_pc; // @[BTB.scala 123:42:@3205.4]
  assign _T_2691 = btb_pc_2 == fb_reg_pc; // @[BTB.scala 123:42:@3206.4]
  assign _T_2692 = btb_pc_3 == fb_reg_pc; // @[BTB.scala 123:42:@3207.4]
  assign _T_2693 = btb_pc_4 == fb_reg_pc; // @[BTB.scala 123:42:@3208.4]
  assign _T_2694 = btb_pc_5 == fb_reg_pc; // @[BTB.scala 123:42:@3209.4]
  assign _T_2695 = btb_pc_6 == fb_reg_pc; // @[BTB.scala 123:42:@3210.4]
  assign _T_2696 = btb_pc_7 == fb_reg_pc; // @[BTB.scala 123:42:@3211.4]
  assign _T_2697 = btb_pc_8 == fb_reg_pc; // @[BTB.scala 123:42:@3212.4]
  assign _T_2698 = btb_pc_9 == fb_reg_pc; // @[BTB.scala 123:42:@3213.4]
  assign _T_2699 = btb_pc_10 == fb_reg_pc; // @[BTB.scala 123:42:@3214.4]
  assign _T_2700 = btb_pc_11 == fb_reg_pc; // @[BTB.scala 123:42:@3215.4]
  assign _T_2701 = btb_pc_12 == fb_reg_pc; // @[BTB.scala 123:42:@3216.4]
  assign _T_2702 = btb_pc_13 == fb_reg_pc; // @[BTB.scala 123:42:@3217.4]
  assign _T_2703 = btb_pc_14 == fb_reg_pc; // @[BTB.scala 123:42:@3218.4]
  assign _T_2704 = btb_pc_15 == fb_reg_pc; // @[BTB.scala 123:42:@3219.4]
  assign _T_2705 = btb_pc_16 == fb_reg_pc; // @[BTB.scala 123:42:@3220.4]
  assign _T_2706 = btb_pc_17 == fb_reg_pc; // @[BTB.scala 123:42:@3221.4]
  assign _T_2707 = btb_pc_18 == fb_reg_pc; // @[BTB.scala 123:42:@3222.4]
  assign _T_2708 = btb_pc_19 == fb_reg_pc; // @[BTB.scala 123:42:@3223.4]
  assign _T_2709 = btb_pc_20 == fb_reg_pc; // @[BTB.scala 123:42:@3224.4]
  assign _T_2710 = btb_pc_21 == fb_reg_pc; // @[BTB.scala 123:42:@3225.4]
  assign _T_2711 = btb_pc_22 == fb_reg_pc; // @[BTB.scala 123:42:@3226.4]
  assign _T_2712 = btb_pc_23 == fb_reg_pc; // @[BTB.scala 123:42:@3227.4]
  assign _T_2713 = btb_pc_24 == fb_reg_pc; // @[BTB.scala 123:42:@3228.4]
  assign _T_2714 = btb_pc_25 == fb_reg_pc; // @[BTB.scala 123:42:@3229.4]
  assign _T_2715 = btb_pc_26 == fb_reg_pc; // @[BTB.scala 123:42:@3230.4]
  assign _T_2716 = btb_pc_27 == fb_reg_pc; // @[BTB.scala 123:42:@3231.4]
  assign _T_2717 = btb_pc_28 == fb_reg_pc; // @[BTB.scala 123:42:@3232.4]
  assign _T_2718 = btb_pc_29 == fb_reg_pc; // @[BTB.scala 123:42:@3233.4]
  assign _T_2719 = btb_pc_30 == fb_reg_pc; // @[BTB.scala 123:42:@3234.4]
  assign _T_2720 = btb_pc_31 == fb_reg_pc; // @[BTB.scala 123:42:@3235.4]
  assign _T_2721 = btb_pc_32 == fb_reg_pc; // @[BTB.scala 123:42:@3236.4]
  assign _T_2722 = btb_pc_33 == fb_reg_pc; // @[BTB.scala 123:42:@3237.4]
  assign _T_2723 = btb_pc_34 == fb_reg_pc; // @[BTB.scala 123:42:@3238.4]
  assign _T_2724 = btb_pc_35 == fb_reg_pc; // @[BTB.scala 123:42:@3239.4]
  assign _T_2725 = btb_pc_36 == fb_reg_pc; // @[BTB.scala 123:42:@3240.4]
  assign _T_2726 = btb_pc_37 == fb_reg_pc; // @[BTB.scala 123:42:@3241.4]
  assign _T_2727 = btb_pc_38 == fb_reg_pc; // @[BTB.scala 123:42:@3242.4]
  assign _T_2728 = btb_pc_39 == fb_reg_pc; // @[BTB.scala 123:42:@3243.4]
  assign _T_2729 = btb_pc_40 == fb_reg_pc; // @[BTB.scala 123:42:@3244.4]
  assign _T_2730 = btb_pc_41 == fb_reg_pc; // @[BTB.scala 123:42:@3245.4]
  assign _T_2731 = btb_pc_42 == fb_reg_pc; // @[BTB.scala 123:42:@3246.4]
  assign _T_2732 = btb_pc_43 == fb_reg_pc; // @[BTB.scala 123:42:@3247.4]
  assign _T_2733 = btb_pc_44 == fb_reg_pc; // @[BTB.scala 123:42:@3248.4]
  assign _T_2734 = btb_pc_45 == fb_reg_pc; // @[BTB.scala 123:42:@3249.4]
  assign _T_2735 = btb_pc_46 == fb_reg_pc; // @[BTB.scala 123:42:@3250.4]
  assign _T_2736 = btb_pc_47 == fb_reg_pc; // @[BTB.scala 123:42:@3251.4]
  assign _T_2737 = btb_pc_48 == fb_reg_pc; // @[BTB.scala 123:42:@3252.4]
  assign _T_2738 = btb_pc_49 == fb_reg_pc; // @[BTB.scala 123:42:@3253.4]
  assign _T_2739 = btb_pc_50 == fb_reg_pc; // @[BTB.scala 123:42:@3254.4]
  assign _T_2740 = btb_pc_51 == fb_reg_pc; // @[BTB.scala 123:42:@3255.4]
  assign _T_2741 = btb_pc_52 == fb_reg_pc; // @[BTB.scala 123:42:@3256.4]
  assign _T_2742 = btb_pc_53 == fb_reg_pc; // @[BTB.scala 123:42:@3257.4]
  assign _T_2743 = btb_pc_54 == fb_reg_pc; // @[BTB.scala 123:42:@3258.4]
  assign _T_2744 = btb_pc_55 == fb_reg_pc; // @[BTB.scala 123:42:@3259.4]
  assign _T_2745 = btb_pc_56 == fb_reg_pc; // @[BTB.scala 123:42:@3260.4]
  assign _T_2746 = btb_pc_57 == fb_reg_pc; // @[BTB.scala 123:42:@3261.4]
  assign _T_2747 = btb_pc_58 == fb_reg_pc; // @[BTB.scala 123:42:@3262.4]
  assign _T_2748 = btb_pc_59 == fb_reg_pc; // @[BTB.scala 123:42:@3263.4]
  assign _T_2749 = btb_pc_60 == fb_reg_pc; // @[BTB.scala 123:42:@3264.4]
  assign _T_2750 = btb_pc_61 == fb_reg_pc; // @[BTB.scala 123:42:@3265.4]
  assign _T_2751 = btb_pc_62 == fb_reg_pc; // @[BTB.scala 123:42:@3266.4]
  assign _T_2752 = btb_pc_63 == fb_reg_pc; // @[BTB.scala 123:42:@3267.4]
  assign _T_2829 = {_T_2696,_T_2695,_T_2694,_T_2693,_T_2692,_T_2691,_T_2690,_T_2689}; // @[BTB.scala 123:58:@3339.4]
  assign _T_2837 = {_T_2704,_T_2703,_T_2702,_T_2701,_T_2700,_T_2699,_T_2698,_T_2697,_T_2829}; // @[BTB.scala 123:58:@3347.4]
  assign _T_2844 = {_T_2712,_T_2711,_T_2710,_T_2709,_T_2708,_T_2707,_T_2706,_T_2705}; // @[BTB.scala 123:58:@3354.4]
  assign _T_2853 = {_T_2720,_T_2719,_T_2718,_T_2717,_T_2716,_T_2715,_T_2714,_T_2713,_T_2844,_T_2837}; // @[BTB.scala 123:58:@3363.4]
  assign _T_2860 = {_T_2728,_T_2727,_T_2726,_T_2725,_T_2724,_T_2723,_T_2722,_T_2721}; // @[BTB.scala 123:58:@3370.4]
  assign _T_2868 = {_T_2736,_T_2735,_T_2734,_T_2733,_T_2732,_T_2731,_T_2730,_T_2729,_T_2860}; // @[BTB.scala 123:58:@3378.4]
  assign _T_2875 = {_T_2744,_T_2743,_T_2742,_T_2741,_T_2740,_T_2739,_T_2738,_T_2737}; // @[BTB.scala 123:58:@3385.4]
  assign _T_2884 = {_T_2752,_T_2751,_T_2750,_T_2749,_T_2748,_T_2747,_T_2746,_T_2745,_T_2875,_T_2868}; // @[BTB.scala 123:58:@3394.4]
  assign _T_2885 = {_T_2884,_T_2853}; // @[BTB.scala 123:58:@3395.4]
  assign fb_wire_lookup = _T_2885 & _T_614; // @[BTB.scala 123:65:@3588.4]
  assign _T_3148 = fb_wire_lookup[0]; // @[Mux.scala 21:36:@3590.4]
  assign _T_3149 = fb_wire_lookup[1]; // @[Mux.scala 21:36:@3591.4]
  assign _T_3150 = fb_wire_lookup[2]; // @[Mux.scala 21:36:@3592.4]
  assign _T_3151 = fb_wire_lookup[3]; // @[Mux.scala 21:36:@3593.4]
  assign _T_3152 = fb_wire_lookup[4]; // @[Mux.scala 21:36:@3594.4]
  assign _T_3153 = fb_wire_lookup[5]; // @[Mux.scala 21:36:@3595.4]
  assign _T_3154 = fb_wire_lookup[6]; // @[Mux.scala 21:36:@3596.4]
  assign _T_3155 = fb_wire_lookup[7]; // @[Mux.scala 21:36:@3597.4]
  assign _T_3156 = fb_wire_lookup[8]; // @[Mux.scala 21:36:@3598.4]
  assign _T_3157 = fb_wire_lookup[9]; // @[Mux.scala 21:36:@3599.4]
  assign _T_3158 = fb_wire_lookup[10]; // @[Mux.scala 21:36:@3600.4]
  assign _T_3159 = fb_wire_lookup[11]; // @[Mux.scala 21:36:@3601.4]
  assign _T_3160 = fb_wire_lookup[12]; // @[Mux.scala 21:36:@3602.4]
  assign _T_3161 = fb_wire_lookup[13]; // @[Mux.scala 21:36:@3603.4]
  assign _T_3162 = fb_wire_lookup[14]; // @[Mux.scala 21:36:@3604.4]
  assign _T_3163 = fb_wire_lookup[15]; // @[Mux.scala 21:36:@3605.4]
  assign _T_3164 = fb_wire_lookup[16]; // @[Mux.scala 21:36:@3606.4]
  assign _T_3165 = fb_wire_lookup[17]; // @[Mux.scala 21:36:@3607.4]
  assign _T_3166 = fb_wire_lookup[18]; // @[Mux.scala 21:36:@3608.4]
  assign _T_3167 = fb_wire_lookup[19]; // @[Mux.scala 21:36:@3609.4]
  assign _T_3168 = fb_wire_lookup[20]; // @[Mux.scala 21:36:@3610.4]
  assign _T_3169 = fb_wire_lookup[21]; // @[Mux.scala 21:36:@3611.4]
  assign _T_3170 = fb_wire_lookup[22]; // @[Mux.scala 21:36:@3612.4]
  assign _T_3171 = fb_wire_lookup[23]; // @[Mux.scala 21:36:@3613.4]
  assign _T_3172 = fb_wire_lookup[24]; // @[Mux.scala 21:36:@3614.4]
  assign _T_3173 = fb_wire_lookup[25]; // @[Mux.scala 21:36:@3615.4]
  assign _T_3174 = fb_wire_lookup[26]; // @[Mux.scala 21:36:@3616.4]
  assign _T_3175 = fb_wire_lookup[27]; // @[Mux.scala 21:36:@3617.4]
  assign _T_3176 = fb_wire_lookup[28]; // @[Mux.scala 21:36:@3618.4]
  assign _T_3177 = fb_wire_lookup[29]; // @[Mux.scala 21:36:@3619.4]
  assign _T_3178 = fb_wire_lookup[30]; // @[Mux.scala 21:36:@3620.4]
  assign _T_3179 = fb_wire_lookup[31]; // @[Mux.scala 21:36:@3621.4]
  assign _T_3180 = fb_wire_lookup[32]; // @[Mux.scala 21:36:@3622.4]
  assign _T_3181 = fb_wire_lookup[33]; // @[Mux.scala 21:36:@3623.4]
  assign _T_3182 = fb_wire_lookup[34]; // @[Mux.scala 21:36:@3624.4]
  assign _T_3183 = fb_wire_lookup[35]; // @[Mux.scala 21:36:@3625.4]
  assign _T_3184 = fb_wire_lookup[36]; // @[Mux.scala 21:36:@3626.4]
  assign _T_3185 = fb_wire_lookup[37]; // @[Mux.scala 21:36:@3627.4]
  assign _T_3186 = fb_wire_lookup[38]; // @[Mux.scala 21:36:@3628.4]
  assign _T_3187 = fb_wire_lookup[39]; // @[Mux.scala 21:36:@3629.4]
  assign _T_3188 = fb_wire_lookup[40]; // @[Mux.scala 21:36:@3630.4]
  assign _T_3189 = fb_wire_lookup[41]; // @[Mux.scala 21:36:@3631.4]
  assign _T_3190 = fb_wire_lookup[42]; // @[Mux.scala 21:36:@3632.4]
  assign _T_3191 = fb_wire_lookup[43]; // @[Mux.scala 21:36:@3633.4]
  assign _T_3192 = fb_wire_lookup[44]; // @[Mux.scala 21:36:@3634.4]
  assign _T_3193 = fb_wire_lookup[45]; // @[Mux.scala 21:36:@3635.4]
  assign _T_3194 = fb_wire_lookup[46]; // @[Mux.scala 21:36:@3636.4]
  assign _T_3195 = fb_wire_lookup[47]; // @[Mux.scala 21:36:@3637.4]
  assign _T_3196 = fb_wire_lookup[48]; // @[Mux.scala 21:36:@3638.4]
  assign _T_3197 = fb_wire_lookup[49]; // @[Mux.scala 21:36:@3639.4]
  assign _T_3198 = fb_wire_lookup[50]; // @[Mux.scala 21:36:@3640.4]
  assign _T_3199 = fb_wire_lookup[51]; // @[Mux.scala 21:36:@3641.4]
  assign _T_3200 = fb_wire_lookup[52]; // @[Mux.scala 21:36:@3642.4]
  assign _T_3201 = fb_wire_lookup[53]; // @[Mux.scala 21:36:@3643.4]
  assign _T_3202 = fb_wire_lookup[54]; // @[Mux.scala 21:36:@3644.4]
  assign _T_3203 = fb_wire_lookup[55]; // @[Mux.scala 21:36:@3645.4]
  assign _T_3204 = fb_wire_lookup[56]; // @[Mux.scala 21:36:@3646.4]
  assign _T_3205 = fb_wire_lookup[57]; // @[Mux.scala 21:36:@3647.4]
  assign _T_3206 = fb_wire_lookup[58]; // @[Mux.scala 21:36:@3648.4]
  assign _T_3207 = fb_wire_lookup[59]; // @[Mux.scala 21:36:@3649.4]
  assign _T_3208 = fb_wire_lookup[60]; // @[Mux.scala 21:36:@3650.4]
  assign _T_3209 = fb_wire_lookup[61]; // @[Mux.scala 21:36:@3651.4]
  assign _T_3210 = fb_wire_lookup[62]; // @[Mux.scala 21:36:@3652.4]
  assign _T_3211 = fb_wire_lookup[63]; // @[Mux.scala 21:36:@3653.4]
  assign _T_3214 = _T_3148 ? btb_hcount_0 : 2'h0; // @[Mux.scala 19:72:@3654.4]
  assign _T_3216 = _T_3149 ? btb_hcount_1 : 2'h0; // @[Mux.scala 19:72:@3655.4]
  assign _T_3218 = _T_3150 ? btb_hcount_2 : 2'h0; // @[Mux.scala 19:72:@3656.4]
  assign _T_3220 = _T_3151 ? btb_hcount_3 : 2'h0; // @[Mux.scala 19:72:@3657.4]
  assign _T_3222 = _T_3152 ? btb_hcount_4 : 2'h0; // @[Mux.scala 19:72:@3658.4]
  assign _T_3224 = _T_3153 ? btb_hcount_5 : 2'h0; // @[Mux.scala 19:72:@3659.4]
  assign _T_3226 = _T_3154 ? btb_hcount_6 : 2'h0; // @[Mux.scala 19:72:@3660.4]
  assign _T_3228 = _T_3155 ? btb_hcount_7 : 2'h0; // @[Mux.scala 19:72:@3661.4]
  assign _T_3230 = _T_3156 ? btb_hcount_8 : 2'h0; // @[Mux.scala 19:72:@3662.4]
  assign _T_3232 = _T_3157 ? btb_hcount_9 : 2'h0; // @[Mux.scala 19:72:@3663.4]
  assign _T_3234 = _T_3158 ? btb_hcount_10 : 2'h0; // @[Mux.scala 19:72:@3664.4]
  assign _T_3236 = _T_3159 ? btb_hcount_11 : 2'h0; // @[Mux.scala 19:72:@3665.4]
  assign _T_3238 = _T_3160 ? btb_hcount_12 : 2'h0; // @[Mux.scala 19:72:@3666.4]
  assign _T_3240 = _T_3161 ? btb_hcount_13 : 2'h0; // @[Mux.scala 19:72:@3667.4]
  assign _T_3242 = _T_3162 ? btb_hcount_14 : 2'h0; // @[Mux.scala 19:72:@3668.4]
  assign _T_3244 = _T_3163 ? btb_hcount_15 : 2'h0; // @[Mux.scala 19:72:@3669.4]
  assign _T_3246 = _T_3164 ? btb_hcount_16 : 2'h0; // @[Mux.scala 19:72:@3670.4]
  assign _T_3248 = _T_3165 ? btb_hcount_17 : 2'h0; // @[Mux.scala 19:72:@3671.4]
  assign _T_3250 = _T_3166 ? btb_hcount_18 : 2'h0; // @[Mux.scala 19:72:@3672.4]
  assign _T_3252 = _T_3167 ? btb_hcount_19 : 2'h0; // @[Mux.scala 19:72:@3673.4]
  assign _T_3254 = _T_3168 ? btb_hcount_20 : 2'h0; // @[Mux.scala 19:72:@3674.4]
  assign _T_3256 = _T_3169 ? btb_hcount_21 : 2'h0; // @[Mux.scala 19:72:@3675.4]
  assign _T_3258 = _T_3170 ? btb_hcount_22 : 2'h0; // @[Mux.scala 19:72:@3676.4]
  assign _T_3260 = _T_3171 ? btb_hcount_23 : 2'h0; // @[Mux.scala 19:72:@3677.4]
  assign _T_3262 = _T_3172 ? btb_hcount_24 : 2'h0; // @[Mux.scala 19:72:@3678.4]
  assign _T_3264 = _T_3173 ? btb_hcount_25 : 2'h0; // @[Mux.scala 19:72:@3679.4]
  assign _T_3266 = _T_3174 ? btb_hcount_26 : 2'h0; // @[Mux.scala 19:72:@3680.4]
  assign _T_3268 = _T_3175 ? btb_hcount_27 : 2'h0; // @[Mux.scala 19:72:@3681.4]
  assign _T_3270 = _T_3176 ? btb_hcount_28 : 2'h0; // @[Mux.scala 19:72:@3682.4]
  assign _T_3272 = _T_3177 ? btb_hcount_29 : 2'h0; // @[Mux.scala 19:72:@3683.4]
  assign _T_3274 = _T_3178 ? btb_hcount_30 : 2'h0; // @[Mux.scala 19:72:@3684.4]
  assign _T_3276 = _T_3179 ? btb_hcount_31 : 2'h0; // @[Mux.scala 19:72:@3685.4]
  assign _T_3278 = _T_3180 ? btb_hcount_32 : 2'h0; // @[Mux.scala 19:72:@3686.4]
  assign _T_3280 = _T_3181 ? btb_hcount_33 : 2'h0; // @[Mux.scala 19:72:@3687.4]
  assign _T_3282 = _T_3182 ? btb_hcount_34 : 2'h0; // @[Mux.scala 19:72:@3688.4]
  assign _T_3284 = _T_3183 ? btb_hcount_35 : 2'h0; // @[Mux.scala 19:72:@3689.4]
  assign _T_3286 = _T_3184 ? btb_hcount_36 : 2'h0; // @[Mux.scala 19:72:@3690.4]
  assign _T_3288 = _T_3185 ? btb_hcount_37 : 2'h0; // @[Mux.scala 19:72:@3691.4]
  assign _T_3290 = _T_3186 ? btb_hcount_38 : 2'h0; // @[Mux.scala 19:72:@3692.4]
  assign _T_3292 = _T_3187 ? btb_hcount_39 : 2'h0; // @[Mux.scala 19:72:@3693.4]
  assign _T_3294 = _T_3188 ? btb_hcount_40 : 2'h0; // @[Mux.scala 19:72:@3694.4]
  assign _T_3296 = _T_3189 ? btb_hcount_41 : 2'h0; // @[Mux.scala 19:72:@3695.4]
  assign _T_3298 = _T_3190 ? btb_hcount_42 : 2'h0; // @[Mux.scala 19:72:@3696.4]
  assign _T_3300 = _T_3191 ? btb_hcount_43 : 2'h0; // @[Mux.scala 19:72:@3697.4]
  assign _T_3302 = _T_3192 ? btb_hcount_44 : 2'h0; // @[Mux.scala 19:72:@3698.4]
  assign _T_3304 = _T_3193 ? btb_hcount_45 : 2'h0; // @[Mux.scala 19:72:@3699.4]
  assign _T_3306 = _T_3194 ? btb_hcount_46 : 2'h0; // @[Mux.scala 19:72:@3700.4]
  assign _T_3308 = _T_3195 ? btb_hcount_47 : 2'h0; // @[Mux.scala 19:72:@3701.4]
  assign _T_3310 = _T_3196 ? btb_hcount_48 : 2'h0; // @[Mux.scala 19:72:@3702.4]
  assign _T_3312 = _T_3197 ? btb_hcount_49 : 2'h0; // @[Mux.scala 19:72:@3703.4]
  assign _T_3314 = _T_3198 ? btb_hcount_50 : 2'h0; // @[Mux.scala 19:72:@3704.4]
  assign _T_3316 = _T_3199 ? btb_hcount_51 : 2'h0; // @[Mux.scala 19:72:@3705.4]
  assign _T_3318 = _T_3200 ? btb_hcount_52 : 2'h0; // @[Mux.scala 19:72:@3706.4]
  assign _T_3320 = _T_3201 ? btb_hcount_53 : 2'h0; // @[Mux.scala 19:72:@3707.4]
  assign _T_3322 = _T_3202 ? btb_hcount_54 : 2'h0; // @[Mux.scala 19:72:@3708.4]
  assign _T_3324 = _T_3203 ? btb_hcount_55 : 2'h0; // @[Mux.scala 19:72:@3709.4]
  assign _T_3326 = _T_3204 ? btb_hcount_56 : 2'h0; // @[Mux.scala 19:72:@3710.4]
  assign _T_3328 = _T_3205 ? btb_hcount_57 : 2'h0; // @[Mux.scala 19:72:@3711.4]
  assign _T_3330 = _T_3206 ? btb_hcount_58 : 2'h0; // @[Mux.scala 19:72:@3712.4]
  assign _T_3332 = _T_3207 ? btb_hcount_59 : 2'h0; // @[Mux.scala 19:72:@3713.4]
  assign _T_3334 = _T_3208 ? btb_hcount_60 : 2'h0; // @[Mux.scala 19:72:@3714.4]
  assign _T_3336 = _T_3209 ? btb_hcount_61 : 2'h0; // @[Mux.scala 19:72:@3715.4]
  assign _T_3338 = _T_3210 ? btb_hcount_62 : 2'h0; // @[Mux.scala 19:72:@3716.4]
  assign _T_3340 = _T_3211 ? btb_hcount_63 : 2'h0; // @[Mux.scala 19:72:@3717.4]
  assign _T_3341 = _T_3214 | _T_3216; // @[Mux.scala 19:72:@3718.4]
  assign _T_3342 = _T_3341 | _T_3218; // @[Mux.scala 19:72:@3719.4]
  assign _T_3343 = _T_3342 | _T_3220; // @[Mux.scala 19:72:@3720.4]
  assign _T_3344 = _T_3343 | _T_3222; // @[Mux.scala 19:72:@3721.4]
  assign _T_3345 = _T_3344 | _T_3224; // @[Mux.scala 19:72:@3722.4]
  assign _T_3346 = _T_3345 | _T_3226; // @[Mux.scala 19:72:@3723.4]
  assign _T_3347 = _T_3346 | _T_3228; // @[Mux.scala 19:72:@3724.4]
  assign _T_3348 = _T_3347 | _T_3230; // @[Mux.scala 19:72:@3725.4]
  assign _T_3349 = _T_3348 | _T_3232; // @[Mux.scala 19:72:@3726.4]
  assign _T_3350 = _T_3349 | _T_3234; // @[Mux.scala 19:72:@3727.4]
  assign _T_3351 = _T_3350 | _T_3236; // @[Mux.scala 19:72:@3728.4]
  assign _T_3352 = _T_3351 | _T_3238; // @[Mux.scala 19:72:@3729.4]
  assign _T_3353 = _T_3352 | _T_3240; // @[Mux.scala 19:72:@3730.4]
  assign _T_3354 = _T_3353 | _T_3242; // @[Mux.scala 19:72:@3731.4]
  assign _T_3355 = _T_3354 | _T_3244; // @[Mux.scala 19:72:@3732.4]
  assign _T_3356 = _T_3355 | _T_3246; // @[Mux.scala 19:72:@3733.4]
  assign _T_3357 = _T_3356 | _T_3248; // @[Mux.scala 19:72:@3734.4]
  assign _T_3358 = _T_3357 | _T_3250; // @[Mux.scala 19:72:@3735.4]
  assign _T_3359 = _T_3358 | _T_3252; // @[Mux.scala 19:72:@3736.4]
  assign _T_3360 = _T_3359 | _T_3254; // @[Mux.scala 19:72:@3737.4]
  assign _T_3361 = _T_3360 | _T_3256; // @[Mux.scala 19:72:@3738.4]
  assign _T_3362 = _T_3361 | _T_3258; // @[Mux.scala 19:72:@3739.4]
  assign _T_3363 = _T_3362 | _T_3260; // @[Mux.scala 19:72:@3740.4]
  assign _T_3364 = _T_3363 | _T_3262; // @[Mux.scala 19:72:@3741.4]
  assign _T_3365 = _T_3364 | _T_3264; // @[Mux.scala 19:72:@3742.4]
  assign _T_3366 = _T_3365 | _T_3266; // @[Mux.scala 19:72:@3743.4]
  assign _T_3367 = _T_3366 | _T_3268; // @[Mux.scala 19:72:@3744.4]
  assign _T_3368 = _T_3367 | _T_3270; // @[Mux.scala 19:72:@3745.4]
  assign _T_3369 = _T_3368 | _T_3272; // @[Mux.scala 19:72:@3746.4]
  assign _T_3370 = _T_3369 | _T_3274; // @[Mux.scala 19:72:@3747.4]
  assign _T_3371 = _T_3370 | _T_3276; // @[Mux.scala 19:72:@3748.4]
  assign _T_3372 = _T_3371 | _T_3278; // @[Mux.scala 19:72:@3749.4]
  assign _T_3373 = _T_3372 | _T_3280; // @[Mux.scala 19:72:@3750.4]
  assign _T_3374 = _T_3373 | _T_3282; // @[Mux.scala 19:72:@3751.4]
  assign _T_3375 = _T_3374 | _T_3284; // @[Mux.scala 19:72:@3752.4]
  assign _T_3376 = _T_3375 | _T_3286; // @[Mux.scala 19:72:@3753.4]
  assign _T_3377 = _T_3376 | _T_3288; // @[Mux.scala 19:72:@3754.4]
  assign _T_3378 = _T_3377 | _T_3290; // @[Mux.scala 19:72:@3755.4]
  assign _T_3379 = _T_3378 | _T_3292; // @[Mux.scala 19:72:@3756.4]
  assign _T_3380 = _T_3379 | _T_3294; // @[Mux.scala 19:72:@3757.4]
  assign _T_3381 = _T_3380 | _T_3296; // @[Mux.scala 19:72:@3758.4]
  assign _T_3382 = _T_3381 | _T_3298; // @[Mux.scala 19:72:@3759.4]
  assign _T_3383 = _T_3382 | _T_3300; // @[Mux.scala 19:72:@3760.4]
  assign _T_3384 = _T_3383 | _T_3302; // @[Mux.scala 19:72:@3761.4]
  assign _T_3385 = _T_3384 | _T_3304; // @[Mux.scala 19:72:@3762.4]
  assign _T_3386 = _T_3385 | _T_3306; // @[Mux.scala 19:72:@3763.4]
  assign _T_3387 = _T_3386 | _T_3308; // @[Mux.scala 19:72:@3764.4]
  assign _T_3388 = _T_3387 | _T_3310; // @[Mux.scala 19:72:@3765.4]
  assign _T_3389 = _T_3388 | _T_3312; // @[Mux.scala 19:72:@3766.4]
  assign _T_3390 = _T_3389 | _T_3314; // @[Mux.scala 19:72:@3767.4]
  assign _T_3391 = _T_3390 | _T_3316; // @[Mux.scala 19:72:@3768.4]
  assign _T_3392 = _T_3391 | _T_3318; // @[Mux.scala 19:72:@3769.4]
  assign _T_3393 = _T_3392 | _T_3320; // @[Mux.scala 19:72:@3770.4]
  assign _T_3394 = _T_3393 | _T_3322; // @[Mux.scala 19:72:@3771.4]
  assign _T_3395 = _T_3394 | _T_3324; // @[Mux.scala 19:72:@3772.4]
  assign _T_3396 = _T_3395 | _T_3326; // @[Mux.scala 19:72:@3773.4]
  assign _T_3397 = _T_3396 | _T_3328; // @[Mux.scala 19:72:@3774.4]
  assign _T_3398 = _T_3397 | _T_3330; // @[Mux.scala 19:72:@3775.4]
  assign _T_3399 = _T_3398 | _T_3332; // @[Mux.scala 19:72:@3776.4]
  assign _T_3400 = _T_3399 | _T_3334; // @[Mux.scala 19:72:@3777.4]
  assign _T_3401 = _T_3400 | _T_3336; // @[Mux.scala 19:72:@3778.4]
  assign _T_3402 = _T_3401 | _T_3338; // @[Mux.scala 19:72:@3779.4]
  assign fb_wire_hcount = _T_3402 | _T_3340; // @[Mux.scala 19:72:@3780.4]
  assign _T_3407 = fb_wire_lookup != 64'h0; // @[BTB.scala 121:30:@3784.4]
  assign _T_3408 = fb_wire_lookup[63:32]; // @[OneHot.scala 26:18:@3785.4]
  assign _T_3409 = fb_wire_lookup[31:0]; // @[OneHot.scala 27:18:@3786.4]
  assign _T_3411 = _T_3408 != 32'h0; // @[OneHot.scala 28:14:@3787.4]
  assign _T_3412 = _T_3408 | _T_3409; // @[OneHot.scala 28:28:@3788.4]
  assign _T_3413 = _T_3412[31:16]; // @[OneHot.scala 26:18:@3789.4]
  assign _T_3414 = _T_3412[15:0]; // @[OneHot.scala 27:18:@3790.4]
  assign _T_3416 = _T_3413 != 16'h0; // @[OneHot.scala 28:14:@3791.4]
  assign _T_3417 = _T_3413 | _T_3414; // @[OneHot.scala 28:28:@3792.4]
  assign _T_3418 = _T_3417[15:8]; // @[OneHot.scala 26:18:@3793.4]
  assign _T_3419 = _T_3417[7:0]; // @[OneHot.scala 27:18:@3794.4]
  assign _T_3421 = _T_3418 != 8'h0; // @[OneHot.scala 28:14:@3795.4]
  assign _T_3422 = _T_3418 | _T_3419; // @[OneHot.scala 28:28:@3796.4]
  assign _T_3423 = _T_3422[7:4]; // @[OneHot.scala 26:18:@3797.4]
  assign _T_3424 = _T_3422[3:0]; // @[OneHot.scala 27:18:@3798.4]
  assign _T_3426 = _T_3423 != 4'h0; // @[OneHot.scala 28:14:@3799.4]
  assign _T_3427 = _T_3423 | _T_3424; // @[OneHot.scala 28:28:@3800.4]
  assign _T_3428 = _T_3427[3:2]; // @[OneHot.scala 26:18:@3801.4]
  assign _T_3429 = _T_3427[1:0]; // @[OneHot.scala 27:18:@3802.4]
  assign _T_3431 = _T_3428 != 2'h0; // @[OneHot.scala 28:14:@3803.4]
  assign _T_3432 = _T_3428 | _T_3429; // @[OneHot.scala 28:28:@3804.4]
  assign _T_3433 = _T_3432[1]; // @[CircuitMath.scala 30:8:@3805.4]
  assign _T_3438 = {_T_3411,_T_3416,_T_3421,_T_3426,_T_3431,_T_3433}; // @[Cat.scala 30:58:@3810.4]
  assign _T_3700 = ~ _T_614; // @[BTB.scala 127:21:@4003.4]
  assign _T_3702 = _T_3700 == 64'h0; // @[BTB.scala 127:21:@4004.4]
  assign _T_3965 = _T_3700[0]; // @[OneHot.scala 39:40:@4198.4]
  assign _T_3966 = _T_3700[1]; // @[OneHot.scala 39:40:@4199.4]
  assign _T_3967 = _T_3700[2]; // @[OneHot.scala 39:40:@4200.4]
  assign _T_3968 = _T_3700[3]; // @[OneHot.scala 39:40:@4201.4]
  assign _T_3969 = _T_3700[4]; // @[OneHot.scala 39:40:@4202.4]
  assign _T_3970 = _T_3700[5]; // @[OneHot.scala 39:40:@4203.4]
  assign _T_3971 = _T_3700[6]; // @[OneHot.scala 39:40:@4204.4]
  assign _T_3972 = _T_3700[7]; // @[OneHot.scala 39:40:@4205.4]
  assign _T_3973 = _T_3700[8]; // @[OneHot.scala 39:40:@4206.4]
  assign _T_3974 = _T_3700[9]; // @[OneHot.scala 39:40:@4207.4]
  assign _T_3975 = _T_3700[10]; // @[OneHot.scala 39:40:@4208.4]
  assign _T_3976 = _T_3700[11]; // @[OneHot.scala 39:40:@4209.4]
  assign _T_3977 = _T_3700[12]; // @[OneHot.scala 39:40:@4210.4]
  assign _T_3978 = _T_3700[13]; // @[OneHot.scala 39:40:@4211.4]
  assign _T_3979 = _T_3700[14]; // @[OneHot.scala 39:40:@4212.4]
  assign _T_3980 = _T_3700[15]; // @[OneHot.scala 39:40:@4213.4]
  assign _T_3981 = _T_3700[16]; // @[OneHot.scala 39:40:@4214.4]
  assign _T_3982 = _T_3700[17]; // @[OneHot.scala 39:40:@4215.4]
  assign _T_3983 = _T_3700[18]; // @[OneHot.scala 39:40:@4216.4]
  assign _T_3984 = _T_3700[19]; // @[OneHot.scala 39:40:@4217.4]
  assign _T_3985 = _T_3700[20]; // @[OneHot.scala 39:40:@4218.4]
  assign _T_3986 = _T_3700[21]; // @[OneHot.scala 39:40:@4219.4]
  assign _T_3987 = _T_3700[22]; // @[OneHot.scala 39:40:@4220.4]
  assign _T_3988 = _T_3700[23]; // @[OneHot.scala 39:40:@4221.4]
  assign _T_3989 = _T_3700[24]; // @[OneHot.scala 39:40:@4222.4]
  assign _T_3990 = _T_3700[25]; // @[OneHot.scala 39:40:@4223.4]
  assign _T_3991 = _T_3700[26]; // @[OneHot.scala 39:40:@4224.4]
  assign _T_3992 = _T_3700[27]; // @[OneHot.scala 39:40:@4225.4]
  assign _T_3993 = _T_3700[28]; // @[OneHot.scala 39:40:@4226.4]
  assign _T_3994 = _T_3700[29]; // @[OneHot.scala 39:40:@4227.4]
  assign _T_3995 = _T_3700[30]; // @[OneHot.scala 39:40:@4228.4]
  assign _T_3996 = _T_3700[31]; // @[OneHot.scala 39:40:@4229.4]
  assign _T_3997 = _T_3700[32]; // @[OneHot.scala 39:40:@4230.4]
  assign _T_3998 = _T_3700[33]; // @[OneHot.scala 39:40:@4231.4]
  assign _T_3999 = _T_3700[34]; // @[OneHot.scala 39:40:@4232.4]
  assign _T_4000 = _T_3700[35]; // @[OneHot.scala 39:40:@4233.4]
  assign _T_4001 = _T_3700[36]; // @[OneHot.scala 39:40:@4234.4]
  assign _T_4002 = _T_3700[37]; // @[OneHot.scala 39:40:@4235.4]
  assign _T_4003 = _T_3700[38]; // @[OneHot.scala 39:40:@4236.4]
  assign _T_4004 = _T_3700[39]; // @[OneHot.scala 39:40:@4237.4]
  assign _T_4005 = _T_3700[40]; // @[OneHot.scala 39:40:@4238.4]
  assign _T_4006 = _T_3700[41]; // @[OneHot.scala 39:40:@4239.4]
  assign _T_4007 = _T_3700[42]; // @[OneHot.scala 39:40:@4240.4]
  assign _T_4008 = _T_3700[43]; // @[OneHot.scala 39:40:@4241.4]
  assign _T_4009 = _T_3700[44]; // @[OneHot.scala 39:40:@4242.4]
  assign _T_4010 = _T_3700[45]; // @[OneHot.scala 39:40:@4243.4]
  assign _T_4011 = _T_3700[46]; // @[OneHot.scala 39:40:@4244.4]
  assign _T_4012 = _T_3700[47]; // @[OneHot.scala 39:40:@4245.4]
  assign _T_4013 = _T_3700[48]; // @[OneHot.scala 39:40:@4246.4]
  assign _T_4014 = _T_3700[49]; // @[OneHot.scala 39:40:@4247.4]
  assign _T_4015 = _T_3700[50]; // @[OneHot.scala 39:40:@4248.4]
  assign _T_4016 = _T_3700[51]; // @[OneHot.scala 39:40:@4249.4]
  assign _T_4017 = _T_3700[52]; // @[OneHot.scala 39:40:@4250.4]
  assign _T_4018 = _T_3700[53]; // @[OneHot.scala 39:40:@4251.4]
  assign _T_4019 = _T_3700[54]; // @[OneHot.scala 39:40:@4252.4]
  assign _T_4020 = _T_3700[55]; // @[OneHot.scala 39:40:@4253.4]
  assign _T_4021 = _T_3700[56]; // @[OneHot.scala 39:40:@4254.4]
  assign _T_4022 = _T_3700[57]; // @[OneHot.scala 39:40:@4255.4]
  assign _T_4023 = _T_3700[58]; // @[OneHot.scala 39:40:@4256.4]
  assign _T_4024 = _T_3700[59]; // @[OneHot.scala 39:40:@4257.4]
  assign _T_4025 = _T_3700[60]; // @[OneHot.scala 39:40:@4258.4]
  assign _T_4026 = _T_3700[61]; // @[OneHot.scala 39:40:@4259.4]
  assign _T_4027 = _T_3700[62]; // @[OneHot.scala 39:40:@4260.4]
  assign _T_4093 = _T_4027 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@4262.4]
  assign _T_4094 = _T_4026 ? 6'h3d : _T_4093; // @[Mux.scala 31:69:@4263.4]
  assign _T_4095 = _T_4025 ? 6'h3c : _T_4094; // @[Mux.scala 31:69:@4264.4]
  assign _T_4096 = _T_4024 ? 6'h3b : _T_4095; // @[Mux.scala 31:69:@4265.4]
  assign _T_4097 = _T_4023 ? 6'h3a : _T_4096; // @[Mux.scala 31:69:@4266.4]
  assign _T_4098 = _T_4022 ? 6'h39 : _T_4097; // @[Mux.scala 31:69:@4267.4]
  assign _T_4099 = _T_4021 ? 6'h38 : _T_4098; // @[Mux.scala 31:69:@4268.4]
  assign _T_4100 = _T_4020 ? 6'h37 : _T_4099; // @[Mux.scala 31:69:@4269.4]
  assign _T_4101 = _T_4019 ? 6'h36 : _T_4100; // @[Mux.scala 31:69:@4270.4]
  assign _T_4102 = _T_4018 ? 6'h35 : _T_4101; // @[Mux.scala 31:69:@4271.4]
  assign _T_4103 = _T_4017 ? 6'h34 : _T_4102; // @[Mux.scala 31:69:@4272.4]
  assign _T_4104 = _T_4016 ? 6'h33 : _T_4103; // @[Mux.scala 31:69:@4273.4]
  assign _T_4105 = _T_4015 ? 6'h32 : _T_4104; // @[Mux.scala 31:69:@4274.4]
  assign _T_4106 = _T_4014 ? 6'h31 : _T_4105; // @[Mux.scala 31:69:@4275.4]
  assign _T_4107 = _T_4013 ? 6'h30 : _T_4106; // @[Mux.scala 31:69:@4276.4]
  assign _T_4108 = _T_4012 ? 6'h2f : _T_4107; // @[Mux.scala 31:69:@4277.4]
  assign _T_4109 = _T_4011 ? 6'h2e : _T_4108; // @[Mux.scala 31:69:@4278.4]
  assign _T_4110 = _T_4010 ? 6'h2d : _T_4109; // @[Mux.scala 31:69:@4279.4]
  assign _T_4111 = _T_4009 ? 6'h2c : _T_4110; // @[Mux.scala 31:69:@4280.4]
  assign _T_4112 = _T_4008 ? 6'h2b : _T_4111; // @[Mux.scala 31:69:@4281.4]
  assign _T_4113 = _T_4007 ? 6'h2a : _T_4112; // @[Mux.scala 31:69:@4282.4]
  assign _T_4114 = _T_4006 ? 6'h29 : _T_4113; // @[Mux.scala 31:69:@4283.4]
  assign _T_4115 = _T_4005 ? 6'h28 : _T_4114; // @[Mux.scala 31:69:@4284.4]
  assign _T_4116 = _T_4004 ? 6'h27 : _T_4115; // @[Mux.scala 31:69:@4285.4]
  assign _T_4117 = _T_4003 ? 6'h26 : _T_4116; // @[Mux.scala 31:69:@4286.4]
  assign _T_4118 = _T_4002 ? 6'h25 : _T_4117; // @[Mux.scala 31:69:@4287.4]
  assign _T_4119 = _T_4001 ? 6'h24 : _T_4118; // @[Mux.scala 31:69:@4288.4]
  assign _T_4120 = _T_4000 ? 6'h23 : _T_4119; // @[Mux.scala 31:69:@4289.4]
  assign _T_4121 = _T_3999 ? 6'h22 : _T_4120; // @[Mux.scala 31:69:@4290.4]
  assign _T_4122 = _T_3998 ? 6'h21 : _T_4121; // @[Mux.scala 31:69:@4291.4]
  assign _T_4123 = _T_3997 ? 6'h20 : _T_4122; // @[Mux.scala 31:69:@4292.4]
  assign _T_4124 = _T_3996 ? 6'h1f : _T_4123; // @[Mux.scala 31:69:@4293.4]
  assign _T_4125 = _T_3995 ? 6'h1e : _T_4124; // @[Mux.scala 31:69:@4294.4]
  assign _T_4126 = _T_3994 ? 6'h1d : _T_4125; // @[Mux.scala 31:69:@4295.4]
  assign _T_4127 = _T_3993 ? 6'h1c : _T_4126; // @[Mux.scala 31:69:@4296.4]
  assign _T_4128 = _T_3992 ? 6'h1b : _T_4127; // @[Mux.scala 31:69:@4297.4]
  assign _T_4129 = _T_3991 ? 6'h1a : _T_4128; // @[Mux.scala 31:69:@4298.4]
  assign _T_4130 = _T_3990 ? 6'h19 : _T_4129; // @[Mux.scala 31:69:@4299.4]
  assign _T_4131 = _T_3989 ? 6'h18 : _T_4130; // @[Mux.scala 31:69:@4300.4]
  assign _T_4132 = _T_3988 ? 6'h17 : _T_4131; // @[Mux.scala 31:69:@4301.4]
  assign _T_4133 = _T_3987 ? 6'h16 : _T_4132; // @[Mux.scala 31:69:@4302.4]
  assign _T_4134 = _T_3986 ? 6'h15 : _T_4133; // @[Mux.scala 31:69:@4303.4]
  assign _T_4135 = _T_3985 ? 6'h14 : _T_4134; // @[Mux.scala 31:69:@4304.4]
  assign _T_4136 = _T_3984 ? 6'h13 : _T_4135; // @[Mux.scala 31:69:@4305.4]
  assign _T_4137 = _T_3983 ? 6'h12 : _T_4136; // @[Mux.scala 31:69:@4306.4]
  assign _T_4138 = _T_3982 ? 6'h11 : _T_4137; // @[Mux.scala 31:69:@4307.4]
  assign _T_4139 = _T_3981 ? 6'h10 : _T_4138; // @[Mux.scala 31:69:@4308.4]
  assign _T_4140 = _T_3980 ? 6'hf : _T_4139; // @[Mux.scala 31:69:@4309.4]
  assign _T_4141 = _T_3979 ? 6'he : _T_4140; // @[Mux.scala 31:69:@4310.4]
  assign _T_4142 = _T_3978 ? 6'hd : _T_4141; // @[Mux.scala 31:69:@4311.4]
  assign _T_4143 = _T_3977 ? 6'hc : _T_4142; // @[Mux.scala 31:69:@4312.4]
  assign _T_4144 = _T_3976 ? 6'hb : _T_4143; // @[Mux.scala 31:69:@4313.4]
  assign _T_4145 = _T_3975 ? 6'ha : _T_4144; // @[Mux.scala 31:69:@4314.4]
  assign _T_4146 = _T_3974 ? 6'h9 : _T_4145; // @[Mux.scala 31:69:@4315.4]
  assign _T_4147 = _T_3973 ? 6'h8 : _T_4146; // @[Mux.scala 31:69:@4316.4]
  assign _T_4148 = _T_3972 ? 6'h7 : _T_4147; // @[Mux.scala 31:69:@4317.4]
  assign _T_4149 = _T_3971 ? 6'h6 : _T_4148; // @[Mux.scala 31:69:@4318.4]
  assign _T_4150 = _T_3970 ? 6'h5 : _T_4149; // @[Mux.scala 31:69:@4319.4]
  assign _T_4151 = _T_3969 ? 6'h4 : _T_4150; // @[Mux.scala 31:69:@4320.4]
  assign _T_4152 = _T_3968 ? 6'h3 : _T_4151; // @[Mux.scala 31:69:@4321.4]
  assign _T_4153 = _T_3967 ? 6'h2 : _T_4152; // @[Mux.scala 31:69:@4322.4]
  assign _T_4154 = _T_3966 ? 6'h1 : _T_4153; // @[Mux.scala 31:69:@4323.4]
  assign _T_4155 = _T_3965 ? 6'h0 : _T_4154; // @[Mux.scala 31:69:@4324.4]
  assign _T_4156 = _T_3702 ? fb_reg_lfsr : _T_4155; // @[BTB.scala 127:10:@4325.4]
  assign fb_wire_bindex = _T_3407 ? _T_3438 : _T_4156; // @[BTB.scala 126:8:@4326.4]
  assign _GEN_0 = 6'h0 == fb_wire_bindex ? fb_reg_pc : btb_pc_0; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_1 = 6'h1 == fb_wire_bindex ? fb_reg_pc : btb_pc_1; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_2 = 6'h2 == fb_wire_bindex ? fb_reg_pc : btb_pc_2; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_3 = 6'h3 == fb_wire_bindex ? fb_reg_pc : btb_pc_3; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_4 = 6'h4 == fb_wire_bindex ? fb_reg_pc : btb_pc_4; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_5 = 6'h5 == fb_wire_bindex ? fb_reg_pc : btb_pc_5; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_6 = 6'h6 == fb_wire_bindex ? fb_reg_pc : btb_pc_6; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_7 = 6'h7 == fb_wire_bindex ? fb_reg_pc : btb_pc_7; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_8 = 6'h8 == fb_wire_bindex ? fb_reg_pc : btb_pc_8; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_9 = 6'h9 == fb_wire_bindex ? fb_reg_pc : btb_pc_9; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_10 = 6'ha == fb_wire_bindex ? fb_reg_pc : btb_pc_10; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_11 = 6'hb == fb_wire_bindex ? fb_reg_pc : btb_pc_11; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_12 = 6'hc == fb_wire_bindex ? fb_reg_pc : btb_pc_12; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_13 = 6'hd == fb_wire_bindex ? fb_reg_pc : btb_pc_13; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_14 = 6'he == fb_wire_bindex ? fb_reg_pc : btb_pc_14; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_15 = 6'hf == fb_wire_bindex ? fb_reg_pc : btb_pc_15; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_16 = 6'h10 == fb_wire_bindex ? fb_reg_pc : btb_pc_16; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_17 = 6'h11 == fb_wire_bindex ? fb_reg_pc : btb_pc_17; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_18 = 6'h12 == fb_wire_bindex ? fb_reg_pc : btb_pc_18; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_19 = 6'h13 == fb_wire_bindex ? fb_reg_pc : btb_pc_19; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_20 = 6'h14 == fb_wire_bindex ? fb_reg_pc : btb_pc_20; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_21 = 6'h15 == fb_wire_bindex ? fb_reg_pc : btb_pc_21; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_22 = 6'h16 == fb_wire_bindex ? fb_reg_pc : btb_pc_22; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_23 = 6'h17 == fb_wire_bindex ? fb_reg_pc : btb_pc_23; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_24 = 6'h18 == fb_wire_bindex ? fb_reg_pc : btb_pc_24; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_25 = 6'h19 == fb_wire_bindex ? fb_reg_pc : btb_pc_25; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_26 = 6'h1a == fb_wire_bindex ? fb_reg_pc : btb_pc_26; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_27 = 6'h1b == fb_wire_bindex ? fb_reg_pc : btb_pc_27; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_28 = 6'h1c == fb_wire_bindex ? fb_reg_pc : btb_pc_28; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_29 = 6'h1d == fb_wire_bindex ? fb_reg_pc : btb_pc_29; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_30 = 6'h1e == fb_wire_bindex ? fb_reg_pc : btb_pc_30; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_31 = 6'h1f == fb_wire_bindex ? fb_reg_pc : btb_pc_31; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_32 = 6'h20 == fb_wire_bindex ? fb_reg_pc : btb_pc_32; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_33 = 6'h21 == fb_wire_bindex ? fb_reg_pc : btb_pc_33; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_34 = 6'h22 == fb_wire_bindex ? fb_reg_pc : btb_pc_34; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_35 = 6'h23 == fb_wire_bindex ? fb_reg_pc : btb_pc_35; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_36 = 6'h24 == fb_wire_bindex ? fb_reg_pc : btb_pc_36; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_37 = 6'h25 == fb_wire_bindex ? fb_reg_pc : btb_pc_37; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_38 = 6'h26 == fb_wire_bindex ? fb_reg_pc : btb_pc_38; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_39 = 6'h27 == fb_wire_bindex ? fb_reg_pc : btb_pc_39; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_40 = 6'h28 == fb_wire_bindex ? fb_reg_pc : btb_pc_40; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_41 = 6'h29 == fb_wire_bindex ? fb_reg_pc : btb_pc_41; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_42 = 6'h2a == fb_wire_bindex ? fb_reg_pc : btb_pc_42; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_43 = 6'h2b == fb_wire_bindex ? fb_reg_pc : btb_pc_43; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_44 = 6'h2c == fb_wire_bindex ? fb_reg_pc : btb_pc_44; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_45 = 6'h2d == fb_wire_bindex ? fb_reg_pc : btb_pc_45; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_46 = 6'h2e == fb_wire_bindex ? fb_reg_pc : btb_pc_46; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_47 = 6'h2f == fb_wire_bindex ? fb_reg_pc : btb_pc_47; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_48 = 6'h30 == fb_wire_bindex ? fb_reg_pc : btb_pc_48; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_49 = 6'h31 == fb_wire_bindex ? fb_reg_pc : btb_pc_49; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_50 = 6'h32 == fb_wire_bindex ? fb_reg_pc : btb_pc_50; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_51 = 6'h33 == fb_wire_bindex ? fb_reg_pc : btb_pc_51; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_52 = 6'h34 == fb_wire_bindex ? fb_reg_pc : btb_pc_52; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_53 = 6'h35 == fb_wire_bindex ? fb_reg_pc : btb_pc_53; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_54 = 6'h36 == fb_wire_bindex ? fb_reg_pc : btb_pc_54; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_55 = 6'h37 == fb_wire_bindex ? fb_reg_pc : btb_pc_55; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_56 = 6'h38 == fb_wire_bindex ? fb_reg_pc : btb_pc_56; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_57 = 6'h39 == fb_wire_bindex ? fb_reg_pc : btb_pc_57; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_58 = 6'h3a == fb_wire_bindex ? fb_reg_pc : btb_pc_58; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_59 = 6'h3b == fb_wire_bindex ? fb_reg_pc : btb_pc_59; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_60 = 6'h3c == fb_wire_bindex ? fb_reg_pc : btb_pc_60; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_61 = 6'h3d == fb_wire_bindex ? fb_reg_pc : btb_pc_61; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_62 = 6'h3e == fb_wire_bindex ? fb_reg_pc : btb_pc_62; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_63 = 6'h3f == fb_wire_bindex ? fb_reg_pc : btb_pc_63; // @[BTB.scala 132:34:@4330.8]
  assign _GEN_64 = 6'h0 == fb_wire_bindex ? fb_reg_target : btb_target_0; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_65 = 6'h1 == fb_wire_bindex ? fb_reg_target : btb_target_1; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_66 = 6'h2 == fb_wire_bindex ? fb_reg_target : btb_target_2; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_67 = 6'h3 == fb_wire_bindex ? fb_reg_target : btb_target_3; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_68 = 6'h4 == fb_wire_bindex ? fb_reg_target : btb_target_4; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_69 = 6'h5 == fb_wire_bindex ? fb_reg_target : btb_target_5; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_70 = 6'h6 == fb_wire_bindex ? fb_reg_target : btb_target_6; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_71 = 6'h7 == fb_wire_bindex ? fb_reg_target : btb_target_7; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_72 = 6'h8 == fb_wire_bindex ? fb_reg_target : btb_target_8; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_73 = 6'h9 == fb_wire_bindex ? fb_reg_target : btb_target_9; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_74 = 6'ha == fb_wire_bindex ? fb_reg_target : btb_target_10; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_75 = 6'hb == fb_wire_bindex ? fb_reg_target : btb_target_11; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_76 = 6'hc == fb_wire_bindex ? fb_reg_target : btb_target_12; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_77 = 6'hd == fb_wire_bindex ? fb_reg_target : btb_target_13; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_78 = 6'he == fb_wire_bindex ? fb_reg_target : btb_target_14; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_79 = 6'hf == fb_wire_bindex ? fb_reg_target : btb_target_15; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_80 = 6'h10 == fb_wire_bindex ? fb_reg_target : btb_target_16; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_81 = 6'h11 == fb_wire_bindex ? fb_reg_target : btb_target_17; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_82 = 6'h12 == fb_wire_bindex ? fb_reg_target : btb_target_18; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_83 = 6'h13 == fb_wire_bindex ? fb_reg_target : btb_target_19; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_84 = 6'h14 == fb_wire_bindex ? fb_reg_target : btb_target_20; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_85 = 6'h15 == fb_wire_bindex ? fb_reg_target : btb_target_21; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_86 = 6'h16 == fb_wire_bindex ? fb_reg_target : btb_target_22; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_87 = 6'h17 == fb_wire_bindex ? fb_reg_target : btb_target_23; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_88 = 6'h18 == fb_wire_bindex ? fb_reg_target : btb_target_24; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_89 = 6'h19 == fb_wire_bindex ? fb_reg_target : btb_target_25; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_90 = 6'h1a == fb_wire_bindex ? fb_reg_target : btb_target_26; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_91 = 6'h1b == fb_wire_bindex ? fb_reg_target : btb_target_27; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_92 = 6'h1c == fb_wire_bindex ? fb_reg_target : btb_target_28; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_93 = 6'h1d == fb_wire_bindex ? fb_reg_target : btb_target_29; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_94 = 6'h1e == fb_wire_bindex ? fb_reg_target : btb_target_30; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_95 = 6'h1f == fb_wire_bindex ? fb_reg_target : btb_target_31; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_96 = 6'h20 == fb_wire_bindex ? fb_reg_target : btb_target_32; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_97 = 6'h21 == fb_wire_bindex ? fb_reg_target : btb_target_33; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_98 = 6'h22 == fb_wire_bindex ? fb_reg_target : btb_target_34; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_99 = 6'h23 == fb_wire_bindex ? fb_reg_target : btb_target_35; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_100 = 6'h24 == fb_wire_bindex ? fb_reg_target : btb_target_36; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_101 = 6'h25 == fb_wire_bindex ? fb_reg_target : btb_target_37; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_102 = 6'h26 == fb_wire_bindex ? fb_reg_target : btb_target_38; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_103 = 6'h27 == fb_wire_bindex ? fb_reg_target : btb_target_39; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_104 = 6'h28 == fb_wire_bindex ? fb_reg_target : btb_target_40; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_105 = 6'h29 == fb_wire_bindex ? fb_reg_target : btb_target_41; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_106 = 6'h2a == fb_wire_bindex ? fb_reg_target : btb_target_42; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_107 = 6'h2b == fb_wire_bindex ? fb_reg_target : btb_target_43; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_108 = 6'h2c == fb_wire_bindex ? fb_reg_target : btb_target_44; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_109 = 6'h2d == fb_wire_bindex ? fb_reg_target : btb_target_45; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_110 = 6'h2e == fb_wire_bindex ? fb_reg_target : btb_target_46; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_111 = 6'h2f == fb_wire_bindex ? fb_reg_target : btb_target_47; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_112 = 6'h30 == fb_wire_bindex ? fb_reg_target : btb_target_48; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_113 = 6'h31 == fb_wire_bindex ? fb_reg_target : btb_target_49; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_114 = 6'h32 == fb_wire_bindex ? fb_reg_target : btb_target_50; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_115 = 6'h33 == fb_wire_bindex ? fb_reg_target : btb_target_51; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_116 = 6'h34 == fb_wire_bindex ? fb_reg_target : btb_target_52; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_117 = 6'h35 == fb_wire_bindex ? fb_reg_target : btb_target_53; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_118 = 6'h36 == fb_wire_bindex ? fb_reg_target : btb_target_54; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_119 = 6'h37 == fb_wire_bindex ? fb_reg_target : btb_target_55; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_120 = 6'h38 == fb_wire_bindex ? fb_reg_target : btb_target_56; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_121 = 6'h39 == fb_wire_bindex ? fb_reg_target : btb_target_57; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_122 = 6'h3a == fb_wire_bindex ? fb_reg_target : btb_target_58; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_123 = 6'h3b == fb_wire_bindex ? fb_reg_target : btb_target_59; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_124 = 6'h3c == fb_wire_bindex ? fb_reg_target : btb_target_60; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_125 = 6'h3d == fb_wire_bindex ? fb_reg_target : btb_target_61; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_126 = 6'h3e == fb_wire_bindex ? fb_reg_target : btb_target_62; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_127 = 6'h3f == fb_wire_bindex ? fb_reg_target : btb_target_63; // @[BTB.scala 133:34:@4331.8]
  assign _GEN_128 = 6'h0 == fb_wire_bindex ? fb_reg_btype : btb_btype_0; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_129 = 6'h1 == fb_wire_bindex ? fb_reg_btype : btb_btype_1; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_130 = 6'h2 == fb_wire_bindex ? fb_reg_btype : btb_btype_2; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_131 = 6'h3 == fb_wire_bindex ? fb_reg_btype : btb_btype_3; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_132 = 6'h4 == fb_wire_bindex ? fb_reg_btype : btb_btype_4; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_133 = 6'h5 == fb_wire_bindex ? fb_reg_btype : btb_btype_5; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_134 = 6'h6 == fb_wire_bindex ? fb_reg_btype : btb_btype_6; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_135 = 6'h7 == fb_wire_bindex ? fb_reg_btype : btb_btype_7; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_136 = 6'h8 == fb_wire_bindex ? fb_reg_btype : btb_btype_8; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_137 = 6'h9 == fb_wire_bindex ? fb_reg_btype : btb_btype_9; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_138 = 6'ha == fb_wire_bindex ? fb_reg_btype : btb_btype_10; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_139 = 6'hb == fb_wire_bindex ? fb_reg_btype : btb_btype_11; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_140 = 6'hc == fb_wire_bindex ? fb_reg_btype : btb_btype_12; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_141 = 6'hd == fb_wire_bindex ? fb_reg_btype : btb_btype_13; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_142 = 6'he == fb_wire_bindex ? fb_reg_btype : btb_btype_14; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_143 = 6'hf == fb_wire_bindex ? fb_reg_btype : btb_btype_15; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_144 = 6'h10 == fb_wire_bindex ? fb_reg_btype : btb_btype_16; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_145 = 6'h11 == fb_wire_bindex ? fb_reg_btype : btb_btype_17; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_146 = 6'h12 == fb_wire_bindex ? fb_reg_btype : btb_btype_18; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_147 = 6'h13 == fb_wire_bindex ? fb_reg_btype : btb_btype_19; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_148 = 6'h14 == fb_wire_bindex ? fb_reg_btype : btb_btype_20; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_149 = 6'h15 == fb_wire_bindex ? fb_reg_btype : btb_btype_21; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_150 = 6'h16 == fb_wire_bindex ? fb_reg_btype : btb_btype_22; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_151 = 6'h17 == fb_wire_bindex ? fb_reg_btype : btb_btype_23; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_152 = 6'h18 == fb_wire_bindex ? fb_reg_btype : btb_btype_24; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_153 = 6'h19 == fb_wire_bindex ? fb_reg_btype : btb_btype_25; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_154 = 6'h1a == fb_wire_bindex ? fb_reg_btype : btb_btype_26; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_155 = 6'h1b == fb_wire_bindex ? fb_reg_btype : btb_btype_27; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_156 = 6'h1c == fb_wire_bindex ? fb_reg_btype : btb_btype_28; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_157 = 6'h1d == fb_wire_bindex ? fb_reg_btype : btb_btype_29; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_158 = 6'h1e == fb_wire_bindex ? fb_reg_btype : btb_btype_30; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_159 = 6'h1f == fb_wire_bindex ? fb_reg_btype : btb_btype_31; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_160 = 6'h20 == fb_wire_bindex ? fb_reg_btype : btb_btype_32; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_161 = 6'h21 == fb_wire_bindex ? fb_reg_btype : btb_btype_33; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_162 = 6'h22 == fb_wire_bindex ? fb_reg_btype : btb_btype_34; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_163 = 6'h23 == fb_wire_bindex ? fb_reg_btype : btb_btype_35; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_164 = 6'h24 == fb_wire_bindex ? fb_reg_btype : btb_btype_36; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_165 = 6'h25 == fb_wire_bindex ? fb_reg_btype : btb_btype_37; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_166 = 6'h26 == fb_wire_bindex ? fb_reg_btype : btb_btype_38; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_167 = 6'h27 == fb_wire_bindex ? fb_reg_btype : btb_btype_39; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_168 = 6'h28 == fb_wire_bindex ? fb_reg_btype : btb_btype_40; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_169 = 6'h29 == fb_wire_bindex ? fb_reg_btype : btb_btype_41; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_170 = 6'h2a == fb_wire_bindex ? fb_reg_btype : btb_btype_42; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_171 = 6'h2b == fb_wire_bindex ? fb_reg_btype : btb_btype_43; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_172 = 6'h2c == fb_wire_bindex ? fb_reg_btype : btb_btype_44; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_173 = 6'h2d == fb_wire_bindex ? fb_reg_btype : btb_btype_45; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_174 = 6'h2e == fb_wire_bindex ? fb_reg_btype : btb_btype_46; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_175 = 6'h2f == fb_wire_bindex ? fb_reg_btype : btb_btype_47; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_176 = 6'h30 == fb_wire_bindex ? fb_reg_btype : btb_btype_48; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_177 = 6'h31 == fb_wire_bindex ? fb_reg_btype : btb_btype_49; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_178 = 6'h32 == fb_wire_bindex ? fb_reg_btype : btb_btype_50; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_179 = 6'h33 == fb_wire_bindex ? fb_reg_btype : btb_btype_51; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_180 = 6'h34 == fb_wire_bindex ? fb_reg_btype : btb_btype_52; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_181 = 6'h35 == fb_wire_bindex ? fb_reg_btype : btb_btype_53; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_182 = 6'h36 == fb_wire_bindex ? fb_reg_btype : btb_btype_54; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_183 = 6'h37 == fb_wire_bindex ? fb_reg_btype : btb_btype_55; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_184 = 6'h38 == fb_wire_bindex ? fb_reg_btype : btb_btype_56; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_185 = 6'h39 == fb_wire_bindex ? fb_reg_btype : btb_btype_57; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_186 = 6'h3a == fb_wire_bindex ? fb_reg_btype : btb_btype_58; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_187 = 6'h3b == fb_wire_bindex ? fb_reg_btype : btb_btype_59; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_188 = 6'h3c == fb_wire_bindex ? fb_reg_btype : btb_btype_60; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_189 = 6'h3d == fb_wire_bindex ? fb_reg_btype : btb_btype_61; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_190 = 6'h3e == fb_wire_bindex ? fb_reg_btype : btb_btype_62; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_191 = 6'h3f == fb_wire_bindex ? fb_reg_btype : btb_btype_63; // @[BTB.scala 134:34:@4332.8]
  assign _GEN_192 = fb_reg_redirect ? _GEN_0 : btb_pc_0; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_193 = fb_reg_redirect ? _GEN_1 : btb_pc_1; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_194 = fb_reg_redirect ? _GEN_2 : btb_pc_2; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_195 = fb_reg_redirect ? _GEN_3 : btb_pc_3; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_196 = fb_reg_redirect ? _GEN_4 : btb_pc_4; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_197 = fb_reg_redirect ? _GEN_5 : btb_pc_5; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_198 = fb_reg_redirect ? _GEN_6 : btb_pc_6; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_199 = fb_reg_redirect ? _GEN_7 : btb_pc_7; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_200 = fb_reg_redirect ? _GEN_8 : btb_pc_8; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_201 = fb_reg_redirect ? _GEN_9 : btb_pc_9; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_202 = fb_reg_redirect ? _GEN_10 : btb_pc_10; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_203 = fb_reg_redirect ? _GEN_11 : btb_pc_11; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_204 = fb_reg_redirect ? _GEN_12 : btb_pc_12; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_205 = fb_reg_redirect ? _GEN_13 : btb_pc_13; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_206 = fb_reg_redirect ? _GEN_14 : btb_pc_14; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_207 = fb_reg_redirect ? _GEN_15 : btb_pc_15; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_208 = fb_reg_redirect ? _GEN_16 : btb_pc_16; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_209 = fb_reg_redirect ? _GEN_17 : btb_pc_17; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_210 = fb_reg_redirect ? _GEN_18 : btb_pc_18; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_211 = fb_reg_redirect ? _GEN_19 : btb_pc_19; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_212 = fb_reg_redirect ? _GEN_20 : btb_pc_20; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_213 = fb_reg_redirect ? _GEN_21 : btb_pc_21; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_214 = fb_reg_redirect ? _GEN_22 : btb_pc_22; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_215 = fb_reg_redirect ? _GEN_23 : btb_pc_23; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_216 = fb_reg_redirect ? _GEN_24 : btb_pc_24; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_217 = fb_reg_redirect ? _GEN_25 : btb_pc_25; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_218 = fb_reg_redirect ? _GEN_26 : btb_pc_26; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_219 = fb_reg_redirect ? _GEN_27 : btb_pc_27; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_220 = fb_reg_redirect ? _GEN_28 : btb_pc_28; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_221 = fb_reg_redirect ? _GEN_29 : btb_pc_29; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_222 = fb_reg_redirect ? _GEN_30 : btb_pc_30; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_223 = fb_reg_redirect ? _GEN_31 : btb_pc_31; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_224 = fb_reg_redirect ? _GEN_32 : btb_pc_32; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_225 = fb_reg_redirect ? _GEN_33 : btb_pc_33; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_226 = fb_reg_redirect ? _GEN_34 : btb_pc_34; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_227 = fb_reg_redirect ? _GEN_35 : btb_pc_35; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_228 = fb_reg_redirect ? _GEN_36 : btb_pc_36; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_229 = fb_reg_redirect ? _GEN_37 : btb_pc_37; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_230 = fb_reg_redirect ? _GEN_38 : btb_pc_38; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_231 = fb_reg_redirect ? _GEN_39 : btb_pc_39; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_232 = fb_reg_redirect ? _GEN_40 : btb_pc_40; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_233 = fb_reg_redirect ? _GEN_41 : btb_pc_41; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_234 = fb_reg_redirect ? _GEN_42 : btb_pc_42; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_235 = fb_reg_redirect ? _GEN_43 : btb_pc_43; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_236 = fb_reg_redirect ? _GEN_44 : btb_pc_44; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_237 = fb_reg_redirect ? _GEN_45 : btb_pc_45; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_238 = fb_reg_redirect ? _GEN_46 : btb_pc_46; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_239 = fb_reg_redirect ? _GEN_47 : btb_pc_47; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_240 = fb_reg_redirect ? _GEN_48 : btb_pc_48; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_241 = fb_reg_redirect ? _GEN_49 : btb_pc_49; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_242 = fb_reg_redirect ? _GEN_50 : btb_pc_50; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_243 = fb_reg_redirect ? _GEN_51 : btb_pc_51; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_244 = fb_reg_redirect ? _GEN_52 : btb_pc_52; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_245 = fb_reg_redirect ? _GEN_53 : btb_pc_53; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_246 = fb_reg_redirect ? _GEN_54 : btb_pc_54; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_247 = fb_reg_redirect ? _GEN_55 : btb_pc_55; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_248 = fb_reg_redirect ? _GEN_56 : btb_pc_56; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_249 = fb_reg_redirect ? _GEN_57 : btb_pc_57; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_250 = fb_reg_redirect ? _GEN_58 : btb_pc_58; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_251 = fb_reg_redirect ? _GEN_59 : btb_pc_59; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_252 = fb_reg_redirect ? _GEN_60 : btb_pc_60; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_253 = fb_reg_redirect ? _GEN_61 : btb_pc_61; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_254 = fb_reg_redirect ? _GEN_62 : btb_pc_62; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_255 = fb_reg_redirect ? _GEN_63 : btb_pc_63; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_256 = fb_reg_redirect ? _GEN_64 : btb_target_0; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_257 = fb_reg_redirect ? _GEN_65 : btb_target_1; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_258 = fb_reg_redirect ? _GEN_66 : btb_target_2; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_259 = fb_reg_redirect ? _GEN_67 : btb_target_3; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_260 = fb_reg_redirect ? _GEN_68 : btb_target_4; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_261 = fb_reg_redirect ? _GEN_69 : btb_target_5; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_262 = fb_reg_redirect ? _GEN_70 : btb_target_6; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_263 = fb_reg_redirect ? _GEN_71 : btb_target_7; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_264 = fb_reg_redirect ? _GEN_72 : btb_target_8; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_265 = fb_reg_redirect ? _GEN_73 : btb_target_9; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_266 = fb_reg_redirect ? _GEN_74 : btb_target_10; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_267 = fb_reg_redirect ? _GEN_75 : btb_target_11; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_268 = fb_reg_redirect ? _GEN_76 : btb_target_12; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_269 = fb_reg_redirect ? _GEN_77 : btb_target_13; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_270 = fb_reg_redirect ? _GEN_78 : btb_target_14; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_271 = fb_reg_redirect ? _GEN_79 : btb_target_15; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_272 = fb_reg_redirect ? _GEN_80 : btb_target_16; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_273 = fb_reg_redirect ? _GEN_81 : btb_target_17; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_274 = fb_reg_redirect ? _GEN_82 : btb_target_18; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_275 = fb_reg_redirect ? _GEN_83 : btb_target_19; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_276 = fb_reg_redirect ? _GEN_84 : btb_target_20; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_277 = fb_reg_redirect ? _GEN_85 : btb_target_21; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_278 = fb_reg_redirect ? _GEN_86 : btb_target_22; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_279 = fb_reg_redirect ? _GEN_87 : btb_target_23; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_280 = fb_reg_redirect ? _GEN_88 : btb_target_24; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_281 = fb_reg_redirect ? _GEN_89 : btb_target_25; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_282 = fb_reg_redirect ? _GEN_90 : btb_target_26; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_283 = fb_reg_redirect ? _GEN_91 : btb_target_27; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_284 = fb_reg_redirect ? _GEN_92 : btb_target_28; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_285 = fb_reg_redirect ? _GEN_93 : btb_target_29; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_286 = fb_reg_redirect ? _GEN_94 : btb_target_30; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_287 = fb_reg_redirect ? _GEN_95 : btb_target_31; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_288 = fb_reg_redirect ? _GEN_96 : btb_target_32; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_289 = fb_reg_redirect ? _GEN_97 : btb_target_33; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_290 = fb_reg_redirect ? _GEN_98 : btb_target_34; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_291 = fb_reg_redirect ? _GEN_99 : btb_target_35; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_292 = fb_reg_redirect ? _GEN_100 : btb_target_36; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_293 = fb_reg_redirect ? _GEN_101 : btb_target_37; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_294 = fb_reg_redirect ? _GEN_102 : btb_target_38; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_295 = fb_reg_redirect ? _GEN_103 : btb_target_39; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_296 = fb_reg_redirect ? _GEN_104 : btb_target_40; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_297 = fb_reg_redirect ? _GEN_105 : btb_target_41; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_298 = fb_reg_redirect ? _GEN_106 : btb_target_42; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_299 = fb_reg_redirect ? _GEN_107 : btb_target_43; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_300 = fb_reg_redirect ? _GEN_108 : btb_target_44; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_301 = fb_reg_redirect ? _GEN_109 : btb_target_45; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_302 = fb_reg_redirect ? _GEN_110 : btb_target_46; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_303 = fb_reg_redirect ? _GEN_111 : btb_target_47; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_304 = fb_reg_redirect ? _GEN_112 : btb_target_48; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_305 = fb_reg_redirect ? _GEN_113 : btb_target_49; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_306 = fb_reg_redirect ? _GEN_114 : btb_target_50; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_307 = fb_reg_redirect ? _GEN_115 : btb_target_51; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_308 = fb_reg_redirect ? _GEN_116 : btb_target_52; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_309 = fb_reg_redirect ? _GEN_117 : btb_target_53; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_310 = fb_reg_redirect ? _GEN_118 : btb_target_54; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_311 = fb_reg_redirect ? _GEN_119 : btb_target_55; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_312 = fb_reg_redirect ? _GEN_120 : btb_target_56; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_313 = fb_reg_redirect ? _GEN_121 : btb_target_57; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_314 = fb_reg_redirect ? _GEN_122 : btb_target_58; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_315 = fb_reg_redirect ? _GEN_123 : btb_target_59; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_316 = fb_reg_redirect ? _GEN_124 : btb_target_60; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_317 = fb_reg_redirect ? _GEN_125 : btb_target_61; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_318 = fb_reg_redirect ? _GEN_126 : btb_target_62; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_319 = fb_reg_redirect ? _GEN_127 : btb_target_63; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_320 = fb_reg_redirect ? _GEN_128 : btb_btype_0; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_321 = fb_reg_redirect ? _GEN_129 : btb_btype_1; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_322 = fb_reg_redirect ? _GEN_130 : btb_btype_2; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_323 = fb_reg_redirect ? _GEN_131 : btb_btype_3; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_324 = fb_reg_redirect ? _GEN_132 : btb_btype_4; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_325 = fb_reg_redirect ? _GEN_133 : btb_btype_5; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_326 = fb_reg_redirect ? _GEN_134 : btb_btype_6; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_327 = fb_reg_redirect ? _GEN_135 : btb_btype_7; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_328 = fb_reg_redirect ? _GEN_136 : btb_btype_8; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_329 = fb_reg_redirect ? _GEN_137 : btb_btype_9; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_330 = fb_reg_redirect ? _GEN_138 : btb_btype_10; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_331 = fb_reg_redirect ? _GEN_139 : btb_btype_11; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_332 = fb_reg_redirect ? _GEN_140 : btb_btype_12; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_333 = fb_reg_redirect ? _GEN_141 : btb_btype_13; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_334 = fb_reg_redirect ? _GEN_142 : btb_btype_14; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_335 = fb_reg_redirect ? _GEN_143 : btb_btype_15; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_336 = fb_reg_redirect ? _GEN_144 : btb_btype_16; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_337 = fb_reg_redirect ? _GEN_145 : btb_btype_17; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_338 = fb_reg_redirect ? _GEN_146 : btb_btype_18; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_339 = fb_reg_redirect ? _GEN_147 : btb_btype_19; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_340 = fb_reg_redirect ? _GEN_148 : btb_btype_20; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_341 = fb_reg_redirect ? _GEN_149 : btb_btype_21; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_342 = fb_reg_redirect ? _GEN_150 : btb_btype_22; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_343 = fb_reg_redirect ? _GEN_151 : btb_btype_23; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_344 = fb_reg_redirect ? _GEN_152 : btb_btype_24; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_345 = fb_reg_redirect ? _GEN_153 : btb_btype_25; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_346 = fb_reg_redirect ? _GEN_154 : btb_btype_26; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_347 = fb_reg_redirect ? _GEN_155 : btb_btype_27; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_348 = fb_reg_redirect ? _GEN_156 : btb_btype_28; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_349 = fb_reg_redirect ? _GEN_157 : btb_btype_29; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_350 = fb_reg_redirect ? _GEN_158 : btb_btype_30; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_351 = fb_reg_redirect ? _GEN_159 : btb_btype_31; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_352 = fb_reg_redirect ? _GEN_160 : btb_btype_32; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_353 = fb_reg_redirect ? _GEN_161 : btb_btype_33; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_354 = fb_reg_redirect ? _GEN_162 : btb_btype_34; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_355 = fb_reg_redirect ? _GEN_163 : btb_btype_35; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_356 = fb_reg_redirect ? _GEN_164 : btb_btype_36; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_357 = fb_reg_redirect ? _GEN_165 : btb_btype_37; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_358 = fb_reg_redirect ? _GEN_166 : btb_btype_38; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_359 = fb_reg_redirect ? _GEN_167 : btb_btype_39; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_360 = fb_reg_redirect ? _GEN_168 : btb_btype_40; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_361 = fb_reg_redirect ? _GEN_169 : btb_btype_41; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_362 = fb_reg_redirect ? _GEN_170 : btb_btype_42; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_363 = fb_reg_redirect ? _GEN_171 : btb_btype_43; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_364 = fb_reg_redirect ? _GEN_172 : btb_btype_44; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_365 = fb_reg_redirect ? _GEN_173 : btb_btype_45; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_366 = fb_reg_redirect ? _GEN_174 : btb_btype_46; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_367 = fb_reg_redirect ? _GEN_175 : btb_btype_47; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_368 = fb_reg_redirect ? _GEN_176 : btb_btype_48; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_369 = fb_reg_redirect ? _GEN_177 : btb_btype_49; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_370 = fb_reg_redirect ? _GEN_178 : btb_btype_50; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_371 = fb_reg_redirect ? _GEN_179 : btb_btype_51; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_372 = fb_reg_redirect ? _GEN_180 : btb_btype_52; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_373 = fb_reg_redirect ? _GEN_181 : btb_btype_53; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_374 = fb_reg_redirect ? _GEN_182 : btb_btype_54; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_375 = fb_reg_redirect ? _GEN_183 : btb_btype_55; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_376 = fb_reg_redirect ? _GEN_184 : btb_btype_56; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_377 = fb_reg_redirect ? _GEN_185 : btb_btype_57; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_378 = fb_reg_redirect ? _GEN_186 : btb_btype_58; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_379 = fb_reg_redirect ? _GEN_187 : btb_btype_59; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_380 = fb_reg_redirect ? _GEN_188 : btb_btype_60; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_381 = fb_reg_redirect ? _GEN_189 : btb_btype_61; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_382 = fb_reg_redirect ? _GEN_190 : btb_btype_62; // @[BTB.scala 131:28:@4329.6]
  assign _GEN_383 = fb_reg_redirect ? _GEN_191 : btb_btype_63; // @[BTB.scala 131:28:@4329.6]
  assign _T_4159 = fb_reg_btype == 2'h2; // @[BTB.scala 136:24:@4334.6]
  assign _T_4163 = fb_wire_hcount != 2'h0; // @[BTB.scala 53:42:@4339.12]
  assign _T_4164 = fb_wire_hcount[1]; // @[BTB.scala 53:49:@4340.12]
  assign _T_4165 = fb_wire_hcount[0]; // @[BTB.scala 53:58:@4341.12]
  assign _T_4167 = _T_4165 == 1'h0; // @[BTB.scala 53:56:@4342.12]
  assign _T_4168 = _T_4164 | _T_4167; // @[BTB.scala 53:53:@4343.12]
  assign _T_4169 = {_T_4163,_T_4168}; // @[Cat.scala 30:58:@4344.12]
  assign _GEN_384 = 6'h0 == fb_wire_bindex ? _T_4169 : btb_hcount_0; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_385 = 6'h1 == fb_wire_bindex ? _T_4169 : btb_hcount_1; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_386 = 6'h2 == fb_wire_bindex ? _T_4169 : btb_hcount_2; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_387 = 6'h3 == fb_wire_bindex ? _T_4169 : btb_hcount_3; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_388 = 6'h4 == fb_wire_bindex ? _T_4169 : btb_hcount_4; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_389 = 6'h5 == fb_wire_bindex ? _T_4169 : btb_hcount_5; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_390 = 6'h6 == fb_wire_bindex ? _T_4169 : btb_hcount_6; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_391 = 6'h7 == fb_wire_bindex ? _T_4169 : btb_hcount_7; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_392 = 6'h8 == fb_wire_bindex ? _T_4169 : btb_hcount_8; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_393 = 6'h9 == fb_wire_bindex ? _T_4169 : btb_hcount_9; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_394 = 6'ha == fb_wire_bindex ? _T_4169 : btb_hcount_10; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_395 = 6'hb == fb_wire_bindex ? _T_4169 : btb_hcount_11; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_396 = 6'hc == fb_wire_bindex ? _T_4169 : btb_hcount_12; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_397 = 6'hd == fb_wire_bindex ? _T_4169 : btb_hcount_13; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_398 = 6'he == fb_wire_bindex ? _T_4169 : btb_hcount_14; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_399 = 6'hf == fb_wire_bindex ? _T_4169 : btb_hcount_15; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_400 = 6'h10 == fb_wire_bindex ? _T_4169 : btb_hcount_16; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_401 = 6'h11 == fb_wire_bindex ? _T_4169 : btb_hcount_17; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_402 = 6'h12 == fb_wire_bindex ? _T_4169 : btb_hcount_18; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_403 = 6'h13 == fb_wire_bindex ? _T_4169 : btb_hcount_19; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_404 = 6'h14 == fb_wire_bindex ? _T_4169 : btb_hcount_20; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_405 = 6'h15 == fb_wire_bindex ? _T_4169 : btb_hcount_21; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_406 = 6'h16 == fb_wire_bindex ? _T_4169 : btb_hcount_22; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_407 = 6'h17 == fb_wire_bindex ? _T_4169 : btb_hcount_23; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_408 = 6'h18 == fb_wire_bindex ? _T_4169 : btb_hcount_24; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_409 = 6'h19 == fb_wire_bindex ? _T_4169 : btb_hcount_25; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_410 = 6'h1a == fb_wire_bindex ? _T_4169 : btb_hcount_26; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_411 = 6'h1b == fb_wire_bindex ? _T_4169 : btb_hcount_27; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_412 = 6'h1c == fb_wire_bindex ? _T_4169 : btb_hcount_28; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_413 = 6'h1d == fb_wire_bindex ? _T_4169 : btb_hcount_29; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_414 = 6'h1e == fb_wire_bindex ? _T_4169 : btb_hcount_30; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_415 = 6'h1f == fb_wire_bindex ? _T_4169 : btb_hcount_31; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_416 = 6'h20 == fb_wire_bindex ? _T_4169 : btb_hcount_32; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_417 = 6'h21 == fb_wire_bindex ? _T_4169 : btb_hcount_33; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_418 = 6'h22 == fb_wire_bindex ? _T_4169 : btb_hcount_34; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_419 = 6'h23 == fb_wire_bindex ? _T_4169 : btb_hcount_35; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_420 = 6'h24 == fb_wire_bindex ? _T_4169 : btb_hcount_36; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_421 = 6'h25 == fb_wire_bindex ? _T_4169 : btb_hcount_37; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_422 = 6'h26 == fb_wire_bindex ? _T_4169 : btb_hcount_38; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_423 = 6'h27 == fb_wire_bindex ? _T_4169 : btb_hcount_39; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_424 = 6'h28 == fb_wire_bindex ? _T_4169 : btb_hcount_40; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_425 = 6'h29 == fb_wire_bindex ? _T_4169 : btb_hcount_41; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_426 = 6'h2a == fb_wire_bindex ? _T_4169 : btb_hcount_42; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_427 = 6'h2b == fb_wire_bindex ? _T_4169 : btb_hcount_43; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_428 = 6'h2c == fb_wire_bindex ? _T_4169 : btb_hcount_44; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_429 = 6'h2d == fb_wire_bindex ? _T_4169 : btb_hcount_45; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_430 = 6'h2e == fb_wire_bindex ? _T_4169 : btb_hcount_46; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_431 = 6'h2f == fb_wire_bindex ? _T_4169 : btb_hcount_47; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_432 = 6'h30 == fb_wire_bindex ? _T_4169 : btb_hcount_48; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_433 = 6'h31 == fb_wire_bindex ? _T_4169 : btb_hcount_49; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_434 = 6'h32 == fb_wire_bindex ? _T_4169 : btb_hcount_50; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_435 = 6'h33 == fb_wire_bindex ? _T_4169 : btb_hcount_51; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_436 = 6'h34 == fb_wire_bindex ? _T_4169 : btb_hcount_52; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_437 = 6'h35 == fb_wire_bindex ? _T_4169 : btb_hcount_53; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_438 = 6'h36 == fb_wire_bindex ? _T_4169 : btb_hcount_54; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_439 = 6'h37 == fb_wire_bindex ? _T_4169 : btb_hcount_55; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_440 = 6'h38 == fb_wire_bindex ? _T_4169 : btb_hcount_56; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_441 = 6'h39 == fb_wire_bindex ? _T_4169 : btb_hcount_57; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_442 = 6'h3a == fb_wire_bindex ? _T_4169 : btb_hcount_58; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_443 = 6'h3b == fb_wire_bindex ? _T_4169 : btb_hcount_59; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_444 = 6'h3c == fb_wire_bindex ? _T_4169 : btb_hcount_60; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_445 = 6'h3d == fb_wire_bindex ? _T_4169 : btb_hcount_61; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_446 = 6'h3e == fb_wire_bindex ? _T_4169 : btb_hcount_62; // @[BTB.scala 139:38:@4345.12]
  assign _GEN_447 = 6'h3f == fb_wire_bindex ? _T_4169 : btb_hcount_63; // @[BTB.scala 139:38:@4345.12]
  assign _T_4170 = ~ fb_wire_hcount; // @[BTB.scala 54:42:@4348.12]
  assign _T_4172 = _T_4170 == 2'h0; // @[BTB.scala 54:42:@4349.12]
  assign _T_4177 = _T_4164 & _T_4167; // @[BTB.scala 54:53:@4353.12]
  assign _T_4178 = {_T_4172,_T_4177}; // @[Cat.scala 30:58:@4354.12]
  assign _GEN_448 = 6'h0 == fb_wire_bindex ? _T_4178 : btb_hcount_0; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_449 = 6'h1 == fb_wire_bindex ? _T_4178 : btb_hcount_1; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_450 = 6'h2 == fb_wire_bindex ? _T_4178 : btb_hcount_2; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_451 = 6'h3 == fb_wire_bindex ? _T_4178 : btb_hcount_3; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_452 = 6'h4 == fb_wire_bindex ? _T_4178 : btb_hcount_4; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_453 = 6'h5 == fb_wire_bindex ? _T_4178 : btb_hcount_5; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_454 = 6'h6 == fb_wire_bindex ? _T_4178 : btb_hcount_6; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_455 = 6'h7 == fb_wire_bindex ? _T_4178 : btb_hcount_7; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_456 = 6'h8 == fb_wire_bindex ? _T_4178 : btb_hcount_8; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_457 = 6'h9 == fb_wire_bindex ? _T_4178 : btb_hcount_9; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_458 = 6'ha == fb_wire_bindex ? _T_4178 : btb_hcount_10; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_459 = 6'hb == fb_wire_bindex ? _T_4178 : btb_hcount_11; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_460 = 6'hc == fb_wire_bindex ? _T_4178 : btb_hcount_12; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_461 = 6'hd == fb_wire_bindex ? _T_4178 : btb_hcount_13; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_462 = 6'he == fb_wire_bindex ? _T_4178 : btb_hcount_14; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_463 = 6'hf == fb_wire_bindex ? _T_4178 : btb_hcount_15; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_464 = 6'h10 == fb_wire_bindex ? _T_4178 : btb_hcount_16; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_465 = 6'h11 == fb_wire_bindex ? _T_4178 : btb_hcount_17; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_466 = 6'h12 == fb_wire_bindex ? _T_4178 : btb_hcount_18; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_467 = 6'h13 == fb_wire_bindex ? _T_4178 : btb_hcount_19; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_468 = 6'h14 == fb_wire_bindex ? _T_4178 : btb_hcount_20; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_469 = 6'h15 == fb_wire_bindex ? _T_4178 : btb_hcount_21; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_470 = 6'h16 == fb_wire_bindex ? _T_4178 : btb_hcount_22; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_471 = 6'h17 == fb_wire_bindex ? _T_4178 : btb_hcount_23; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_472 = 6'h18 == fb_wire_bindex ? _T_4178 : btb_hcount_24; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_473 = 6'h19 == fb_wire_bindex ? _T_4178 : btb_hcount_25; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_474 = 6'h1a == fb_wire_bindex ? _T_4178 : btb_hcount_26; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_475 = 6'h1b == fb_wire_bindex ? _T_4178 : btb_hcount_27; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_476 = 6'h1c == fb_wire_bindex ? _T_4178 : btb_hcount_28; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_477 = 6'h1d == fb_wire_bindex ? _T_4178 : btb_hcount_29; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_478 = 6'h1e == fb_wire_bindex ? _T_4178 : btb_hcount_30; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_479 = 6'h1f == fb_wire_bindex ? _T_4178 : btb_hcount_31; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_480 = 6'h20 == fb_wire_bindex ? _T_4178 : btb_hcount_32; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_481 = 6'h21 == fb_wire_bindex ? _T_4178 : btb_hcount_33; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_482 = 6'h22 == fb_wire_bindex ? _T_4178 : btb_hcount_34; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_483 = 6'h23 == fb_wire_bindex ? _T_4178 : btb_hcount_35; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_484 = 6'h24 == fb_wire_bindex ? _T_4178 : btb_hcount_36; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_485 = 6'h25 == fb_wire_bindex ? _T_4178 : btb_hcount_37; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_486 = 6'h26 == fb_wire_bindex ? _T_4178 : btb_hcount_38; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_487 = 6'h27 == fb_wire_bindex ? _T_4178 : btb_hcount_39; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_488 = 6'h28 == fb_wire_bindex ? _T_4178 : btb_hcount_40; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_489 = 6'h29 == fb_wire_bindex ? _T_4178 : btb_hcount_41; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_490 = 6'h2a == fb_wire_bindex ? _T_4178 : btb_hcount_42; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_491 = 6'h2b == fb_wire_bindex ? _T_4178 : btb_hcount_43; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_492 = 6'h2c == fb_wire_bindex ? _T_4178 : btb_hcount_44; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_493 = 6'h2d == fb_wire_bindex ? _T_4178 : btb_hcount_45; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_494 = 6'h2e == fb_wire_bindex ? _T_4178 : btb_hcount_46; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_495 = 6'h2f == fb_wire_bindex ? _T_4178 : btb_hcount_47; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_496 = 6'h30 == fb_wire_bindex ? _T_4178 : btb_hcount_48; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_497 = 6'h31 == fb_wire_bindex ? _T_4178 : btb_hcount_49; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_498 = 6'h32 == fb_wire_bindex ? _T_4178 : btb_hcount_50; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_499 = 6'h33 == fb_wire_bindex ? _T_4178 : btb_hcount_51; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_500 = 6'h34 == fb_wire_bindex ? _T_4178 : btb_hcount_52; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_501 = 6'h35 == fb_wire_bindex ? _T_4178 : btb_hcount_53; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_502 = 6'h36 == fb_wire_bindex ? _T_4178 : btb_hcount_54; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_503 = 6'h37 == fb_wire_bindex ? _T_4178 : btb_hcount_55; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_504 = 6'h38 == fb_wire_bindex ? _T_4178 : btb_hcount_56; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_505 = 6'h39 == fb_wire_bindex ? _T_4178 : btb_hcount_57; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_506 = 6'h3a == fb_wire_bindex ? _T_4178 : btb_hcount_58; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_507 = 6'h3b == fb_wire_bindex ? _T_4178 : btb_hcount_59; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_508 = 6'h3c == fb_wire_bindex ? _T_4178 : btb_hcount_60; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_509 = 6'h3d == fb_wire_bindex ? _T_4178 : btb_hcount_61; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_510 = 6'h3e == fb_wire_bindex ? _T_4178 : btb_hcount_62; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_511 = 6'h3f == fb_wire_bindex ? _T_4178 : btb_hcount_63; // @[BTB.scala 141:38:@4355.12]
  assign _GEN_512 = fb_reg_redirect ? _GEN_384 : _GEN_448; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_513 = fb_reg_redirect ? _GEN_385 : _GEN_449; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_514 = fb_reg_redirect ? _GEN_386 : _GEN_450; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_515 = fb_reg_redirect ? _GEN_387 : _GEN_451; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_516 = fb_reg_redirect ? _GEN_388 : _GEN_452; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_517 = fb_reg_redirect ? _GEN_389 : _GEN_453; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_518 = fb_reg_redirect ? _GEN_390 : _GEN_454; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_519 = fb_reg_redirect ? _GEN_391 : _GEN_455; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_520 = fb_reg_redirect ? _GEN_392 : _GEN_456; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_521 = fb_reg_redirect ? _GEN_393 : _GEN_457; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_522 = fb_reg_redirect ? _GEN_394 : _GEN_458; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_523 = fb_reg_redirect ? _GEN_395 : _GEN_459; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_524 = fb_reg_redirect ? _GEN_396 : _GEN_460; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_525 = fb_reg_redirect ? _GEN_397 : _GEN_461; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_526 = fb_reg_redirect ? _GEN_398 : _GEN_462; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_527 = fb_reg_redirect ? _GEN_399 : _GEN_463; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_528 = fb_reg_redirect ? _GEN_400 : _GEN_464; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_529 = fb_reg_redirect ? _GEN_401 : _GEN_465; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_530 = fb_reg_redirect ? _GEN_402 : _GEN_466; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_531 = fb_reg_redirect ? _GEN_403 : _GEN_467; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_532 = fb_reg_redirect ? _GEN_404 : _GEN_468; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_533 = fb_reg_redirect ? _GEN_405 : _GEN_469; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_534 = fb_reg_redirect ? _GEN_406 : _GEN_470; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_535 = fb_reg_redirect ? _GEN_407 : _GEN_471; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_536 = fb_reg_redirect ? _GEN_408 : _GEN_472; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_537 = fb_reg_redirect ? _GEN_409 : _GEN_473; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_538 = fb_reg_redirect ? _GEN_410 : _GEN_474; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_539 = fb_reg_redirect ? _GEN_411 : _GEN_475; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_540 = fb_reg_redirect ? _GEN_412 : _GEN_476; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_541 = fb_reg_redirect ? _GEN_413 : _GEN_477; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_542 = fb_reg_redirect ? _GEN_414 : _GEN_478; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_543 = fb_reg_redirect ? _GEN_415 : _GEN_479; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_544 = fb_reg_redirect ? _GEN_416 : _GEN_480; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_545 = fb_reg_redirect ? _GEN_417 : _GEN_481; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_546 = fb_reg_redirect ? _GEN_418 : _GEN_482; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_547 = fb_reg_redirect ? _GEN_419 : _GEN_483; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_548 = fb_reg_redirect ? _GEN_420 : _GEN_484; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_549 = fb_reg_redirect ? _GEN_421 : _GEN_485; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_550 = fb_reg_redirect ? _GEN_422 : _GEN_486; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_551 = fb_reg_redirect ? _GEN_423 : _GEN_487; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_552 = fb_reg_redirect ? _GEN_424 : _GEN_488; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_553 = fb_reg_redirect ? _GEN_425 : _GEN_489; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_554 = fb_reg_redirect ? _GEN_426 : _GEN_490; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_555 = fb_reg_redirect ? _GEN_427 : _GEN_491; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_556 = fb_reg_redirect ? _GEN_428 : _GEN_492; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_557 = fb_reg_redirect ? _GEN_429 : _GEN_493; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_558 = fb_reg_redirect ? _GEN_430 : _GEN_494; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_559 = fb_reg_redirect ? _GEN_431 : _GEN_495; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_560 = fb_reg_redirect ? _GEN_432 : _GEN_496; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_561 = fb_reg_redirect ? _GEN_433 : _GEN_497; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_562 = fb_reg_redirect ? _GEN_434 : _GEN_498; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_563 = fb_reg_redirect ? _GEN_435 : _GEN_499; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_564 = fb_reg_redirect ? _GEN_436 : _GEN_500; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_565 = fb_reg_redirect ? _GEN_437 : _GEN_501; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_566 = fb_reg_redirect ? _GEN_438 : _GEN_502; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_567 = fb_reg_redirect ? _GEN_439 : _GEN_503; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_568 = fb_reg_redirect ? _GEN_440 : _GEN_504; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_569 = fb_reg_redirect ? _GEN_441 : _GEN_505; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_570 = fb_reg_redirect ? _GEN_442 : _GEN_506; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_571 = fb_reg_redirect ? _GEN_443 : _GEN_507; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_572 = fb_reg_redirect ? _GEN_444 : _GEN_508; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_573 = fb_reg_redirect ? _GEN_445 : _GEN_509; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_574 = fb_reg_redirect ? _GEN_446 : _GEN_510; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_575 = fb_reg_redirect ? _GEN_447 : _GEN_511; // @[BTB.scala 138:32:@4338.10]
  assign _GEN_576 = 6'h0 == fb_wire_bindex ? 2'h2 : btb_hcount_0; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_577 = 6'h1 == fb_wire_bindex ? 2'h2 : btb_hcount_1; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_578 = 6'h2 == fb_wire_bindex ? 2'h2 : btb_hcount_2; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_579 = 6'h3 == fb_wire_bindex ? 2'h2 : btb_hcount_3; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_580 = 6'h4 == fb_wire_bindex ? 2'h2 : btb_hcount_4; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_581 = 6'h5 == fb_wire_bindex ? 2'h2 : btb_hcount_5; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_582 = 6'h6 == fb_wire_bindex ? 2'h2 : btb_hcount_6; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_583 = 6'h7 == fb_wire_bindex ? 2'h2 : btb_hcount_7; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_584 = 6'h8 == fb_wire_bindex ? 2'h2 : btb_hcount_8; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_585 = 6'h9 == fb_wire_bindex ? 2'h2 : btb_hcount_9; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_586 = 6'ha == fb_wire_bindex ? 2'h2 : btb_hcount_10; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_587 = 6'hb == fb_wire_bindex ? 2'h2 : btb_hcount_11; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_588 = 6'hc == fb_wire_bindex ? 2'h2 : btb_hcount_12; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_589 = 6'hd == fb_wire_bindex ? 2'h2 : btb_hcount_13; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_590 = 6'he == fb_wire_bindex ? 2'h2 : btb_hcount_14; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_591 = 6'hf == fb_wire_bindex ? 2'h2 : btb_hcount_15; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_592 = 6'h10 == fb_wire_bindex ? 2'h2 : btb_hcount_16; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_593 = 6'h11 == fb_wire_bindex ? 2'h2 : btb_hcount_17; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_594 = 6'h12 == fb_wire_bindex ? 2'h2 : btb_hcount_18; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_595 = 6'h13 == fb_wire_bindex ? 2'h2 : btb_hcount_19; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_596 = 6'h14 == fb_wire_bindex ? 2'h2 : btb_hcount_20; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_597 = 6'h15 == fb_wire_bindex ? 2'h2 : btb_hcount_21; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_598 = 6'h16 == fb_wire_bindex ? 2'h2 : btb_hcount_22; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_599 = 6'h17 == fb_wire_bindex ? 2'h2 : btb_hcount_23; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_600 = 6'h18 == fb_wire_bindex ? 2'h2 : btb_hcount_24; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_601 = 6'h19 == fb_wire_bindex ? 2'h2 : btb_hcount_25; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_602 = 6'h1a == fb_wire_bindex ? 2'h2 : btb_hcount_26; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_603 = 6'h1b == fb_wire_bindex ? 2'h2 : btb_hcount_27; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_604 = 6'h1c == fb_wire_bindex ? 2'h2 : btb_hcount_28; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_605 = 6'h1d == fb_wire_bindex ? 2'h2 : btb_hcount_29; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_606 = 6'h1e == fb_wire_bindex ? 2'h2 : btb_hcount_30; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_607 = 6'h1f == fb_wire_bindex ? 2'h2 : btb_hcount_31; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_608 = 6'h20 == fb_wire_bindex ? 2'h2 : btb_hcount_32; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_609 = 6'h21 == fb_wire_bindex ? 2'h2 : btb_hcount_33; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_610 = 6'h22 == fb_wire_bindex ? 2'h2 : btb_hcount_34; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_611 = 6'h23 == fb_wire_bindex ? 2'h2 : btb_hcount_35; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_612 = 6'h24 == fb_wire_bindex ? 2'h2 : btb_hcount_36; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_613 = 6'h25 == fb_wire_bindex ? 2'h2 : btb_hcount_37; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_614 = 6'h26 == fb_wire_bindex ? 2'h2 : btb_hcount_38; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_615 = 6'h27 == fb_wire_bindex ? 2'h2 : btb_hcount_39; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_616 = 6'h28 == fb_wire_bindex ? 2'h2 : btb_hcount_40; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_617 = 6'h29 == fb_wire_bindex ? 2'h2 : btb_hcount_41; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_618 = 6'h2a == fb_wire_bindex ? 2'h2 : btb_hcount_42; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_619 = 6'h2b == fb_wire_bindex ? 2'h2 : btb_hcount_43; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_620 = 6'h2c == fb_wire_bindex ? 2'h2 : btb_hcount_44; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_621 = 6'h2d == fb_wire_bindex ? 2'h2 : btb_hcount_45; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_622 = 6'h2e == fb_wire_bindex ? 2'h2 : btb_hcount_46; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_623 = 6'h2f == fb_wire_bindex ? 2'h2 : btb_hcount_47; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_624 = 6'h30 == fb_wire_bindex ? 2'h2 : btb_hcount_48; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_625 = 6'h31 == fb_wire_bindex ? 2'h2 : btb_hcount_49; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_626 = 6'h32 == fb_wire_bindex ? 2'h2 : btb_hcount_50; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_627 = 6'h33 == fb_wire_bindex ? 2'h2 : btb_hcount_51; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_628 = 6'h34 == fb_wire_bindex ? 2'h2 : btb_hcount_52; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_629 = 6'h35 == fb_wire_bindex ? 2'h2 : btb_hcount_53; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_630 = 6'h36 == fb_wire_bindex ? 2'h2 : btb_hcount_54; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_631 = 6'h37 == fb_wire_bindex ? 2'h2 : btb_hcount_55; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_632 = 6'h38 == fb_wire_bindex ? 2'h2 : btb_hcount_56; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_633 = 6'h39 == fb_wire_bindex ? 2'h2 : btb_hcount_57; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_634 = 6'h3a == fb_wire_bindex ? 2'h2 : btb_hcount_58; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_635 = 6'h3b == fb_wire_bindex ? 2'h2 : btb_hcount_59; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_636 = 6'h3c == fb_wire_bindex ? 2'h2 : btb_hcount_60; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_637 = 6'h3d == fb_wire_bindex ? 2'h2 : btb_hcount_61; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_638 = 6'h3e == fb_wire_bindex ? 2'h2 : btb_hcount_62; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_639 = 6'h3f == fb_wire_bindex ? 2'h2 : btb_hcount_63; // @[BTB.scala 144:36:@4360.12]
  assign _GEN_640 = fb_reg_redirect ? _GEN_576 : btb_hcount_0; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_641 = fb_reg_redirect ? _GEN_577 : btb_hcount_1; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_642 = fb_reg_redirect ? _GEN_578 : btb_hcount_2; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_643 = fb_reg_redirect ? _GEN_579 : btb_hcount_3; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_644 = fb_reg_redirect ? _GEN_580 : btb_hcount_4; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_645 = fb_reg_redirect ? _GEN_581 : btb_hcount_5; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_646 = fb_reg_redirect ? _GEN_582 : btb_hcount_6; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_647 = fb_reg_redirect ? _GEN_583 : btb_hcount_7; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_648 = fb_reg_redirect ? _GEN_584 : btb_hcount_8; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_649 = fb_reg_redirect ? _GEN_585 : btb_hcount_9; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_650 = fb_reg_redirect ? _GEN_586 : btb_hcount_10; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_651 = fb_reg_redirect ? _GEN_587 : btb_hcount_11; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_652 = fb_reg_redirect ? _GEN_588 : btb_hcount_12; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_653 = fb_reg_redirect ? _GEN_589 : btb_hcount_13; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_654 = fb_reg_redirect ? _GEN_590 : btb_hcount_14; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_655 = fb_reg_redirect ? _GEN_591 : btb_hcount_15; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_656 = fb_reg_redirect ? _GEN_592 : btb_hcount_16; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_657 = fb_reg_redirect ? _GEN_593 : btb_hcount_17; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_658 = fb_reg_redirect ? _GEN_594 : btb_hcount_18; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_659 = fb_reg_redirect ? _GEN_595 : btb_hcount_19; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_660 = fb_reg_redirect ? _GEN_596 : btb_hcount_20; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_661 = fb_reg_redirect ? _GEN_597 : btb_hcount_21; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_662 = fb_reg_redirect ? _GEN_598 : btb_hcount_22; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_663 = fb_reg_redirect ? _GEN_599 : btb_hcount_23; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_664 = fb_reg_redirect ? _GEN_600 : btb_hcount_24; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_665 = fb_reg_redirect ? _GEN_601 : btb_hcount_25; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_666 = fb_reg_redirect ? _GEN_602 : btb_hcount_26; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_667 = fb_reg_redirect ? _GEN_603 : btb_hcount_27; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_668 = fb_reg_redirect ? _GEN_604 : btb_hcount_28; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_669 = fb_reg_redirect ? _GEN_605 : btb_hcount_29; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_670 = fb_reg_redirect ? _GEN_606 : btb_hcount_30; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_671 = fb_reg_redirect ? _GEN_607 : btb_hcount_31; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_672 = fb_reg_redirect ? _GEN_608 : btb_hcount_32; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_673 = fb_reg_redirect ? _GEN_609 : btb_hcount_33; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_674 = fb_reg_redirect ? _GEN_610 : btb_hcount_34; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_675 = fb_reg_redirect ? _GEN_611 : btb_hcount_35; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_676 = fb_reg_redirect ? _GEN_612 : btb_hcount_36; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_677 = fb_reg_redirect ? _GEN_613 : btb_hcount_37; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_678 = fb_reg_redirect ? _GEN_614 : btb_hcount_38; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_679 = fb_reg_redirect ? _GEN_615 : btb_hcount_39; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_680 = fb_reg_redirect ? _GEN_616 : btb_hcount_40; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_681 = fb_reg_redirect ? _GEN_617 : btb_hcount_41; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_682 = fb_reg_redirect ? _GEN_618 : btb_hcount_42; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_683 = fb_reg_redirect ? _GEN_619 : btb_hcount_43; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_684 = fb_reg_redirect ? _GEN_620 : btb_hcount_44; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_685 = fb_reg_redirect ? _GEN_621 : btb_hcount_45; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_686 = fb_reg_redirect ? _GEN_622 : btb_hcount_46; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_687 = fb_reg_redirect ? _GEN_623 : btb_hcount_47; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_688 = fb_reg_redirect ? _GEN_624 : btb_hcount_48; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_689 = fb_reg_redirect ? _GEN_625 : btb_hcount_49; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_690 = fb_reg_redirect ? _GEN_626 : btb_hcount_50; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_691 = fb_reg_redirect ? _GEN_627 : btb_hcount_51; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_692 = fb_reg_redirect ? _GEN_628 : btb_hcount_52; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_693 = fb_reg_redirect ? _GEN_629 : btb_hcount_53; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_694 = fb_reg_redirect ? _GEN_630 : btb_hcount_54; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_695 = fb_reg_redirect ? _GEN_631 : btb_hcount_55; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_696 = fb_reg_redirect ? _GEN_632 : btb_hcount_56; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_697 = fb_reg_redirect ? _GEN_633 : btb_hcount_57; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_698 = fb_reg_redirect ? _GEN_634 : btb_hcount_58; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_699 = fb_reg_redirect ? _GEN_635 : btb_hcount_59; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_700 = fb_reg_redirect ? _GEN_636 : btb_hcount_60; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_701 = fb_reg_redirect ? _GEN_637 : btb_hcount_61; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_702 = fb_reg_redirect ? _GEN_638 : btb_hcount_62; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_703 = fb_reg_redirect ? _GEN_639 : btb_hcount_63; // @[BTB.scala 143:35:@4359.10]
  assign _GEN_704 = _T_3407 ? _GEN_512 : _GEN_640; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_705 = _T_3407 ? _GEN_513 : _GEN_641; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_706 = _T_3407 ? _GEN_514 : _GEN_642; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_707 = _T_3407 ? _GEN_515 : _GEN_643; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_708 = _T_3407 ? _GEN_516 : _GEN_644; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_709 = _T_3407 ? _GEN_517 : _GEN_645; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_710 = _T_3407 ? _GEN_518 : _GEN_646; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_711 = _T_3407 ? _GEN_519 : _GEN_647; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_712 = _T_3407 ? _GEN_520 : _GEN_648; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_713 = _T_3407 ? _GEN_521 : _GEN_649; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_714 = _T_3407 ? _GEN_522 : _GEN_650; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_715 = _T_3407 ? _GEN_523 : _GEN_651; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_716 = _T_3407 ? _GEN_524 : _GEN_652; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_717 = _T_3407 ? _GEN_525 : _GEN_653; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_718 = _T_3407 ? _GEN_526 : _GEN_654; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_719 = _T_3407 ? _GEN_527 : _GEN_655; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_720 = _T_3407 ? _GEN_528 : _GEN_656; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_721 = _T_3407 ? _GEN_529 : _GEN_657; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_722 = _T_3407 ? _GEN_530 : _GEN_658; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_723 = _T_3407 ? _GEN_531 : _GEN_659; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_724 = _T_3407 ? _GEN_532 : _GEN_660; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_725 = _T_3407 ? _GEN_533 : _GEN_661; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_726 = _T_3407 ? _GEN_534 : _GEN_662; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_727 = _T_3407 ? _GEN_535 : _GEN_663; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_728 = _T_3407 ? _GEN_536 : _GEN_664; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_729 = _T_3407 ? _GEN_537 : _GEN_665; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_730 = _T_3407 ? _GEN_538 : _GEN_666; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_731 = _T_3407 ? _GEN_539 : _GEN_667; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_732 = _T_3407 ? _GEN_540 : _GEN_668; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_733 = _T_3407 ? _GEN_541 : _GEN_669; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_734 = _T_3407 ? _GEN_542 : _GEN_670; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_735 = _T_3407 ? _GEN_543 : _GEN_671; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_736 = _T_3407 ? _GEN_544 : _GEN_672; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_737 = _T_3407 ? _GEN_545 : _GEN_673; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_738 = _T_3407 ? _GEN_546 : _GEN_674; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_739 = _T_3407 ? _GEN_547 : _GEN_675; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_740 = _T_3407 ? _GEN_548 : _GEN_676; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_741 = _T_3407 ? _GEN_549 : _GEN_677; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_742 = _T_3407 ? _GEN_550 : _GEN_678; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_743 = _T_3407 ? _GEN_551 : _GEN_679; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_744 = _T_3407 ? _GEN_552 : _GEN_680; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_745 = _T_3407 ? _GEN_553 : _GEN_681; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_746 = _T_3407 ? _GEN_554 : _GEN_682; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_747 = _T_3407 ? _GEN_555 : _GEN_683; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_748 = _T_3407 ? _GEN_556 : _GEN_684; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_749 = _T_3407 ? _GEN_557 : _GEN_685; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_750 = _T_3407 ? _GEN_558 : _GEN_686; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_751 = _T_3407 ? _GEN_559 : _GEN_687; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_752 = _T_3407 ? _GEN_560 : _GEN_688; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_753 = _T_3407 ? _GEN_561 : _GEN_689; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_754 = _T_3407 ? _GEN_562 : _GEN_690; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_755 = _T_3407 ? _GEN_563 : _GEN_691; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_756 = _T_3407 ? _GEN_564 : _GEN_692; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_757 = _T_3407 ? _GEN_565 : _GEN_693; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_758 = _T_3407 ? _GEN_566 : _GEN_694; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_759 = _T_3407 ? _GEN_567 : _GEN_695; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_760 = _T_3407 ? _GEN_568 : _GEN_696; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_761 = _T_3407 ? _GEN_569 : _GEN_697; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_762 = _T_3407 ? _GEN_570 : _GEN_698; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_763 = _T_3407 ? _GEN_571 : _GEN_699; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_764 = _T_3407 ? _GEN_572 : _GEN_700; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_765 = _T_3407 ? _GEN_573 : _GEN_701; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_766 = _T_3407 ? _GEN_574 : _GEN_702; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_767 = _T_3407 ? _GEN_575 : _GEN_703; // @[BTB.scala 137:28:@4337.8]
  assign _GEN_768 = _T_4159 ? _GEN_704 : btb_hcount_0; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_769 = _T_4159 ? _GEN_705 : btb_hcount_1; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_770 = _T_4159 ? _GEN_706 : btb_hcount_2; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_771 = _T_4159 ? _GEN_707 : btb_hcount_3; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_772 = _T_4159 ? _GEN_708 : btb_hcount_4; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_773 = _T_4159 ? _GEN_709 : btb_hcount_5; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_774 = _T_4159 ? _GEN_710 : btb_hcount_6; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_775 = _T_4159 ? _GEN_711 : btb_hcount_7; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_776 = _T_4159 ? _GEN_712 : btb_hcount_8; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_777 = _T_4159 ? _GEN_713 : btb_hcount_9; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_778 = _T_4159 ? _GEN_714 : btb_hcount_10; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_779 = _T_4159 ? _GEN_715 : btb_hcount_11; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_780 = _T_4159 ? _GEN_716 : btb_hcount_12; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_781 = _T_4159 ? _GEN_717 : btb_hcount_13; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_782 = _T_4159 ? _GEN_718 : btb_hcount_14; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_783 = _T_4159 ? _GEN_719 : btb_hcount_15; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_784 = _T_4159 ? _GEN_720 : btb_hcount_16; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_785 = _T_4159 ? _GEN_721 : btb_hcount_17; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_786 = _T_4159 ? _GEN_722 : btb_hcount_18; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_787 = _T_4159 ? _GEN_723 : btb_hcount_19; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_788 = _T_4159 ? _GEN_724 : btb_hcount_20; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_789 = _T_4159 ? _GEN_725 : btb_hcount_21; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_790 = _T_4159 ? _GEN_726 : btb_hcount_22; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_791 = _T_4159 ? _GEN_727 : btb_hcount_23; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_792 = _T_4159 ? _GEN_728 : btb_hcount_24; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_793 = _T_4159 ? _GEN_729 : btb_hcount_25; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_794 = _T_4159 ? _GEN_730 : btb_hcount_26; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_795 = _T_4159 ? _GEN_731 : btb_hcount_27; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_796 = _T_4159 ? _GEN_732 : btb_hcount_28; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_797 = _T_4159 ? _GEN_733 : btb_hcount_29; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_798 = _T_4159 ? _GEN_734 : btb_hcount_30; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_799 = _T_4159 ? _GEN_735 : btb_hcount_31; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_800 = _T_4159 ? _GEN_736 : btb_hcount_32; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_801 = _T_4159 ? _GEN_737 : btb_hcount_33; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_802 = _T_4159 ? _GEN_738 : btb_hcount_34; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_803 = _T_4159 ? _GEN_739 : btb_hcount_35; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_804 = _T_4159 ? _GEN_740 : btb_hcount_36; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_805 = _T_4159 ? _GEN_741 : btb_hcount_37; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_806 = _T_4159 ? _GEN_742 : btb_hcount_38; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_807 = _T_4159 ? _GEN_743 : btb_hcount_39; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_808 = _T_4159 ? _GEN_744 : btb_hcount_40; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_809 = _T_4159 ? _GEN_745 : btb_hcount_41; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_810 = _T_4159 ? _GEN_746 : btb_hcount_42; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_811 = _T_4159 ? _GEN_747 : btb_hcount_43; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_812 = _T_4159 ? _GEN_748 : btb_hcount_44; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_813 = _T_4159 ? _GEN_749 : btb_hcount_45; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_814 = _T_4159 ? _GEN_750 : btb_hcount_46; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_815 = _T_4159 ? _GEN_751 : btb_hcount_47; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_816 = _T_4159 ? _GEN_752 : btb_hcount_48; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_817 = _T_4159 ? _GEN_753 : btb_hcount_49; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_818 = _T_4159 ? _GEN_754 : btb_hcount_50; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_819 = _T_4159 ? _GEN_755 : btb_hcount_51; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_820 = _T_4159 ? _GEN_756 : btb_hcount_52; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_821 = _T_4159 ? _GEN_757 : btb_hcount_53; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_822 = _T_4159 ? _GEN_758 : btb_hcount_54; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_823 = _T_4159 ? _GEN_759 : btb_hcount_55; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_824 = _T_4159 ? _GEN_760 : btb_hcount_56; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_825 = _T_4159 ? _GEN_761 : btb_hcount_57; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_826 = _T_4159 ? _GEN_762 : btb_hcount_58; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_827 = _T_4159 ? _GEN_763 : btb_hcount_59; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_828 = _T_4159 ? _GEN_764 : btb_hcount_60; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_829 = _T_4159 ? _GEN_765 : btb_hcount_61; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_830 = _T_4159 ? _GEN_766 : btb_hcount_62; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_831 = _T_4159 ? _GEN_767 : btb_hcount_63; // @[BTB.scala 136:46:@4335.6]
  assign _GEN_832 = fb_reg_valid ? _GEN_192 : btb_pc_0; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_833 = fb_reg_valid ? _GEN_193 : btb_pc_1; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_834 = fb_reg_valid ? _GEN_194 : btb_pc_2; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_835 = fb_reg_valid ? _GEN_195 : btb_pc_3; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_836 = fb_reg_valid ? _GEN_196 : btb_pc_4; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_837 = fb_reg_valid ? _GEN_197 : btb_pc_5; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_838 = fb_reg_valid ? _GEN_198 : btb_pc_6; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_839 = fb_reg_valid ? _GEN_199 : btb_pc_7; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_840 = fb_reg_valid ? _GEN_200 : btb_pc_8; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_841 = fb_reg_valid ? _GEN_201 : btb_pc_9; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_842 = fb_reg_valid ? _GEN_202 : btb_pc_10; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_843 = fb_reg_valid ? _GEN_203 : btb_pc_11; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_844 = fb_reg_valid ? _GEN_204 : btb_pc_12; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_845 = fb_reg_valid ? _GEN_205 : btb_pc_13; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_846 = fb_reg_valid ? _GEN_206 : btb_pc_14; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_847 = fb_reg_valid ? _GEN_207 : btb_pc_15; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_848 = fb_reg_valid ? _GEN_208 : btb_pc_16; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_849 = fb_reg_valid ? _GEN_209 : btb_pc_17; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_850 = fb_reg_valid ? _GEN_210 : btb_pc_18; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_851 = fb_reg_valid ? _GEN_211 : btb_pc_19; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_852 = fb_reg_valid ? _GEN_212 : btb_pc_20; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_853 = fb_reg_valid ? _GEN_213 : btb_pc_21; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_854 = fb_reg_valid ? _GEN_214 : btb_pc_22; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_855 = fb_reg_valid ? _GEN_215 : btb_pc_23; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_856 = fb_reg_valid ? _GEN_216 : btb_pc_24; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_857 = fb_reg_valid ? _GEN_217 : btb_pc_25; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_858 = fb_reg_valid ? _GEN_218 : btb_pc_26; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_859 = fb_reg_valid ? _GEN_219 : btb_pc_27; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_860 = fb_reg_valid ? _GEN_220 : btb_pc_28; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_861 = fb_reg_valid ? _GEN_221 : btb_pc_29; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_862 = fb_reg_valid ? _GEN_222 : btb_pc_30; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_863 = fb_reg_valid ? _GEN_223 : btb_pc_31; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_864 = fb_reg_valid ? _GEN_224 : btb_pc_32; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_865 = fb_reg_valid ? _GEN_225 : btb_pc_33; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_866 = fb_reg_valid ? _GEN_226 : btb_pc_34; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_867 = fb_reg_valid ? _GEN_227 : btb_pc_35; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_868 = fb_reg_valid ? _GEN_228 : btb_pc_36; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_869 = fb_reg_valid ? _GEN_229 : btb_pc_37; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_870 = fb_reg_valid ? _GEN_230 : btb_pc_38; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_871 = fb_reg_valid ? _GEN_231 : btb_pc_39; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_872 = fb_reg_valid ? _GEN_232 : btb_pc_40; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_873 = fb_reg_valid ? _GEN_233 : btb_pc_41; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_874 = fb_reg_valid ? _GEN_234 : btb_pc_42; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_875 = fb_reg_valid ? _GEN_235 : btb_pc_43; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_876 = fb_reg_valid ? _GEN_236 : btb_pc_44; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_877 = fb_reg_valid ? _GEN_237 : btb_pc_45; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_878 = fb_reg_valid ? _GEN_238 : btb_pc_46; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_879 = fb_reg_valid ? _GEN_239 : btb_pc_47; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_880 = fb_reg_valid ? _GEN_240 : btb_pc_48; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_881 = fb_reg_valid ? _GEN_241 : btb_pc_49; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_882 = fb_reg_valid ? _GEN_242 : btb_pc_50; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_883 = fb_reg_valid ? _GEN_243 : btb_pc_51; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_884 = fb_reg_valid ? _GEN_244 : btb_pc_52; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_885 = fb_reg_valid ? _GEN_245 : btb_pc_53; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_886 = fb_reg_valid ? _GEN_246 : btb_pc_54; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_887 = fb_reg_valid ? _GEN_247 : btb_pc_55; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_888 = fb_reg_valid ? _GEN_248 : btb_pc_56; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_889 = fb_reg_valid ? _GEN_249 : btb_pc_57; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_890 = fb_reg_valid ? _GEN_250 : btb_pc_58; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_891 = fb_reg_valid ? _GEN_251 : btb_pc_59; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_892 = fb_reg_valid ? _GEN_252 : btb_pc_60; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_893 = fb_reg_valid ? _GEN_253 : btb_pc_61; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_894 = fb_reg_valid ? _GEN_254 : btb_pc_62; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_895 = fb_reg_valid ? _GEN_255 : btb_pc_63; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_896 = fb_reg_valid ? _GEN_256 : btb_target_0; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_897 = fb_reg_valid ? _GEN_257 : btb_target_1; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_898 = fb_reg_valid ? _GEN_258 : btb_target_2; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_899 = fb_reg_valid ? _GEN_259 : btb_target_3; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_900 = fb_reg_valid ? _GEN_260 : btb_target_4; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_901 = fb_reg_valid ? _GEN_261 : btb_target_5; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_902 = fb_reg_valid ? _GEN_262 : btb_target_6; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_903 = fb_reg_valid ? _GEN_263 : btb_target_7; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_904 = fb_reg_valid ? _GEN_264 : btb_target_8; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_905 = fb_reg_valid ? _GEN_265 : btb_target_9; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_906 = fb_reg_valid ? _GEN_266 : btb_target_10; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_907 = fb_reg_valid ? _GEN_267 : btb_target_11; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_908 = fb_reg_valid ? _GEN_268 : btb_target_12; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_909 = fb_reg_valid ? _GEN_269 : btb_target_13; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_910 = fb_reg_valid ? _GEN_270 : btb_target_14; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_911 = fb_reg_valid ? _GEN_271 : btb_target_15; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_912 = fb_reg_valid ? _GEN_272 : btb_target_16; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_913 = fb_reg_valid ? _GEN_273 : btb_target_17; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_914 = fb_reg_valid ? _GEN_274 : btb_target_18; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_915 = fb_reg_valid ? _GEN_275 : btb_target_19; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_916 = fb_reg_valid ? _GEN_276 : btb_target_20; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_917 = fb_reg_valid ? _GEN_277 : btb_target_21; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_918 = fb_reg_valid ? _GEN_278 : btb_target_22; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_919 = fb_reg_valid ? _GEN_279 : btb_target_23; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_920 = fb_reg_valid ? _GEN_280 : btb_target_24; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_921 = fb_reg_valid ? _GEN_281 : btb_target_25; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_922 = fb_reg_valid ? _GEN_282 : btb_target_26; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_923 = fb_reg_valid ? _GEN_283 : btb_target_27; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_924 = fb_reg_valid ? _GEN_284 : btb_target_28; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_925 = fb_reg_valid ? _GEN_285 : btb_target_29; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_926 = fb_reg_valid ? _GEN_286 : btb_target_30; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_927 = fb_reg_valid ? _GEN_287 : btb_target_31; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_928 = fb_reg_valid ? _GEN_288 : btb_target_32; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_929 = fb_reg_valid ? _GEN_289 : btb_target_33; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_930 = fb_reg_valid ? _GEN_290 : btb_target_34; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_931 = fb_reg_valid ? _GEN_291 : btb_target_35; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_932 = fb_reg_valid ? _GEN_292 : btb_target_36; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_933 = fb_reg_valid ? _GEN_293 : btb_target_37; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_934 = fb_reg_valid ? _GEN_294 : btb_target_38; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_935 = fb_reg_valid ? _GEN_295 : btb_target_39; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_936 = fb_reg_valid ? _GEN_296 : btb_target_40; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_937 = fb_reg_valid ? _GEN_297 : btb_target_41; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_938 = fb_reg_valid ? _GEN_298 : btb_target_42; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_939 = fb_reg_valid ? _GEN_299 : btb_target_43; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_940 = fb_reg_valid ? _GEN_300 : btb_target_44; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_941 = fb_reg_valid ? _GEN_301 : btb_target_45; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_942 = fb_reg_valid ? _GEN_302 : btb_target_46; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_943 = fb_reg_valid ? _GEN_303 : btb_target_47; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_944 = fb_reg_valid ? _GEN_304 : btb_target_48; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_945 = fb_reg_valid ? _GEN_305 : btb_target_49; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_946 = fb_reg_valid ? _GEN_306 : btb_target_50; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_947 = fb_reg_valid ? _GEN_307 : btb_target_51; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_948 = fb_reg_valid ? _GEN_308 : btb_target_52; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_949 = fb_reg_valid ? _GEN_309 : btb_target_53; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_950 = fb_reg_valid ? _GEN_310 : btb_target_54; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_951 = fb_reg_valid ? _GEN_311 : btb_target_55; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_952 = fb_reg_valid ? _GEN_312 : btb_target_56; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_953 = fb_reg_valid ? _GEN_313 : btb_target_57; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_954 = fb_reg_valid ? _GEN_314 : btb_target_58; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_955 = fb_reg_valid ? _GEN_315 : btb_target_59; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_956 = fb_reg_valid ? _GEN_316 : btb_target_60; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_957 = fb_reg_valid ? _GEN_317 : btb_target_61; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_958 = fb_reg_valid ? _GEN_318 : btb_target_62; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_959 = fb_reg_valid ? _GEN_319 : btb_target_63; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_960 = fb_reg_valid ? _GEN_320 : btb_btype_0; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_961 = fb_reg_valid ? _GEN_321 : btb_btype_1; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_962 = fb_reg_valid ? _GEN_322 : btb_btype_2; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_963 = fb_reg_valid ? _GEN_323 : btb_btype_3; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_964 = fb_reg_valid ? _GEN_324 : btb_btype_4; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_965 = fb_reg_valid ? _GEN_325 : btb_btype_5; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_966 = fb_reg_valid ? _GEN_326 : btb_btype_6; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_967 = fb_reg_valid ? _GEN_327 : btb_btype_7; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_968 = fb_reg_valid ? _GEN_328 : btb_btype_8; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_969 = fb_reg_valid ? _GEN_329 : btb_btype_9; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_970 = fb_reg_valid ? _GEN_330 : btb_btype_10; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_971 = fb_reg_valid ? _GEN_331 : btb_btype_11; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_972 = fb_reg_valid ? _GEN_332 : btb_btype_12; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_973 = fb_reg_valid ? _GEN_333 : btb_btype_13; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_974 = fb_reg_valid ? _GEN_334 : btb_btype_14; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_975 = fb_reg_valid ? _GEN_335 : btb_btype_15; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_976 = fb_reg_valid ? _GEN_336 : btb_btype_16; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_977 = fb_reg_valid ? _GEN_337 : btb_btype_17; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_978 = fb_reg_valid ? _GEN_338 : btb_btype_18; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_979 = fb_reg_valid ? _GEN_339 : btb_btype_19; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_980 = fb_reg_valid ? _GEN_340 : btb_btype_20; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_981 = fb_reg_valid ? _GEN_341 : btb_btype_21; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_982 = fb_reg_valid ? _GEN_342 : btb_btype_22; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_983 = fb_reg_valid ? _GEN_343 : btb_btype_23; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_984 = fb_reg_valid ? _GEN_344 : btb_btype_24; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_985 = fb_reg_valid ? _GEN_345 : btb_btype_25; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_986 = fb_reg_valid ? _GEN_346 : btb_btype_26; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_987 = fb_reg_valid ? _GEN_347 : btb_btype_27; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_988 = fb_reg_valid ? _GEN_348 : btb_btype_28; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_989 = fb_reg_valid ? _GEN_349 : btb_btype_29; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_990 = fb_reg_valid ? _GEN_350 : btb_btype_30; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_991 = fb_reg_valid ? _GEN_351 : btb_btype_31; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_992 = fb_reg_valid ? _GEN_352 : btb_btype_32; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_993 = fb_reg_valid ? _GEN_353 : btb_btype_33; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_994 = fb_reg_valid ? _GEN_354 : btb_btype_34; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_995 = fb_reg_valid ? _GEN_355 : btb_btype_35; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_996 = fb_reg_valid ? _GEN_356 : btb_btype_36; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_997 = fb_reg_valid ? _GEN_357 : btb_btype_37; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_998 = fb_reg_valid ? _GEN_358 : btb_btype_38; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_999 = fb_reg_valid ? _GEN_359 : btb_btype_39; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1000 = fb_reg_valid ? _GEN_360 : btb_btype_40; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1001 = fb_reg_valid ? _GEN_361 : btb_btype_41; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1002 = fb_reg_valid ? _GEN_362 : btb_btype_42; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1003 = fb_reg_valid ? _GEN_363 : btb_btype_43; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1004 = fb_reg_valid ? _GEN_364 : btb_btype_44; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1005 = fb_reg_valid ? _GEN_365 : btb_btype_45; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1006 = fb_reg_valid ? _GEN_366 : btb_btype_46; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1007 = fb_reg_valid ? _GEN_367 : btb_btype_47; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1008 = fb_reg_valid ? _GEN_368 : btb_btype_48; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1009 = fb_reg_valid ? _GEN_369 : btb_btype_49; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1010 = fb_reg_valid ? _GEN_370 : btb_btype_50; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1011 = fb_reg_valid ? _GEN_371 : btb_btype_51; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1012 = fb_reg_valid ? _GEN_372 : btb_btype_52; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1013 = fb_reg_valid ? _GEN_373 : btb_btype_53; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1014 = fb_reg_valid ? _GEN_374 : btb_btype_54; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1015 = fb_reg_valid ? _GEN_375 : btb_btype_55; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1016 = fb_reg_valid ? _GEN_376 : btb_btype_56; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1017 = fb_reg_valid ? _GEN_377 : btb_btype_57; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1018 = fb_reg_valid ? _GEN_378 : btb_btype_58; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1019 = fb_reg_valid ? _GEN_379 : btb_btype_59; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1020 = fb_reg_valid ? _GEN_380 : btb_btype_60; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1021 = fb_reg_valid ? _GEN_381 : btb_btype_61; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1022 = fb_reg_valid ? _GEN_382 : btb_btype_62; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1023 = fb_reg_valid ? _GEN_383 : btb_btype_63; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1024 = fb_reg_valid ? _GEN_768 : btb_hcount_0; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1025 = fb_reg_valid ? _GEN_769 : btb_hcount_1; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1026 = fb_reg_valid ? _GEN_770 : btb_hcount_2; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1027 = fb_reg_valid ? _GEN_771 : btb_hcount_3; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1028 = fb_reg_valid ? _GEN_772 : btb_hcount_4; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1029 = fb_reg_valid ? _GEN_773 : btb_hcount_5; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1030 = fb_reg_valid ? _GEN_774 : btb_hcount_6; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1031 = fb_reg_valid ? _GEN_775 : btb_hcount_7; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1032 = fb_reg_valid ? _GEN_776 : btb_hcount_8; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1033 = fb_reg_valid ? _GEN_777 : btb_hcount_9; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1034 = fb_reg_valid ? _GEN_778 : btb_hcount_10; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1035 = fb_reg_valid ? _GEN_779 : btb_hcount_11; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1036 = fb_reg_valid ? _GEN_780 : btb_hcount_12; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1037 = fb_reg_valid ? _GEN_781 : btb_hcount_13; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1038 = fb_reg_valid ? _GEN_782 : btb_hcount_14; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1039 = fb_reg_valid ? _GEN_783 : btb_hcount_15; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1040 = fb_reg_valid ? _GEN_784 : btb_hcount_16; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1041 = fb_reg_valid ? _GEN_785 : btb_hcount_17; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1042 = fb_reg_valid ? _GEN_786 : btb_hcount_18; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1043 = fb_reg_valid ? _GEN_787 : btb_hcount_19; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1044 = fb_reg_valid ? _GEN_788 : btb_hcount_20; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1045 = fb_reg_valid ? _GEN_789 : btb_hcount_21; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1046 = fb_reg_valid ? _GEN_790 : btb_hcount_22; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1047 = fb_reg_valid ? _GEN_791 : btb_hcount_23; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1048 = fb_reg_valid ? _GEN_792 : btb_hcount_24; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1049 = fb_reg_valid ? _GEN_793 : btb_hcount_25; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1050 = fb_reg_valid ? _GEN_794 : btb_hcount_26; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1051 = fb_reg_valid ? _GEN_795 : btb_hcount_27; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1052 = fb_reg_valid ? _GEN_796 : btb_hcount_28; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1053 = fb_reg_valid ? _GEN_797 : btb_hcount_29; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1054 = fb_reg_valid ? _GEN_798 : btb_hcount_30; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1055 = fb_reg_valid ? _GEN_799 : btb_hcount_31; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1056 = fb_reg_valid ? _GEN_800 : btb_hcount_32; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1057 = fb_reg_valid ? _GEN_801 : btb_hcount_33; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1058 = fb_reg_valid ? _GEN_802 : btb_hcount_34; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1059 = fb_reg_valid ? _GEN_803 : btb_hcount_35; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1060 = fb_reg_valid ? _GEN_804 : btb_hcount_36; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1061 = fb_reg_valid ? _GEN_805 : btb_hcount_37; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1062 = fb_reg_valid ? _GEN_806 : btb_hcount_38; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1063 = fb_reg_valid ? _GEN_807 : btb_hcount_39; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1064 = fb_reg_valid ? _GEN_808 : btb_hcount_40; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1065 = fb_reg_valid ? _GEN_809 : btb_hcount_41; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1066 = fb_reg_valid ? _GEN_810 : btb_hcount_42; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1067 = fb_reg_valid ? _GEN_811 : btb_hcount_43; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1068 = fb_reg_valid ? _GEN_812 : btb_hcount_44; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1069 = fb_reg_valid ? _GEN_813 : btb_hcount_45; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1070 = fb_reg_valid ? _GEN_814 : btb_hcount_46; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1071 = fb_reg_valid ? _GEN_815 : btb_hcount_47; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1072 = fb_reg_valid ? _GEN_816 : btb_hcount_48; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1073 = fb_reg_valid ? _GEN_817 : btb_hcount_49; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1074 = fb_reg_valid ? _GEN_818 : btb_hcount_50; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1075 = fb_reg_valid ? _GEN_819 : btb_hcount_51; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1076 = fb_reg_valid ? _GEN_820 : btb_hcount_52; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1077 = fb_reg_valid ? _GEN_821 : btb_hcount_53; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1078 = fb_reg_valid ? _GEN_822 : btb_hcount_54; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1079 = fb_reg_valid ? _GEN_823 : btb_hcount_55; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1080 = fb_reg_valid ? _GEN_824 : btb_hcount_56; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1081 = fb_reg_valid ? _GEN_825 : btb_hcount_57; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1082 = fb_reg_valid ? _GEN_826 : btb_hcount_58; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1083 = fb_reg_valid ? _GEN_827 : btb_hcount_59; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1084 = fb_reg_valid ? _GEN_828 : btb_hcount_60; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1085 = fb_reg_valid ? _GEN_829 : btb_hcount_61; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1086 = fb_reg_valid ? _GEN_830 : btb_hcount_62; // @[BTB.scala 130:23:@4328.4]
  assign _GEN_1087 = fb_reg_valid ? _GEN_831 : btb_hcount_63; // @[BTB.scala 130:23:@4328.4]
  assign io_pred_pc_0 = _T_1391 ? io_ras_peek : _T_1403; // @[BTB.scala 80:20:@2184.4]
  assign io_pred_pc_1 = _T_2644 ? io_ras_peek : _T_2656; // @[BTB.scala 80:20:@3167.4]
  assign io_split = _T_1402 & _T_2675; // @[BTB.scala 85:12:@3183.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_pc_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  btb_pc_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  btb_pc_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  btb_pc_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  btb_pc_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  btb_pc_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  btb_pc_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  btb_pc_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  btb_pc_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  btb_pc_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  btb_pc_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  btb_pc_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  btb_pc_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  btb_pc_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  btb_pc_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  btb_pc_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  btb_pc_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  btb_pc_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  btb_pc_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  btb_pc_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  btb_pc_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  btb_pc_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  btb_pc_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  btb_pc_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  btb_pc_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  btb_pc_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  btb_pc_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  btb_pc_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  btb_pc_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  btb_pc_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  btb_pc_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  btb_pc_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  btb_pc_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  btb_pc_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  btb_pc_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  btb_pc_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  btb_pc_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  btb_pc_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  btb_pc_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  btb_pc_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  btb_pc_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  btb_pc_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  btb_pc_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  btb_pc_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  btb_pc_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  btb_pc_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  btb_pc_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  btb_pc_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  btb_pc_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  btb_pc_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  btb_pc_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  btb_pc_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  btb_pc_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  btb_pc_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  btb_pc_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  btb_pc_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  btb_pc_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  btb_pc_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  btb_pc_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  btb_pc_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  btb_pc_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  btb_pc_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  btb_pc_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  btb_pc_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  btb_target_0 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  btb_target_1 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  btb_target_2 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  btb_target_3 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  btb_target_4 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  btb_target_5 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  btb_target_6 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  btb_target_7 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  btb_target_8 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  btb_target_9 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  btb_target_10 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  btb_target_11 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  btb_target_12 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  btb_target_13 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  btb_target_14 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  btb_target_15 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  btb_target_16 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  btb_target_17 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  btb_target_18 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  btb_target_19 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  btb_target_20 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  btb_target_21 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  btb_target_22 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  btb_target_23 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  btb_target_24 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  btb_target_25 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  btb_target_26 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  btb_target_27 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  btb_target_28 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  btb_target_29 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  btb_target_30 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  btb_target_31 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  btb_target_32 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  btb_target_33 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  btb_target_34 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  btb_target_35 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  btb_target_36 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  btb_target_37 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  btb_target_38 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  btb_target_39 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  btb_target_40 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  btb_target_41 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  btb_target_42 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  btb_target_43 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  btb_target_44 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  btb_target_45 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  btb_target_46 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  btb_target_47 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  btb_target_48 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  btb_target_49 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  btb_target_50 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  btb_target_51 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  btb_target_52 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  btb_target_53 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  btb_target_54 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  btb_target_55 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  btb_target_56 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  btb_target_57 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  btb_target_58 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  btb_target_59 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  btb_target_60 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  btb_target_61 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  btb_target_62 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  btb_target_63 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  btb_hcount_0 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  btb_hcount_1 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  btb_hcount_2 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  btb_hcount_3 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  btb_hcount_4 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  btb_hcount_5 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  btb_hcount_6 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  btb_hcount_7 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  btb_hcount_8 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  btb_hcount_9 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  btb_hcount_10 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  btb_hcount_11 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  btb_hcount_12 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  btb_hcount_13 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  btb_hcount_14 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  btb_hcount_15 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  btb_hcount_16 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  btb_hcount_17 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  btb_hcount_18 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  btb_hcount_19 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  btb_hcount_20 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  btb_hcount_21 = _RAND_149[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  btb_hcount_22 = _RAND_150[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  btb_hcount_23 = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  btb_hcount_24 = _RAND_152[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  btb_hcount_25 = _RAND_153[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  btb_hcount_26 = _RAND_154[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  btb_hcount_27 = _RAND_155[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  btb_hcount_28 = _RAND_156[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  btb_hcount_29 = _RAND_157[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  btb_hcount_30 = _RAND_158[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  btb_hcount_31 = _RAND_159[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  btb_hcount_32 = _RAND_160[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  btb_hcount_33 = _RAND_161[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  btb_hcount_34 = _RAND_162[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  btb_hcount_35 = _RAND_163[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  btb_hcount_36 = _RAND_164[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  btb_hcount_37 = _RAND_165[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  btb_hcount_38 = _RAND_166[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  btb_hcount_39 = _RAND_167[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  btb_hcount_40 = _RAND_168[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  btb_hcount_41 = _RAND_169[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  btb_hcount_42 = _RAND_170[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  btb_hcount_43 = _RAND_171[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  btb_hcount_44 = _RAND_172[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  btb_hcount_45 = _RAND_173[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  btb_hcount_46 = _RAND_174[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  btb_hcount_47 = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  btb_hcount_48 = _RAND_176[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  btb_hcount_49 = _RAND_177[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  btb_hcount_50 = _RAND_178[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  btb_hcount_51 = _RAND_179[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  btb_hcount_52 = _RAND_180[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  btb_hcount_53 = _RAND_181[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  btb_hcount_54 = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  btb_hcount_55 = _RAND_183[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  btb_hcount_56 = _RAND_184[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  btb_hcount_57 = _RAND_185[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  btb_hcount_58 = _RAND_186[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  btb_hcount_59 = _RAND_187[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  btb_hcount_60 = _RAND_188[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  btb_hcount_61 = _RAND_189[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  btb_hcount_62 = _RAND_190[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  btb_hcount_63 = _RAND_191[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  btb_btype_0 = _RAND_192[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  btb_btype_1 = _RAND_193[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  btb_btype_2 = _RAND_194[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  btb_btype_3 = _RAND_195[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  btb_btype_4 = _RAND_196[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  btb_btype_5 = _RAND_197[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  btb_btype_6 = _RAND_198[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  btb_btype_7 = _RAND_199[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  btb_btype_8 = _RAND_200[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  btb_btype_9 = _RAND_201[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  btb_btype_10 = _RAND_202[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  btb_btype_11 = _RAND_203[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  btb_btype_12 = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  btb_btype_13 = _RAND_205[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  btb_btype_14 = _RAND_206[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  btb_btype_15 = _RAND_207[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  btb_btype_16 = _RAND_208[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  btb_btype_17 = _RAND_209[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  btb_btype_18 = _RAND_210[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  btb_btype_19 = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  btb_btype_20 = _RAND_212[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  btb_btype_21 = _RAND_213[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  btb_btype_22 = _RAND_214[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  btb_btype_23 = _RAND_215[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  btb_btype_24 = _RAND_216[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  btb_btype_25 = _RAND_217[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  btb_btype_26 = _RAND_218[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  btb_btype_27 = _RAND_219[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  btb_btype_28 = _RAND_220[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  btb_btype_29 = _RAND_221[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  btb_btype_30 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  btb_btype_31 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  btb_btype_32 = _RAND_224[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  btb_btype_33 = _RAND_225[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  btb_btype_34 = _RAND_226[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  btb_btype_35 = _RAND_227[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  btb_btype_36 = _RAND_228[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  btb_btype_37 = _RAND_229[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  btb_btype_38 = _RAND_230[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  btb_btype_39 = _RAND_231[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  btb_btype_40 = _RAND_232[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  btb_btype_41 = _RAND_233[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  btb_btype_42 = _RAND_234[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  btb_btype_43 = _RAND_235[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  btb_btype_44 = _RAND_236[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  btb_btype_45 = _RAND_237[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  btb_btype_46 = _RAND_238[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  btb_btype_47 = _RAND_239[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  btb_btype_48 = _RAND_240[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  btb_btype_49 = _RAND_241[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  btb_btype_50 = _RAND_242[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  btb_btype_51 = _RAND_243[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  btb_btype_52 = _RAND_244[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  btb_btype_53 = _RAND_245[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  btb_btype_54 = _RAND_246[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  btb_btype_55 = _RAND_247[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  btb_btype_56 = _RAND_248[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  btb_btype_57 = _RAND_249[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  btb_btype_58 = _RAND_250[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  btb_btype_59 = _RAND_251[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  btb_btype_60 = _RAND_252[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  btb_btype_61 = _RAND_253[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  btb_btype_62 = _RAND_254[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  btb_btype_63 = _RAND_255[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  fb_reg_valid = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  fb_reg_redirect = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  fb_reg_lfsr = _RAND_258[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  fb_reg_pc = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  fb_reg_target = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  fb_reg_btype = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      btb_pc_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_pc_0 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_pc_1 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_pc_2 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_pc_3 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_pc_4 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_pc_5 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_pc_6 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_pc_7 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_pc_8 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_pc_9 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_pc_10 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_pc_11 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_pc_12 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_pc_13 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_pc_14 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_pc_15 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_pc_16 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_pc_17 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_pc_18 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_pc_19 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_pc_20 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_pc_21 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_pc_22 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_pc_23 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_pc_24 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_pc_25 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_pc_26 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_pc_27 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_pc_28 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_pc_29 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_pc_30 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_pc_31 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_pc_32 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_pc_33 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_pc_34 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_pc_35 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_pc_36 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_pc_37 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_pc_38 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_pc_39 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_pc_40 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_pc_41 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_pc_42 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_pc_43 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_pc_44 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_pc_45 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_pc_46 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_pc_47 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_pc_48 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_pc_49 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_pc_50 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_pc_51 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_pc_52 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_pc_53 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_pc_54 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_pc_55 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_pc_56 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_pc_57 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_pc_58 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_pc_59 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_pc_60 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_pc_61 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_pc_62 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_pc_63 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_target_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_target_0 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_target_1 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_target_2 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_target_3 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_target_4 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_target_5 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_target_6 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_target_7 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_target_8 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_target_9 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_target_10 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_target_11 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_target_12 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_target_13 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_target_14 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_target_15 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_target_16 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_target_17 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_target_18 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_target_19 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_target_20 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_target_21 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_target_22 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_target_23 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_target_24 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_target_25 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_target_26 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_target_27 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_target_28 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_target_29 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_target_30 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_target_31 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_target_32 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_target_33 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_target_34 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_target_35 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_target_36 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_target_37 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_target_38 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_target_39 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_target_40 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_target_41 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_target_42 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_target_43 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_target_44 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_target_45 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_target_46 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_target_47 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_target_48 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_target_49 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_target_50 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_target_51 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_target_52 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_target_53 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_target_54 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_target_55 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_target_56 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_target_57 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_target_58 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_target_59 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_target_60 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_target_61 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_target_62 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_target_63 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= _T_4169;
              end
            end else begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= _T_4169;
              end
            end else begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= _T_4169;
              end
            end else begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= _T_4169;
              end
            end else begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= _T_4169;
              end
            end else begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= _T_4169;
              end
            end else begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= _T_4169;
              end
            end else begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= _T_4169;
              end
            end else begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= _T_4169;
              end
            end else begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= _T_4169;
              end
            end else begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= _T_4169;
              end
            end else begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= _T_4169;
              end
            end else begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= _T_4169;
              end
            end else begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= _T_4169;
              end
            end else begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= _T_4169;
              end
            end else begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= _T_4169;
              end
            end else begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= _T_4169;
              end
            end else begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= _T_4169;
              end
            end else begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= _T_4169;
              end
            end else begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= _T_4169;
              end
            end else begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= _T_4169;
              end
            end else begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= _T_4169;
              end
            end else begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= _T_4169;
              end
            end else begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= _T_4169;
              end
            end else begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= _T_4169;
              end
            end else begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= _T_4169;
              end
            end else begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= _T_4169;
              end
            end else begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= _T_4169;
              end
            end else begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= _T_4169;
              end
            end else begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= _T_4169;
              end
            end else begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= _T_4169;
              end
            end else begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= _T_4169;
              end
            end else begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= _T_4169;
              end
            end else begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= _T_4169;
              end
            end else begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= _T_4169;
              end
            end else begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= _T_4169;
              end
            end else begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= _T_4169;
              end
            end else begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= _T_4169;
              end
            end else begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= _T_4169;
              end
            end else begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= _T_4169;
              end
            end else begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= _T_4169;
              end
            end else begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= _T_4169;
              end
            end else begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= _T_4169;
              end
            end else begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= _T_4169;
              end
            end else begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= _T_4169;
              end
            end else begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= _T_4169;
              end
            end else begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= _T_4169;
              end
            end else begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= _T_4169;
              end
            end else begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= _T_4169;
              end
            end else begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= _T_4169;
              end
            end else begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= _T_4169;
              end
            end else begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= _T_4169;
              end
            end else begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= _T_4169;
              end
            end else begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= _T_4169;
              end
            end else begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= _T_4169;
              end
            end else begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= _T_4169;
              end
            end else begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= _T_4169;
              end
            end else begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= _T_4169;
              end
            end else begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= _T_4169;
              end
            end else begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= _T_4169;
              end
            end else begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= _T_4169;
              end
            end else begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= _T_4169;
              end
            end else begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= _T_4169;
              end
            end else begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_4159) begin
          if (_T_3407) begin
            if (fb_reg_redirect) begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= _T_4169;
              end
            end else begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= _T_4178;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_btype_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_btype_0 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_btype_1 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_btype_2 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_btype_3 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_btype_4 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_btype_5 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_btype_6 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_btype_7 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_btype_8 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_btype_9 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_btype_10 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_btype_11 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_btype_12 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_btype_13 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_btype_14 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_btype_15 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_btype_16 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_btype_17 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_btype_18 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_btype_19 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_btype_20 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_btype_21 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_btype_22 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_btype_23 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_btype_24 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_btype_25 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_btype_26 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_btype_27 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_btype_28 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_btype_29 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_btype_30 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_btype_31 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_btype_32 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_btype_33 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_btype_34 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_btype_35 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_btype_36 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_btype_37 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_btype_38 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_btype_39 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_btype_40 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_btype_41 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_btype_42 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_btype_43 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_btype_44 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_btype_45 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_btype_46 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_btype_47 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_btype_48 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_btype_49 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_btype_50 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_btype_51 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_btype_52 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_btype_53 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_btype_54 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_btype_55 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_btype_56 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_btype_57 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_btype_58 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_btype_59 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_btype_60 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_btype_61 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_btype_62 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_btype_63 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      fb_reg_valid <= 1'h0;
    end else begin
      fb_reg_valid <= io_feedBack_valid;
    end
    if (reset) begin
      fb_reg_redirect <= 1'h0;
    end else begin
      fb_reg_redirect <= io_feedBack_bits_redirect;
    end
    if (reset) begin
      fb_reg_lfsr <= 6'h1;
    end else begin
      fb_reg_lfsr <= _T_2687;
    end
    if (reset) begin
      fb_reg_pc <= 32'h0;
    end else begin
      fb_reg_pc <= io_fb_pc;
    end
    if (reset) begin
      fb_reg_target <= 32'h0;
    end else begin
      fb_reg_target <= io_feedBack_bits_tgt;
    end
    if (reset) begin
      fb_reg_btype <= 2'h0;
    end else begin
      fb_reg_btype <= io_fb_type;
    end
  end
endmodule
module RAS( // @[:@4365.2]
  input         clock, // @[:@4366.4]
  input         reset, // @[:@4367.4]
  input         io_push_valid, // @[:@4368.4]
  input  [31:0] io_push_bits, // @[:@4368.4]
  input         io_pop, // @[:@4368.4]
  output [31:0] io_peek // @[:@4368.4]
);
  reg [31:0] stack [0:15]; // @[RAS.scala 13:18:@4370.4]
  reg [31:0] _RAND_0;
  wire [31:0] stack__T_23_data; // @[RAS.scala 13:18:@4370.4]
  wire [3:0] stack__T_23_addr; // @[RAS.scala 13:18:@4370.4]
  wire [31:0] stack__T_24_data; // @[RAS.scala 13:18:@4370.4]
  wire [3:0] stack__T_24_addr; // @[RAS.scala 13:18:@4370.4]
  wire  stack__T_24_mask; // @[RAS.scala 13:18:@4370.4]
  wire  stack__T_24_en; // @[RAS.scala 13:18:@4370.4]
  wire [31:0] stack__T_25_data; // @[RAS.scala 13:18:@4370.4]
  wire [3:0] stack__T_25_addr; // @[RAS.scala 13:18:@4370.4]
  wire  stack__T_25_mask; // @[RAS.scala 13:18:@4370.4]
  wire  stack__T_25_en; // @[RAS.scala 13:18:@4370.4]
  reg [3:0] pos; // @[RAS.scala 14:22:@4371.4]
  reg [31:0] _RAND_1;
  reg [3:0] next; // @[RAS.scala 15:22:@4372.4]
  reg [31:0] _RAND_2;
  wire  _GEN_7; // @[RAS.scala 19:18:@4376.6]
  wire  _T_27; // @[RAS.scala 26:26:@4385.4]
  wire  _T_28; // @[RAS.scala 26:23:@4386.4]
  wire [4:0] _T_30; // @[RAS.scala 27:18:@4388.6]
  wire [3:0] _T_31; // @[RAS.scala 27:18:@4389.6]
  wire [4:0] _T_33; // @[RAS.scala 28:18:@4391.6]
  wire [3:0] _T_34; // @[RAS.scala 28:18:@4392.6]
  wire [4:0] _T_36; // @[RAS.scala 31:18:@4397.8]
  wire [4:0] _T_37; // @[RAS.scala 31:18:@4398.8]
  wire [3:0] _T_38; // @[RAS.scala 31:18:@4399.8]
  wire [4:0] _T_40; // @[RAS.scala 32:18:@4401.8]
  wire [4:0] _T_41; // @[RAS.scala 32:18:@4402.8]
  wire [3:0] _T_42; // @[RAS.scala 32:18:@4403.8]
  wire [3:0] _GEN_20; // @[RAS.scala 29:22:@4396.6]
  wire [3:0] _GEN_21; // @[RAS.scala 29:22:@4396.6]
  wire [3:0] _GEN_22; // @[RAS.scala 26:35:@4387.4]
  wire [3:0] _GEN_23; // @[RAS.scala 26:35:@4387.4]
  assign stack__T_23_addr = pos;
  assign stack__T_23_data = stack[stack__T_23_addr]; // @[RAS.scala 13:18:@4370.4]
  assign stack__T_24_data = io_push_bits;
  assign stack__T_24_addr = pos;
  assign stack__T_24_mask = 1'h1;
  assign stack__T_24_en = io_push_valid ? io_pop : 1'h0;
  assign stack__T_25_data = io_push_bits;
  assign stack__T_25_addr = next;
  assign stack__T_25_mask = 1'h1;
  assign stack__T_25_en = io_push_valid ? _GEN_7 : 1'h0;
  assign _GEN_7 = io_pop ? 1'h0 : 1'h1; // @[RAS.scala 19:18:@4376.6]
  assign _T_27 = io_pop == 1'h0; // @[RAS.scala 26:26:@4385.4]
  assign _T_28 = io_push_valid & _T_27; // @[RAS.scala 26:23:@4386.4]
  assign _T_30 = pos + 4'h1; // @[RAS.scala 27:18:@4388.6]
  assign _T_31 = pos + 4'h1; // @[RAS.scala 27:18:@4389.6]
  assign _T_33 = next + 4'h1; // @[RAS.scala 28:18:@4391.6]
  assign _T_34 = next + 4'h1; // @[RAS.scala 28:18:@4392.6]
  assign _T_36 = pos - 4'h1; // @[RAS.scala 31:18:@4397.8]
  assign _T_37 = $unsigned(_T_36); // @[RAS.scala 31:18:@4398.8]
  assign _T_38 = _T_37[3:0]; // @[RAS.scala 31:18:@4399.8]
  assign _T_40 = next - 4'h1; // @[RAS.scala 32:18:@4401.8]
  assign _T_41 = $unsigned(_T_40); // @[RAS.scala 32:18:@4402.8]
  assign _T_42 = _T_41[3:0]; // @[RAS.scala 32:18:@4403.8]
  assign _GEN_20 = io_pop ? _T_38 : pos; // @[RAS.scala 29:22:@4396.6]
  assign _GEN_21 = io_pop ? _T_42 : next; // @[RAS.scala 29:22:@4396.6]
  assign _GEN_22 = _T_28 ? _T_31 : _GEN_20; // @[RAS.scala 26:35:@4387.4]
  assign _GEN_23 = _T_28 ? _T_34 : _GEN_21; // @[RAS.scala 26:35:@4387.4]
  assign io_peek = stack__T_23_data; // @[RAS.scala 16:11:@4374.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    stack[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pos = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  next = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(stack__T_24_en & stack__T_24_mask) begin
      stack[stack__T_24_addr] <= stack__T_24_data; // @[RAS.scala 13:18:@4370.4]
    end
    if(stack__T_25_en & stack__T_25_mask) begin
      stack[stack__T_25_addr] <= stack__T_25_data; // @[RAS.scala 13:18:@4370.4]
    end
    if (reset) begin
      pos <= 4'hf;
    end else begin
      if (_T_28) begin
        pos <= _T_31;
      end else begin
        if (io_pop) begin
          pos <= _T_38;
        end
      end
    end
    if (reset) begin
      next <= 4'h0;
    end else begin
      if (_T_28) begin
        next <= _T_34;
      end else begin
        if (io_pop) begin
          next <= _T_42;
        end
      end
    end
  end
endmodule
module FrontEnd( // @[:@4407.2]
  input         clock, // @[:@4408.4]
  input         reset, // @[:@4409.4]
  input  [31:0] io_cyc, // @[:@4410.4]
  input         io_mem_addr_ready, // @[:@4410.4]
  output        io_mem_addr_valid, // @[:@4410.4]
  output [31:0] io_mem_addr_bits, // @[:@4410.4]
  input         io_mem_inst_0_valid, // @[:@4410.4]
  input  [31:0] io_mem_inst_0_bits, // @[:@4410.4]
  input         io_mem_inst_1_valid, // @[:@4410.4]
  input  [31:0] io_mem_inst_1_bits, // @[:@4410.4]
  input         io_back_xcpt_valid, // @[:@4410.4]
  input  [31:0] io_back_xcpt_bits, // @[:@4410.4]
  input         io_back_kill, // @[:@4410.4]
  input         io_back_fence, // @[:@4410.4]
  input         io_back_ras_pop, // @[:@4410.4]
  input         io_back_ras_push_valid, // @[:@4410.4]
  input  [31:0] io_back_ras_push_bits, // @[:@4410.4]
  input  [31:0] io_back_fb_pc, // @[:@4410.4]
  input  [1:0]  io_back_fb_type, // @[:@4410.4]
  input         io_back_feedBack_valid, // @[:@4410.4]
  input         io_back_feedBack_bits_redirect, // @[:@4410.4]
  input  [31:0] io_back_feedBack_bits_tgt, // @[:@4410.4]
  input         io_back_forward_0, // @[:@4410.4]
  input         io_back_forward_1, // @[:@4410.4]
  output        io_back_inst_0_valid, // @[:@4410.4]
  output [31:0] io_back_inst_0_bits, // @[:@4410.4]
  output        io_back_inst_1_valid, // @[:@4410.4]
  output [31:0] io_back_inst_1_bits, // @[:@4410.4]
  output [31:0] io_back_pc_0, // @[:@4410.4]
  output [31:0] io_back_pc_1, // @[:@4410.4]
  output [31:0] io_back_pred_0, // @[:@4410.4]
  output [31:0] io_back_pred_1 // @[:@4410.4]
);
  wire  FetchInst_clock; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_reset; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_cyc; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_mem_addr_ready; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_mem_addr_valid; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_mem_addr_bits; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_mem_inst_0_valid; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_mem_inst_0_bits; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_mem_inst_1_valid; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_mem_inst_1_bits; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_if_kill; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_if_fence; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_if_target; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_if_split; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_btb_target; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_forward_0; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_forward_1; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_kill_0; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_kill_1; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_if_pc; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_if_forward_0; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_if_forward_1; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_inst_0_valid; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_dec_inst_0_bits; // @[FrontEnd.scala 18:22:@4412.4]
  wire  FetchInst_io_dec_inst_1_valid; // @[FrontEnd.scala 18:22:@4412.4]
  wire [31:0] FetchInst_io_dec_inst_1_bits; // @[FrontEnd.scala 18:22:@4412.4]
  wire  BTB_clock; // @[FrontEnd.scala 20:22:@4416.4]
  wire  BTB_reset; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_if_pc; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_ras_peek; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_pred_pc_0; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_pred_pc_1; // @[FrontEnd.scala 20:22:@4416.4]
  wire  BTB_io_split; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_fb_pc; // @[FrontEnd.scala 20:22:@4416.4]
  wire [1:0] BTB_io_fb_type; // @[FrontEnd.scala 20:22:@4416.4]
  wire  BTB_io_feedBack_valid; // @[FrontEnd.scala 20:22:@4416.4]
  wire  BTB_io_feedBack_bits_redirect; // @[FrontEnd.scala 20:22:@4416.4]
  wire [31:0] BTB_io_feedBack_bits_tgt; // @[FrontEnd.scala 20:22:@4416.4]
  wire  RAS_clock; // @[FrontEnd.scala 22:22:@4420.4]
  wire  RAS_reset; // @[FrontEnd.scala 22:22:@4420.4]
  wire  RAS_io_push_valid; // @[FrontEnd.scala 22:22:@4420.4]
  wire [31:0] RAS_io_push_bits; // @[FrontEnd.scala 22:22:@4420.4]
  wire  RAS_io_pop; // @[FrontEnd.scala 22:22:@4420.4]
  wire [31:0] RAS_io_peek; // @[FrontEnd.scala 22:22:@4420.4]
  reg [31:0] dec_reg_pc_0; // @[FrontEnd.scala 45:23:@4453.4]
  reg [31:0] _RAND_0;
  reg [31:0] dec_reg_pc_1; // @[FrontEnd.scala 45:23:@4453.4]
  reg [31:0] _RAND_1;
  reg [31:0] dec_reg_pred_0; // @[FrontEnd.scala 46:25:@4454.4]
  reg [31:0] _RAND_2;
  reg [31:0] dec_reg_pred_1; // @[FrontEnd.scala 46:25:@4454.4]
  reg [31:0] _RAND_3;
  wire [28:0] _T_179; // @[FrontEnd.scala 9:13:@4456.6]
  wire [31:0] _T_183; // @[Cat.scala 30:58:@4458.6]
  wire [31:0] _T_188; // @[Cat.scala 30:58:@4465.6]
  FetchInst FetchInst ( // @[FrontEnd.scala 18:22:@4412.4]
    .clock(FetchInst_clock),
    .reset(FetchInst_reset),
    .io_cyc(FetchInst_io_cyc),
    .io_mem_addr_ready(FetchInst_io_mem_addr_ready),
    .io_mem_addr_valid(FetchInst_io_mem_addr_valid),
    .io_mem_addr_bits(FetchInst_io_mem_addr_bits),
    .io_mem_inst_0_valid(FetchInst_io_mem_inst_0_valid),
    .io_mem_inst_0_bits(FetchInst_io_mem_inst_0_bits),
    .io_mem_inst_1_valid(FetchInst_io_mem_inst_1_valid),
    .io_mem_inst_1_bits(FetchInst_io_mem_inst_1_bits),
    .io_if_kill(FetchInst_io_if_kill),
    .io_if_fence(FetchInst_io_if_fence),
    .io_if_target(FetchInst_io_if_target),
    .io_if_split(FetchInst_io_if_split),
    .io_btb_target(FetchInst_io_btb_target),
    .io_dec_forward_0(FetchInst_io_dec_forward_0),
    .io_dec_forward_1(FetchInst_io_dec_forward_1),
    .io_dec_kill_0(FetchInst_io_dec_kill_0),
    .io_dec_kill_1(FetchInst_io_dec_kill_1),
    .io_if_pc(FetchInst_io_if_pc),
    .io_if_forward_0(FetchInst_io_if_forward_0),
    .io_if_forward_1(FetchInst_io_if_forward_1),
    .io_dec_inst_0_valid(FetchInst_io_dec_inst_0_valid),
    .io_dec_inst_0_bits(FetchInst_io_dec_inst_0_bits),
    .io_dec_inst_1_valid(FetchInst_io_dec_inst_1_valid),
    .io_dec_inst_1_bits(FetchInst_io_dec_inst_1_bits)
  );
  BTB BTB ( // @[FrontEnd.scala 20:22:@4416.4]
    .clock(BTB_clock),
    .reset(BTB_reset),
    .io_if_pc(BTB_io_if_pc),
    .io_ras_peek(BTB_io_ras_peek),
    .io_pred_pc_0(BTB_io_pred_pc_0),
    .io_pred_pc_1(BTB_io_pred_pc_1),
    .io_split(BTB_io_split),
    .io_fb_pc(BTB_io_fb_pc),
    .io_fb_type(BTB_io_fb_type),
    .io_feedBack_valid(BTB_io_feedBack_valid),
    .io_feedBack_bits_redirect(BTB_io_feedBack_bits_redirect),
    .io_feedBack_bits_tgt(BTB_io_feedBack_bits_tgt)
  );
  RAS RAS ( // @[FrontEnd.scala 22:22:@4420.4]
    .clock(RAS_clock),
    .reset(RAS_reset),
    .io_push_valid(RAS_io_push_valid),
    .io_push_bits(RAS_io_push_bits),
    .io_pop(RAS_io_pop),
    .io_peek(RAS_io_peek)
  );
  assign _T_179 = FetchInst_io_if_pc[31:3]; // @[FrontEnd.scala 9:13:@4456.6]
  assign _T_183 = {_T_179,1'h0,2'h0}; // @[Cat.scala 30:58:@4458.6]
  assign _T_188 = {_T_179,1'h1,2'h0}; // @[Cat.scala 30:58:@4465.6]
  assign io_mem_addr_valid = FetchInst_io_mem_addr_valid; // @[FrontEnd.scala 24:14:@4428.4]
  assign io_mem_addr_bits = FetchInst_io_mem_addr_bits; // @[FrontEnd.scala 24:14:@4427.4]
  assign io_back_inst_0_valid = FetchInst_io_dec_inst_0_valid; // @[FrontEnd.scala 57:16:@4474.4]
  assign io_back_inst_0_bits = FetchInst_io_dec_inst_0_bits; // @[FrontEnd.scala 57:16:@4473.4]
  assign io_back_inst_1_valid = FetchInst_io_dec_inst_1_valid; // @[FrontEnd.scala 57:16:@4476.4]
  assign io_back_inst_1_bits = FetchInst_io_dec_inst_1_bits; // @[FrontEnd.scala 57:16:@4475.4]
  assign io_back_pc_0 = dec_reg_pc_0; // @[FrontEnd.scala 55:16:@4469.4]
  assign io_back_pc_1 = dec_reg_pc_1; // @[FrontEnd.scala 55:16:@4470.4]
  assign io_back_pred_0 = dec_reg_pred_0; // @[FrontEnd.scala 56:16:@4471.4]
  assign io_back_pred_1 = dec_reg_pred_1; // @[FrontEnd.scala 56:16:@4472.4]
  assign FetchInst_clock = clock; // @[:@4413.4]
  assign FetchInst_reset = reset; // @[:@4414.4]
  assign FetchInst_io_cyc = io_cyc; // @[FrontEnd.scala 19:14:@4415.4]
  assign FetchInst_io_mem_addr_ready = io_mem_addr_ready; // @[FrontEnd.scala 24:14:@4429.4]
  assign FetchInst_io_mem_inst_0_valid = io_mem_inst_0_valid; // @[FrontEnd.scala 24:14:@4424.4]
  assign FetchInst_io_mem_inst_0_bits = io_mem_inst_0_bits; // @[FrontEnd.scala 24:14:@4423.4]
  assign FetchInst_io_mem_inst_1_valid = io_mem_inst_1_valid; // @[FrontEnd.scala 24:14:@4426.4]
  assign FetchInst_io_mem_inst_1_bits = io_mem_inst_1_bits; // @[FrontEnd.scala 24:14:@4425.4]
  assign FetchInst_io_if_kill = FetchInst_io_dec_kill_1; // @[FrontEnd.scala 26:22:@4430.4]
  assign FetchInst_io_if_fence = io_back_fence; // @[FrontEnd.scala 27:22:@4431.4]
  assign FetchInst_io_if_target = io_back_xcpt_valid ? io_back_xcpt_bits : io_back_feedBack_bits_tgt; // @[FrontEnd.scala 28:22:@4433.4]
  assign FetchInst_io_if_split = BTB_io_split; // @[FrontEnd.scala 30:22:@4436.4]
  assign FetchInst_io_btb_target = BTB_io_split ? BTB_io_pred_pc_0 : BTB_io_pred_pc_1; // @[FrontEnd.scala 29:22:@4435.4]
  assign FetchInst_io_dec_forward_0 = io_back_forward_0; // @[FrontEnd.scala 32:22:@4437.4]
  assign FetchInst_io_dec_forward_1 = io_back_forward_1; // @[FrontEnd.scala 32:22:@4438.4]
  assign FetchInst_io_dec_kill_0 = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 33:22:@4440.4]
  assign FetchInst_io_dec_kill_1 = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 34:22:@4442.4]
  assign BTB_clock = clock; // @[:@4417.4]
  assign BTB_reset = reset; // @[:@4418.4]
  assign BTB_io_if_pc = FetchInst_io_if_pc; // @[FrontEnd.scala 39:16:@4446.4]
  assign BTB_io_ras_peek = RAS_io_peek; // @[FrontEnd.scala 40:16:@4447.4]
  assign BTB_io_fb_pc = io_back_fb_pc; // @[FrontEnd.scala 41:16:@4448.4]
  assign BTB_io_fb_type = io_back_fb_type; // @[FrontEnd.scala 42:16:@4449.4]
  assign BTB_io_feedBack_valid = io_back_feedBack_valid; // @[FrontEnd.scala 43:16:@4452.4]
  assign BTB_io_feedBack_bits_redirect = io_back_feedBack_bits_redirect; // @[FrontEnd.scala 43:16:@4451.4]
  assign BTB_io_feedBack_bits_tgt = io_back_feedBack_bits_tgt; // @[FrontEnd.scala 43:16:@4450.4]
  assign RAS_clock = clock; // @[:@4421.4]
  assign RAS_reset = reset; // @[:@4422.4]
  assign RAS_io_push_valid = io_back_ras_push_valid; // @[FrontEnd.scala 37:12:@4445.4]
  assign RAS_io_push_bits = io_back_ras_push_bits; // @[FrontEnd.scala 37:12:@4444.4]
  assign RAS_io_pop = io_back_ras_pop; // @[FrontEnd.scala 36:12:@4443.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dec_reg_pc_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dec_reg_pc_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  dec_reg_pred_0 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  dec_reg_pred_1 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (FetchInst_io_if_forward_0) begin
      dec_reg_pc_0 <= _T_183;
    end
    if (FetchInst_io_if_forward_1) begin
      dec_reg_pc_1 <= _T_188;
    end
    if (FetchInst_io_if_forward_0) begin
      dec_reg_pred_0 <= BTB_io_pred_pc_0;
    end
    if (FetchInst_io_if_forward_1) begin
      dec_reg_pred_1 <= BTB_io_pred_pc_1;
    end
  end
endmodule
module CSRFile( // @[:@4478.2]
  input         clock, // @[:@4479.4]
  input         reset, // @[:@4480.4]
  input  [2:0]  io_rw_cmd, // @[:@4481.4]
  input  [11:0] io_rw_addr, // @[:@4481.4]
  output [31:0] io_rw_rdata, // @[:@4481.4]
  input  [31:0] io_rw_wdata, // @[:@4481.4]
  output        io_eret, // @[:@4481.4]
  output [1:0]  io_status_prv, // @[:@4481.4]
  output [13:0] io_status_unimp5, // @[:@4481.4]
  output        io_status_mprv, // @[:@4481.4]
  output [1:0]  io_status_unimp4, // @[:@4481.4]
  output [1:0]  io_status_mpp, // @[:@4481.4]
  output [2:0]  io_status_unimp3, // @[:@4481.4]
  output        io_status_mpie, // @[:@4481.4]
  output [2:0]  io_status_unimp2, // @[:@4481.4]
  output        io_status_mie, // @[:@4481.4]
  output [2:0]  io_status_unimp1, // @[:@4481.4]
  input         io_xcpt, // @[:@4481.4]
  input  [31:0] io_cause, // @[:@4481.4]
  input  [31:0] io_tval, // @[:@4481.4]
  output [31:0] io_evec, // @[:@4481.4]
  input         io_illegal, // @[:@4481.4]
  input  [1:0]  io_retire, // @[:@4481.4]
  input  [31:0] io_pc, // @[:@4481.4]
  output [31:0] io_time // @[:@4481.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 112:28:@4608.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 112:28:@4608.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 112:28:@4608.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[CSR.scala 113:21:@4609.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[CSR.scala 114:23:@4610.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[CSR.scala 115:22:@4611.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[CSR.scala 116:25:@4612.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[CSR.scala 118:24:@4614.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[CSR.scala 120:24:@4632.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[CSR.scala 120:24:@4632.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[CSR.scala 121:24:@4650.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[CSR.scala 121:24:@4650.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_240; // @[Util.scala 112:41:@4653.4]
  reg [31:0] _RAND_12;
  wire [6:0] _T_241; // @[Util.scala 113:33:@4654.4]
  reg [57:0] _T_244; // @[Util.scala 117:31:@4656.4]
  reg [63:0] _RAND_13;
  wire  _T_245; // @[Util.scala 118:20:@4657.4]
  wire [58:0] _T_247; // @[Util.scala 118:43:@4659.6]
  wire [57:0] _T_248; // @[Util.scala 118:43:@4660.6]
  wire [57:0] _GEN_0; // @[Util.scala 118:34:@4658.4]
  wire [63:0] _T_249; // @[Cat.scala 30:58:@4663.4]
  reg [5:0] _T_252; // @[Util.scala 112:41:@4664.4]
  reg [31:0] _RAND_14;
  wire [5:0] _GEN_147; // @[Util.scala 113:33:@4665.4]
  wire [6:0] _T_253; // @[Util.scala 113:33:@4665.4]
  reg [57:0] _T_256; // @[Util.scala 117:31:@4667.4]
  reg [63:0] _RAND_15;
  wire  _T_257; // @[Util.scala 118:20:@4668.4]
  wire [58:0] _T_259; // @[Util.scala 118:43:@4670.6]
  wire [57:0] _T_260; // @[Util.scala 118:43:@4671.6]
  wire [57:0] _GEN_1; // @[Util.scala 118:34:@4669.4]
  wire [63:0] _T_261; // @[Cat.scala 30:58:@4674.4]
  reg [39:0] _T_264; // @[Util.scala 112:74:@4676.4]
  reg [63:0] _RAND_16;
  wire [40:0] _T_265; // @[Util.scala 113:33:@4677.4]
  reg [39:0] _T_267; // @[Util.scala 112:74:@4679.4]
  reg [63:0] _RAND_17;
  wire [40:0] _T_268; // @[Util.scala 113:33:@4680.4]
  reg [39:0] _T_270; // @[Util.scala 112:74:@4682.4]
  reg [63:0] _RAND_18;
  wire [40:0] _T_271; // @[Util.scala 113:33:@4683.4]
  reg [39:0] _T_273; // @[Util.scala 112:74:@4685.4]
  reg [63:0] _RAND_19;
  wire [40:0] _T_274; // @[Util.scala 113:33:@4686.4]
  reg [39:0] _T_276; // @[Util.scala 112:74:@4688.4]
  reg [63:0] _RAND_20;
  wire [40:0] _T_277; // @[Util.scala 113:33:@4689.4]
  reg [39:0] _T_279; // @[Util.scala 112:74:@4691.4]
  reg [63:0] _RAND_21;
  wire [40:0] _T_280; // @[Util.scala 113:33:@4692.4]
  reg [39:0] _T_282; // @[Util.scala 112:74:@4694.4]
  reg [63:0] _RAND_22;
  wire [40:0] _T_283; // @[Util.scala 113:33:@4695.4]
  reg [39:0] _T_285; // @[Util.scala 112:74:@4697.4]
  reg [63:0] _RAND_23;
  wire [40:0] _T_286; // @[Util.scala 113:33:@4698.4]
  reg [39:0] _T_288; // @[Util.scala 112:74:@4700.4]
  reg [63:0] _RAND_24;
  wire [40:0] _T_289; // @[Util.scala 113:33:@4701.4]
  reg [39:0] _T_291; // @[Util.scala 112:74:@4703.4]
  reg [63:0] _RAND_25;
  wire [40:0] _T_292; // @[Util.scala 113:33:@4704.4]
  reg [39:0] _T_294; // @[Util.scala 112:74:@4706.4]
  reg [63:0] _RAND_26;
  wire [40:0] _T_295; // @[Util.scala 113:33:@4707.4]
  reg [39:0] _T_297; // @[Util.scala 112:74:@4709.4]
  reg [63:0] _RAND_27;
  wire [40:0] _T_298; // @[Util.scala 113:33:@4710.4]
  reg [39:0] _T_300; // @[Util.scala 112:74:@4712.4]
  reg [63:0] _RAND_28;
  wire [40:0] _T_301; // @[Util.scala 113:33:@4713.4]
  reg [39:0] _T_303; // @[Util.scala 112:74:@4715.4]
  reg [63:0] _RAND_29;
  wire [40:0] _T_304; // @[Util.scala 113:33:@4716.4]
  reg [39:0] _T_306; // @[Util.scala 112:74:@4718.4]
  reg [63:0] _RAND_30;
  wire [40:0] _T_307; // @[Util.scala 113:33:@4719.4]
  reg [39:0] _T_309; // @[Util.scala 112:74:@4721.4]
  reg [63:0] _RAND_31;
  wire [40:0] _T_310; // @[Util.scala 113:33:@4722.4]
  reg [39:0] _T_312; // @[Util.scala 112:74:@4724.4]
  reg [63:0] _RAND_32;
  wire [40:0] _T_313; // @[Util.scala 113:33:@4725.4]
  reg [39:0] _T_315; // @[Util.scala 112:74:@4727.4]
  reg [63:0] _RAND_33;
  wire [40:0] _T_316; // @[Util.scala 113:33:@4728.4]
  reg [39:0] _T_318; // @[Util.scala 112:74:@4730.4]
  reg [63:0] _RAND_34;
  wire [40:0] _T_319; // @[Util.scala 113:33:@4731.4]
  reg [39:0] _T_321; // @[Util.scala 112:74:@4733.4]
  reg [63:0] _RAND_35;
  wire [40:0] _T_322; // @[Util.scala 113:33:@4734.4]
  reg [39:0] _T_324; // @[Util.scala 112:74:@4736.4]
  reg [63:0] _RAND_36;
  wire [40:0] _T_325; // @[Util.scala 113:33:@4737.4]
  reg [39:0] _T_327; // @[Util.scala 112:74:@4739.4]
  reg [63:0] _RAND_37;
  wire [40:0] _T_328; // @[Util.scala 113:33:@4740.4]
  reg [39:0] _T_330; // @[Util.scala 112:74:@4742.4]
  reg [63:0] _RAND_38;
  wire [40:0] _T_331; // @[Util.scala 113:33:@4743.4]
  reg [39:0] _T_333; // @[Util.scala 112:74:@4745.4]
  reg [63:0] _RAND_39;
  wire [40:0] _T_334; // @[Util.scala 113:33:@4746.4]
  reg [39:0] _T_336; // @[Util.scala 112:74:@4748.4]
  reg [63:0] _RAND_40;
  wire [40:0] _T_337; // @[Util.scala 113:33:@4749.4]
  reg [39:0] _T_339; // @[Util.scala 112:74:@4751.4]
  reg [63:0] _RAND_41;
  wire [40:0] _T_340; // @[Util.scala 113:33:@4752.4]
  reg [39:0] _T_342; // @[Util.scala 112:74:@4754.4]
  reg [63:0] _RAND_42;
  wire [40:0] _T_343; // @[Util.scala 113:33:@4755.4]
  reg [39:0] _T_345; // @[Util.scala 112:74:@4757.4]
  reg [63:0] _RAND_43;
  wire [40:0] _T_346; // @[Util.scala 113:33:@4758.4]
  reg [39:0] _T_348; // @[Util.scala 112:74:@4760.4]
  reg [63:0] _RAND_44;
  wire [40:0] _T_349; // @[Util.scala 113:33:@4761.4]
  reg [39:0] _T_351; // @[Util.scala 112:74:@4763.4]
  reg [63:0] _RAND_45;
  wire [40:0] _T_352; // @[Util.scala 113:33:@4764.4]
  reg [39:0] _T_354; // @[Util.scala 112:74:@4766.4]
  reg [63:0] _RAND_46;
  wire [40:0] _T_355; // @[Util.scala 113:33:@4767.4]
  reg [39:0] _T_357; // @[Util.scala 112:74:@4769.4]
  reg [63:0] _RAND_47;
  wire [40:0] _T_358; // @[Util.scala 113:33:@4770.4]
  reg [31:0] reg_dscratch; // @[CSR.scala 134:25:@4859.4]
  reg [31:0] _RAND_48;
  wire  system_insn; // @[CSR.scala 137:31:@4861.4]
  wire  _T_446; // @[CSR.scala 138:27:@4862.4]
  wire  _T_448; // @[CSR.scala 138:40:@4863.4]
  wire  cpu_ren; // @[CSR.scala 138:37:@4864.4]
  wire [31:0] read_mstatus; // @[CSR.scala 140:32:@4873.4]
  wire [15:0] _T_468; // @[CSR.scala 156:25:@4879.4]
  wire [15:0] _T_474; // @[CSR.scala 157:25:@4885.4]
  wire  _T_478; // @[CSR.scala 177:73:@4886.4]
  wire  _T_480; // @[CSR.scala 177:73:@4887.4]
  wire  _T_482; // @[CSR.scala 177:73:@4888.4]
  wire  _T_488; // @[CSR.scala 177:73:@4891.4]
  wire  _T_490; // @[CSR.scala 177:73:@4892.4]
  wire  _T_492; // @[CSR.scala 177:73:@4893.4]
  wire  _T_494; // @[CSR.scala 177:73:@4894.4]
  wire  _T_496; // @[CSR.scala 177:73:@4895.4]
  wire  _T_498; // @[CSR.scala 177:73:@4896.4]
  wire  _T_500; // @[CSR.scala 177:73:@4897.4]
  wire  _T_502; // @[CSR.scala 177:73:@4898.4]
  wire  _T_504; // @[CSR.scala 177:73:@4899.4]
  wire  _T_508; // @[CSR.scala 177:73:@4901.4]
  wire  _T_510; // @[CSR.scala 177:73:@4902.4]
  wire  _T_512; // @[CSR.scala 177:73:@4903.4]
  wire  _T_514; // @[CSR.scala 177:73:@4904.4]
  wire  _T_516; // @[CSR.scala 177:73:@4905.4]
  wire  _T_518; // @[CSR.scala 177:73:@4906.4]
  wire  _T_520; // @[CSR.scala 177:73:@4907.4]
  wire  _T_522; // @[CSR.scala 177:73:@4908.4]
  wire  _T_524; // @[CSR.scala 177:73:@4909.4]
  wire  _T_526; // @[CSR.scala 177:73:@4910.4]
  wire  _T_528; // @[CSR.scala 177:73:@4911.4]
  wire  _T_530; // @[CSR.scala 177:73:@4912.4]
  wire  _T_532; // @[CSR.scala 177:73:@4913.4]
  wire  _T_534; // @[CSR.scala 177:73:@4914.4]
  wire  _T_536; // @[CSR.scala 177:73:@4915.4]
  wire  _T_538; // @[CSR.scala 177:73:@4916.4]
  wire  _T_540; // @[CSR.scala 177:73:@4917.4]
  wire  _T_542; // @[CSR.scala 177:73:@4918.4]
  wire  _T_544; // @[CSR.scala 177:73:@4919.4]
  wire  _T_546; // @[CSR.scala 177:73:@4920.4]
  wire  _T_548; // @[CSR.scala 177:73:@4921.4]
  wire  _T_550; // @[CSR.scala 177:73:@4922.4]
  wire  _T_552; // @[CSR.scala 177:73:@4923.4]
  wire  _T_554; // @[CSR.scala 177:73:@4924.4]
  wire  _T_556; // @[CSR.scala 177:73:@4925.4]
  wire  _T_558; // @[CSR.scala 177:73:@4926.4]
  wire  _T_560; // @[CSR.scala 177:73:@4927.4]
  wire  _T_562; // @[CSR.scala 177:73:@4928.4]
  wire  _T_564; // @[CSR.scala 177:73:@4929.4]
  wire  _T_566; // @[CSR.scala 177:73:@4930.4]
  wire  _T_568; // @[CSR.scala 177:73:@4931.4]
  wire  _T_570; // @[CSR.scala 177:73:@4932.4]
  wire  _T_572; // @[CSR.scala 177:73:@4933.4]
  wire  _T_574; // @[CSR.scala 177:73:@4934.4]
  wire  _T_576; // @[CSR.scala 177:73:@4935.4]
  wire  _T_578; // @[CSR.scala 177:73:@4936.4]
  wire  _T_580; // @[CSR.scala 177:73:@4937.4]
  wire  _T_582; // @[CSR.scala 177:73:@4938.4]
  wire  _T_584; // @[CSR.scala 177:73:@4939.4]
  wire  _T_586; // @[CSR.scala 177:73:@4940.4]
  wire  _T_588; // @[CSR.scala 177:73:@4941.4]
  wire  _T_590; // @[CSR.scala 177:73:@4942.4]
  wire  _T_592; // @[CSR.scala 177:73:@4943.4]
  wire  _T_594; // @[CSR.scala 177:73:@4944.4]
  wire  _T_596; // @[CSR.scala 177:73:@4945.4]
  wire  _T_598; // @[CSR.scala 177:73:@4946.4]
  wire  _T_600; // @[CSR.scala 177:73:@4947.4]
  wire  _T_602; // @[CSR.scala 177:73:@4948.4]
  wire  _T_604; // @[CSR.scala 177:73:@4949.4]
  wire  _T_606; // @[CSR.scala 177:73:@4950.4]
  wire  _T_608; // @[CSR.scala 177:73:@4951.4]
  wire  _T_610; // @[CSR.scala 177:73:@4952.4]
  wire  _T_612; // @[CSR.scala 177:73:@4953.4]
  wire  _T_614; // @[CSR.scala 177:73:@4954.4]
  wire  _T_616; // @[CSR.scala 177:73:@4955.4]
  wire  _T_618; // @[CSR.scala 177:73:@4956.4]
  wire  _T_620; // @[CSR.scala 177:73:@4957.4]
  wire  _T_622; // @[CSR.scala 177:73:@4958.4]
  wire  _T_624; // @[CSR.scala 177:73:@4959.4]
  wire  _T_626; // @[CSR.scala 177:73:@4960.4]
  wire  _T_628; // @[CSR.scala 177:73:@4961.4]
  wire  _T_630; // @[CSR.scala 177:73:@4962.4]
  wire  _T_632; // @[CSR.scala 177:73:@4963.4]
  wire  _T_634; // @[CSR.scala 177:73:@4964.4]
  wire  _T_636; // @[CSR.scala 177:73:@4965.4]
  wire  _T_638; // @[CSR.scala 177:73:@4966.4]
  wire  _T_640; // @[CSR.scala 177:73:@4967.4]
  wire  _T_642; // @[CSR.scala 177:73:@4968.4]
  wire [1:0] _T_643; // @[CSR.scala 179:54:@4969.4]
  wire  priv_sufficient; // @[CSR.scala 179:41:@4970.4]
  wire [1:0] _T_644; // @[CSR.scala 180:29:@4971.4]
  wire [1:0] _T_645; // @[CSR.scala 180:37:@4972.4]
  wire  read_only; // @[CSR.scala 180:37:@4973.4]
  wire  _T_647; // @[CSR.scala 181:38:@4974.4]
  wire  _T_648; // @[CSR.scala 181:25:@4975.4]
  wire  cpu_wen; // @[CSR.scala 181:48:@4976.4]
  wire  _T_650; // @[CSR.scala 182:24:@4977.4]
  wire  wen; // @[CSR.scala 182:21:@4978.4]
  wire  _T_651; // @[Util.scala 23:47:@4979.4]
  wire  _T_652; // @[Util.scala 23:47:@4980.4]
  wire  _T_653; // @[Util.scala 23:62:@4981.4]
  wire [31:0] _T_655; // @[CSR.scala 281:9:@4982.4]
  wire [31:0] _T_656; // @[CSR.scala 281:49:@4983.4]
  wire [31:0] _T_659; // @[CSR.scala 281:64:@4985.4]
  wire [31:0] _T_660; // @[CSR.scala 281:60:@4986.4]
  wire [31:0] wdata; // @[CSR.scala 281:58:@4987.4]
  wire [2:0] _T_662; // @[CSR.scala 185:33:@4988.4]
  wire [7:0] opcode; // @[CSR.scala 185:20:@4989.4]
  wire  _T_663; // @[CSR.scala 186:40:@4990.4]
  wire  insn_call; // @[CSR.scala 186:31:@4991.4]
  wire  _T_664; // @[CSR.scala 187:41:@4992.4]
  wire  insn_break; // @[CSR.scala 187:32:@4993.4]
  wire  _T_665; // @[CSR.scala 188:39:@4994.4]
  wire  _T_666; // @[CSR.scala 188:30:@4995.4]
  wire  insn_ret; // @[CSR.scala 188:43:@4996.4]
  wire  _T_940; // @[CSR.scala 199:24:@5195.4]
  wire [1:0] _T_942; // @[Bitwise.scala 48:55:@5198.4]
  wire  _T_944; // @[CSR.scala 201:50:@5199.4]
  wire  _T_946; // @[CSR.scala 201:9:@5201.4]
  wire  _T_948; // @[CSR.scala 201:9:@5202.4]
  wire  _T_951; // @[CSR.scala 208:32:@5211.4]
  wire  _T_953; // @[CSR.scala 208:21:@5212.4]
  wire  _T_954; // @[CSR.scala 208:18:@5213.4]
  wire  _GEN_3; // @[CSR.scala 208:38:@5214.4]
  wire  _GEN_4; // @[CSR.scala 208:38:@5214.4]
  wire [1:0] new_prv; // @[CSR.scala 208:38:@5214.4]
  wire [3:0] _GEN_148; // @[CSR.scala 218:35:@5222.6]
  wire [4:0] _T_958; // @[CSR.scala 218:35:@5222.6]
  wire [3:0] _T_959; // @[CSR.scala 218:35:@5223.6]
  wire [31:0] _GEN_7; // @[CSR.scala 216:18:@5220.4]
  wire [31:0] _GEN_8; // @[CSR.scala 216:18:@5220.4]
  wire [31:0] _GEN_9; // @[CSR.scala 216:18:@5220.4]
  wire [31:0] _GEN_10; // @[CSR.scala 223:19:@5227.4]
  wire [31:0] _GEN_11; // @[CSR.scala 223:19:@5227.4]
  wire [31:0] _GEN_12; // @[CSR.scala 223:19:@5227.4]
  wire [31:0] _GEN_14; // @[CSR.scala 229:17:@5232.4]
  wire [31:0] _GEN_15; // @[CSR.scala 229:17:@5232.4]
  wire [31:0] _GEN_16; // @[CSR.scala 229:17:@5232.4]
  wire [63:0] _T_965; // @[Mux.scala 19:72:@5240.4]
  wire [63:0] _T_967; // @[Mux.scala 19:72:@5241.4]
  wire [15:0] _T_969; // @[Mux.scala 19:72:@5242.4]
  wire [30:0] _T_975; // @[Mux.scala 19:72:@5245.4]
  wire [31:0] _T_977; // @[Mux.scala 19:72:@5246.4]
  wire [8:0] _T_979; // @[Mux.scala 19:72:@5247.4]
  wire [15:0] _T_981; // @[Mux.scala 19:72:@5248.4]
  wire [15:0] _T_983; // @[Mux.scala 19:72:@5249.4]
  wire [31:0] _T_985; // @[Mux.scala 19:72:@5250.4]
  wire [31:0] _T_987; // @[Mux.scala 19:72:@5251.4]
  wire [31:0] _T_989; // @[Mux.scala 19:72:@5252.4]
  wire [31:0] _T_991; // @[Mux.scala 19:72:@5253.4]
  wire [31:0] _T_995; // @[Mux.scala 19:72:@5255.4]
  wire [31:0] _T_997; // @[Mux.scala 19:72:@5256.4]
  wire [39:0] _T_999; // @[Mux.scala 19:72:@5257.4]
  wire [39:0] _T_1001; // @[Mux.scala 19:72:@5258.4]
  wire [39:0] _T_1003; // @[Mux.scala 19:72:@5259.4]
  wire [39:0] _T_1005; // @[Mux.scala 19:72:@5260.4]
  wire [39:0] _T_1007; // @[Mux.scala 19:72:@5261.4]
  wire [39:0] _T_1009; // @[Mux.scala 19:72:@5262.4]
  wire [39:0] _T_1011; // @[Mux.scala 19:72:@5263.4]
  wire [39:0] _T_1013; // @[Mux.scala 19:72:@5264.4]
  wire [39:0] _T_1015; // @[Mux.scala 19:72:@5265.4]
  wire [39:0] _T_1017; // @[Mux.scala 19:72:@5266.4]
  wire [39:0] _T_1019; // @[Mux.scala 19:72:@5267.4]
  wire [39:0] _T_1021; // @[Mux.scala 19:72:@5268.4]
  wire [39:0] _T_1023; // @[Mux.scala 19:72:@5269.4]
  wire [39:0] _T_1025; // @[Mux.scala 19:72:@5270.4]
  wire [39:0] _T_1027; // @[Mux.scala 19:72:@5271.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:@5272.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:@5273.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:@5274.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:@5275.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:@5276.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:@5277.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:@5278.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:@5279.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:@5280.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:@5281.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:@5282.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:@5283.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:@5284.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:@5285.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:@5286.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:@5287.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:@5288.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:@5289.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:@5290.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:@5291.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:@5292.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:@5293.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:@5294.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:@5295.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:@5296.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:@5297.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:@5298.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:@5299.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:@5300.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:@5301.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:@5302.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:@5303.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:@5304.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:@5305.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:@5306.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:@5307.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:@5308.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:@5309.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:@5310.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:@5311.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:@5312.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:@5313.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:@5314.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:@5315.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:@5316.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:@5317.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:@5318.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:@5319.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:@5320.4]
  wire [63:0] _T_1130; // @[Mux.scala 19:72:@5323.4]
  wire [63:0] _GEN_149; // @[Mux.scala 19:72:@5324.4]
  wire [63:0] _T_1131; // @[Mux.scala 19:72:@5324.4]
  wire [63:0] _GEN_150; // @[Mux.scala 19:72:@5327.4]
  wire [63:0] _T_1134; // @[Mux.scala 19:72:@5327.4]
  wire [63:0] _GEN_151; // @[Mux.scala 19:72:@5328.4]
  wire [63:0] _T_1135; // @[Mux.scala 19:72:@5328.4]
  wire [63:0] _GEN_152; // @[Mux.scala 19:72:@5329.4]
  wire [63:0] _T_1136; // @[Mux.scala 19:72:@5329.4]
  wire [63:0] _GEN_153; // @[Mux.scala 19:72:@5330.4]
  wire [63:0] _T_1137; // @[Mux.scala 19:72:@5330.4]
  wire [63:0] _GEN_154; // @[Mux.scala 19:72:@5331.4]
  wire [63:0] _T_1138; // @[Mux.scala 19:72:@5331.4]
  wire [63:0] _GEN_155; // @[Mux.scala 19:72:@5332.4]
  wire [63:0] _T_1139; // @[Mux.scala 19:72:@5332.4]
  wire [63:0] _GEN_156; // @[Mux.scala 19:72:@5333.4]
  wire [63:0] _T_1140; // @[Mux.scala 19:72:@5333.4]
  wire [63:0] _GEN_157; // @[Mux.scala 19:72:@5334.4]
  wire [63:0] _T_1141; // @[Mux.scala 19:72:@5334.4]
  wire [63:0] _GEN_158; // @[Mux.scala 19:72:@5335.4]
  wire [63:0] _T_1142; // @[Mux.scala 19:72:@5335.4]
  wire [63:0] _GEN_159; // @[Mux.scala 19:72:@5337.4]
  wire [63:0] _T_1144; // @[Mux.scala 19:72:@5337.4]
  wire [63:0] _GEN_160; // @[Mux.scala 19:72:@5338.4]
  wire [63:0] _T_1145; // @[Mux.scala 19:72:@5338.4]
  wire [63:0] _GEN_161; // @[Mux.scala 19:72:@5339.4]
  wire [63:0] _T_1146; // @[Mux.scala 19:72:@5339.4]
  wire [63:0] _GEN_162; // @[Mux.scala 19:72:@5340.4]
  wire [63:0] _T_1147; // @[Mux.scala 19:72:@5340.4]
  wire [63:0] _GEN_163; // @[Mux.scala 19:72:@5341.4]
  wire [63:0] _T_1148; // @[Mux.scala 19:72:@5341.4]
  wire [63:0] _GEN_164; // @[Mux.scala 19:72:@5342.4]
  wire [63:0] _T_1149; // @[Mux.scala 19:72:@5342.4]
  wire [63:0] _GEN_165; // @[Mux.scala 19:72:@5343.4]
  wire [63:0] _T_1150; // @[Mux.scala 19:72:@5343.4]
  wire [63:0] _GEN_166; // @[Mux.scala 19:72:@5344.4]
  wire [63:0] _T_1151; // @[Mux.scala 19:72:@5344.4]
  wire [63:0] _GEN_167; // @[Mux.scala 19:72:@5345.4]
  wire [63:0] _T_1152; // @[Mux.scala 19:72:@5345.4]
  wire [63:0] _GEN_168; // @[Mux.scala 19:72:@5346.4]
  wire [63:0] _T_1153; // @[Mux.scala 19:72:@5346.4]
  wire [63:0] _GEN_169; // @[Mux.scala 19:72:@5347.4]
  wire [63:0] _T_1154; // @[Mux.scala 19:72:@5347.4]
  wire [63:0] _GEN_170; // @[Mux.scala 19:72:@5348.4]
  wire [63:0] _T_1155; // @[Mux.scala 19:72:@5348.4]
  wire [63:0] _GEN_171; // @[Mux.scala 19:72:@5349.4]
  wire [63:0] _T_1156; // @[Mux.scala 19:72:@5349.4]
  wire [63:0] _GEN_172; // @[Mux.scala 19:72:@5350.4]
  wire [63:0] _T_1157; // @[Mux.scala 19:72:@5350.4]
  wire [63:0] _GEN_173; // @[Mux.scala 19:72:@5351.4]
  wire [63:0] _T_1158; // @[Mux.scala 19:72:@5351.4]
  wire [63:0] _GEN_174; // @[Mux.scala 19:72:@5352.4]
  wire [63:0] _T_1159; // @[Mux.scala 19:72:@5352.4]
  wire [63:0] _GEN_175; // @[Mux.scala 19:72:@5353.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:@5353.4]
  wire [63:0] _GEN_176; // @[Mux.scala 19:72:@5354.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:@5354.4]
  wire [63:0] _GEN_177; // @[Mux.scala 19:72:@5355.4]
  wire [63:0] _T_1162; // @[Mux.scala 19:72:@5355.4]
  wire [63:0] _GEN_178; // @[Mux.scala 19:72:@5356.4]
  wire [63:0] _T_1163; // @[Mux.scala 19:72:@5356.4]
  wire [63:0] _GEN_179; // @[Mux.scala 19:72:@5357.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:@5357.4]
  wire [63:0] _GEN_180; // @[Mux.scala 19:72:@5358.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:@5358.4]
  wire [63:0] _GEN_181; // @[Mux.scala 19:72:@5359.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:@5359.4]
  wire [63:0] _GEN_182; // @[Mux.scala 19:72:@5360.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:@5360.4]
  wire [63:0] _GEN_183; // @[Mux.scala 19:72:@5361.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:@5361.4]
  wire [63:0] _GEN_184; // @[Mux.scala 19:72:@5362.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:@5362.4]
  wire [63:0] _GEN_185; // @[Mux.scala 19:72:@5363.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:@5363.4]
  wire [63:0] _GEN_186; // @[Mux.scala 19:72:@5364.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:@5364.4]
  wire [63:0] _GEN_187; // @[Mux.scala 19:72:@5365.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:@5365.4]
  wire [63:0] _GEN_188; // @[Mux.scala 19:72:@5366.4]
  wire [63:0] _T_1173; // @[Mux.scala 19:72:@5366.4]
  wire [63:0] _GEN_189; // @[Mux.scala 19:72:@5367.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:@5367.4]
  wire [63:0] _GEN_190; // @[Mux.scala 19:72:@5368.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:@5368.4]
  wire [63:0] _GEN_191; // @[Mux.scala 19:72:@5369.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:@5369.4]
  wire [63:0] _GEN_192; // @[Mux.scala 19:72:@5370.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:@5370.4]
  wire [63:0] _GEN_193; // @[Mux.scala 19:72:@5371.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:@5371.4]
  wire [63:0] _GEN_194; // @[Mux.scala 19:72:@5372.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:@5372.4]
  wire [63:0] _GEN_195; // @[Mux.scala 19:72:@5373.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:@5373.4]
  wire [63:0] _GEN_196; // @[Mux.scala 19:72:@5374.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:@5374.4]
  wire [63:0] _GEN_197; // @[Mux.scala 19:72:@5375.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:@5375.4]
  wire [63:0] _GEN_198; // @[Mux.scala 19:72:@5376.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:@5376.4]
  wire [63:0] _GEN_199; // @[Mux.scala 19:72:@5377.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:@5377.4]
  wire [63:0] _GEN_200; // @[Mux.scala 19:72:@5378.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:@5378.4]
  wire [63:0] _GEN_201; // @[Mux.scala 19:72:@5379.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:@5379.4]
  wire [63:0] _GEN_202; // @[Mux.scala 19:72:@5380.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:@5380.4]
  wire [63:0] _GEN_203; // @[Mux.scala 19:72:@5381.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:@5381.4]
  wire [63:0] _GEN_204; // @[Mux.scala 19:72:@5382.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:@5382.4]
  wire [63:0] _GEN_205; // @[Mux.scala 19:72:@5383.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:@5383.4]
  wire [63:0] _GEN_206; // @[Mux.scala 19:72:@5384.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:@5384.4]
  wire [63:0] _GEN_207; // @[Mux.scala 19:72:@5385.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:@5385.4]
  wire [63:0] _GEN_208; // @[Mux.scala 19:72:@5386.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:@5386.4]
  wire [63:0] _GEN_209; // @[Mux.scala 19:72:@5387.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:@5387.4]
  wire [63:0] _GEN_210; // @[Mux.scala 19:72:@5388.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:@5388.4]
  wire [63:0] _GEN_211; // @[Mux.scala 19:72:@5389.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:@5389.4]
  wire [63:0] _GEN_212; // @[Mux.scala 19:72:@5390.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:@5390.4]
  wire [63:0] _GEN_213; // @[Mux.scala 19:72:@5391.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:@5391.4]
  wire [63:0] _GEN_214; // @[Mux.scala 19:72:@5392.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:@5392.4]
  wire [63:0] _GEN_215; // @[Mux.scala 19:72:@5393.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:@5393.4]
  wire [63:0] _GEN_216; // @[Mux.scala 19:72:@5394.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:@5394.4]
  wire [63:0] _GEN_217; // @[Mux.scala 19:72:@5395.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:@5395.4]
  wire [63:0] _GEN_218; // @[Mux.scala 19:72:@5396.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:@5396.4]
  wire [63:0] _GEN_219; // @[Mux.scala 19:72:@5397.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:@5397.4]
  wire [63:0] _GEN_220; // @[Mux.scala 19:72:@5398.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:@5398.4]
  wire [63:0] _GEN_221; // @[Mux.scala 19:72:@5399.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:@5399.4]
  wire [63:0] _GEN_222; // @[Mux.scala 19:72:@5400.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:@5400.4]
  wire [63:0] _GEN_223; // @[Mux.scala 19:72:@5401.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:@5401.4]
  wire [63:0] _GEN_224; // @[Mux.scala 19:72:@5402.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:@5402.4]
  wire  _T_1220; // @[CSR.scala 245:39:@5415.8]
  wire  _T_1222; // @[CSR.scala 245:39:@5419.8]
  wire  _GEN_17; // @[CSR.scala 244:39:@5409.6]
  wire  _GEN_18; // @[CSR.scala 244:39:@5409.6]
  wire [15:0] _T_1233; // @[:@5438.8 :@5439.8]
  wire  _T_1235; // @[CSR.scala 250:35:@5442.8]
  wire  _T_1237; // @[CSR.scala 250:35:@5446.8]
  wire  _GEN_19; // @[CSR.scala 249:35:@5436.6]
  wire  _GEN_20; // @[CSR.scala 253:35:@5456.6]
  wire  _GEN_21; // @[CSR.scala 253:35:@5456.6]
  wire [7:0] _T_1253; // @[CSR.scala 277:47:@5478.8]
  wire [31:0] _T_1254; // @[CSR.scala 277:72:@5479.8]
  wire [39:0] _T_1255; // @[Cat.scala 30:58:@5480.8]
  wire [40:0] _GEN_22; // @[CSR.scala 277:29:@5477.6]
  wire [7:0] _T_1256; // @[CSR.scala 278:45:@5484.8]
  wire [39:0] _T_1257; // @[Cat.scala 30:58:@5485.8]
  wire [40:0] _GEN_23; // @[CSR.scala 278:29:@5483.6]
  wire [31:0] _T_1259; // @[CSR.scala 277:72:@5490.8]
  wire [39:0] _T_1260; // @[Cat.scala 30:58:@5491.8]
  wire [40:0] _GEN_24; // @[CSR.scala 277:29:@5488.6]
  wire [7:0] _T_1261; // @[CSR.scala 278:45:@5495.8]
  wire [39:0] _T_1262; // @[Cat.scala 30:58:@5496.8]
  wire [40:0] _GEN_25; // @[CSR.scala 278:29:@5494.6]
  wire [31:0] _T_1264; // @[CSR.scala 277:72:@5501.8]
  wire [39:0] _T_1265; // @[Cat.scala 30:58:@5502.8]
  wire [40:0] _GEN_26; // @[CSR.scala 277:29:@5499.6]
  wire [7:0] _T_1266; // @[CSR.scala 278:45:@5506.8]
  wire [39:0] _T_1267; // @[Cat.scala 30:58:@5507.8]
  wire [40:0] _GEN_27; // @[CSR.scala 278:29:@5505.6]
  wire [31:0] _T_1269; // @[CSR.scala 277:72:@5512.8]
  wire [39:0] _T_1270; // @[Cat.scala 30:58:@5513.8]
  wire [40:0] _GEN_28; // @[CSR.scala 277:29:@5510.6]
  wire [7:0] _T_1271; // @[CSR.scala 278:45:@5517.8]
  wire [39:0] _T_1272; // @[Cat.scala 30:58:@5518.8]
  wire [40:0] _GEN_29; // @[CSR.scala 278:29:@5516.6]
  wire [31:0] _T_1274; // @[CSR.scala 277:72:@5523.8]
  wire [39:0] _T_1275; // @[Cat.scala 30:58:@5524.8]
  wire [40:0] _GEN_30; // @[CSR.scala 277:29:@5521.6]
  wire [7:0] _T_1276; // @[CSR.scala 278:45:@5528.8]
  wire [39:0] _T_1277; // @[Cat.scala 30:58:@5529.8]
  wire [40:0] _GEN_31; // @[CSR.scala 278:29:@5527.6]
  wire [31:0] _T_1279; // @[CSR.scala 277:72:@5534.8]
  wire [39:0] _T_1280; // @[Cat.scala 30:58:@5535.8]
  wire [40:0] _GEN_32; // @[CSR.scala 277:29:@5532.6]
  wire [7:0] _T_1281; // @[CSR.scala 278:45:@5539.8]
  wire [39:0] _T_1282; // @[Cat.scala 30:58:@5540.8]
  wire [40:0] _GEN_33; // @[CSR.scala 278:29:@5538.6]
  wire [31:0] _T_1284; // @[CSR.scala 277:72:@5545.8]
  wire [39:0] _T_1285; // @[Cat.scala 30:58:@5546.8]
  wire [40:0] _GEN_34; // @[CSR.scala 277:29:@5543.6]
  wire [7:0] _T_1286; // @[CSR.scala 278:45:@5550.8]
  wire [39:0] _T_1287; // @[Cat.scala 30:58:@5551.8]
  wire [40:0] _GEN_35; // @[CSR.scala 278:29:@5549.6]
  wire [31:0] _T_1289; // @[CSR.scala 277:72:@5556.8]
  wire [39:0] _T_1290; // @[Cat.scala 30:58:@5557.8]
  wire [40:0] _GEN_36; // @[CSR.scala 277:29:@5554.6]
  wire [7:0] _T_1291; // @[CSR.scala 278:45:@5561.8]
  wire [39:0] _T_1292; // @[Cat.scala 30:58:@5562.8]
  wire [40:0] _GEN_37; // @[CSR.scala 278:29:@5560.6]
  wire [31:0] _T_1294; // @[CSR.scala 277:72:@5567.8]
  wire [39:0] _T_1295; // @[Cat.scala 30:58:@5568.8]
  wire [40:0] _GEN_38; // @[CSR.scala 277:29:@5565.6]
  wire [7:0] _T_1296; // @[CSR.scala 278:45:@5572.8]
  wire [39:0] _T_1297; // @[Cat.scala 30:58:@5573.8]
  wire [40:0] _GEN_39; // @[CSR.scala 278:29:@5571.6]
  wire [31:0] _T_1299; // @[CSR.scala 277:72:@5578.8]
  wire [39:0] _T_1300; // @[Cat.scala 30:58:@5579.8]
  wire [40:0] _GEN_40; // @[CSR.scala 277:29:@5576.6]
  wire [7:0] _T_1301; // @[CSR.scala 278:45:@5583.8]
  wire [39:0] _T_1302; // @[Cat.scala 30:58:@5584.8]
  wire [40:0] _GEN_41; // @[CSR.scala 278:29:@5582.6]
  wire [31:0] _T_1304; // @[CSR.scala 277:72:@5589.8]
  wire [39:0] _T_1305; // @[Cat.scala 30:58:@5590.8]
  wire [40:0] _GEN_42; // @[CSR.scala 277:29:@5587.6]
  wire [7:0] _T_1306; // @[CSR.scala 278:45:@5594.8]
  wire [39:0] _T_1307; // @[Cat.scala 30:58:@5595.8]
  wire [40:0] _GEN_43; // @[CSR.scala 278:29:@5593.6]
  wire [31:0] _T_1309; // @[CSR.scala 277:72:@5600.8]
  wire [39:0] _T_1310; // @[Cat.scala 30:58:@5601.8]
  wire [40:0] _GEN_44; // @[CSR.scala 277:29:@5598.6]
  wire [7:0] _T_1311; // @[CSR.scala 278:45:@5605.8]
  wire [39:0] _T_1312; // @[Cat.scala 30:58:@5606.8]
  wire [40:0] _GEN_45; // @[CSR.scala 278:29:@5604.6]
  wire [31:0] _T_1314; // @[CSR.scala 277:72:@5611.8]
  wire [39:0] _T_1315; // @[Cat.scala 30:58:@5612.8]
  wire [40:0] _GEN_46; // @[CSR.scala 277:29:@5609.6]
  wire [7:0] _T_1316; // @[CSR.scala 278:45:@5616.8]
  wire [39:0] _T_1317; // @[Cat.scala 30:58:@5617.8]
  wire [40:0] _GEN_47; // @[CSR.scala 278:29:@5615.6]
  wire [31:0] _T_1319; // @[CSR.scala 277:72:@5622.8]
  wire [39:0] _T_1320; // @[Cat.scala 30:58:@5623.8]
  wire [40:0] _GEN_48; // @[CSR.scala 277:29:@5620.6]
  wire [7:0] _T_1321; // @[CSR.scala 278:45:@5627.8]
  wire [39:0] _T_1322; // @[Cat.scala 30:58:@5628.8]
  wire [40:0] _GEN_49; // @[CSR.scala 278:29:@5626.6]
  wire [31:0] _T_1324; // @[CSR.scala 277:72:@5633.8]
  wire [39:0] _T_1325; // @[Cat.scala 30:58:@5634.8]
  wire [40:0] _GEN_50; // @[CSR.scala 277:29:@5631.6]
  wire [7:0] _T_1326; // @[CSR.scala 278:45:@5638.8]
  wire [39:0] _T_1327; // @[Cat.scala 30:58:@5639.8]
  wire [40:0] _GEN_51; // @[CSR.scala 278:29:@5637.6]
  wire [31:0] _T_1329; // @[CSR.scala 277:72:@5644.8]
  wire [39:0] _T_1330; // @[Cat.scala 30:58:@5645.8]
  wire [40:0] _GEN_52; // @[CSR.scala 277:29:@5642.6]
  wire [7:0] _T_1331; // @[CSR.scala 278:45:@5649.8]
  wire [39:0] _T_1332; // @[Cat.scala 30:58:@5650.8]
  wire [40:0] _GEN_53; // @[CSR.scala 278:29:@5648.6]
  wire [31:0] _T_1334; // @[CSR.scala 277:72:@5655.8]
  wire [39:0] _T_1335; // @[Cat.scala 30:58:@5656.8]
  wire [40:0] _GEN_54; // @[CSR.scala 277:29:@5653.6]
  wire [7:0] _T_1336; // @[CSR.scala 278:45:@5660.8]
  wire [39:0] _T_1337; // @[Cat.scala 30:58:@5661.8]
  wire [40:0] _GEN_55; // @[CSR.scala 278:29:@5659.6]
  wire [31:0] _T_1339; // @[CSR.scala 277:72:@5666.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:@5667.8]
  wire [40:0] _GEN_56; // @[CSR.scala 277:29:@5664.6]
  wire [7:0] _T_1341; // @[CSR.scala 278:45:@5671.8]
  wire [39:0] _T_1342; // @[Cat.scala 30:58:@5672.8]
  wire [40:0] _GEN_57; // @[CSR.scala 278:29:@5670.6]
  wire [31:0] _T_1344; // @[CSR.scala 277:72:@5677.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:@5678.8]
  wire [40:0] _GEN_58; // @[CSR.scala 277:29:@5675.6]
  wire [7:0] _T_1346; // @[CSR.scala 278:45:@5682.8]
  wire [39:0] _T_1347; // @[Cat.scala 30:58:@5683.8]
  wire [40:0] _GEN_59; // @[CSR.scala 278:29:@5681.6]
  wire [31:0] _T_1349; // @[CSR.scala 277:72:@5688.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:@5689.8]
  wire [40:0] _GEN_60; // @[CSR.scala 277:29:@5686.6]
  wire [7:0] _T_1351; // @[CSR.scala 278:45:@5693.8]
  wire [39:0] _T_1352; // @[Cat.scala 30:58:@5694.8]
  wire [40:0] _GEN_61; // @[CSR.scala 278:29:@5692.6]
  wire [31:0] _T_1354; // @[CSR.scala 277:72:@5699.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:@5700.8]
  wire [40:0] _GEN_62; // @[CSR.scala 277:29:@5697.6]
  wire [7:0] _T_1356; // @[CSR.scala 278:45:@5704.8]
  wire [39:0] _T_1357; // @[Cat.scala 30:58:@5705.8]
  wire [40:0] _GEN_63; // @[CSR.scala 278:29:@5703.6]
  wire [31:0] _T_1359; // @[CSR.scala 277:72:@5710.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:@5711.8]
  wire [40:0] _GEN_64; // @[CSR.scala 277:29:@5708.6]
  wire [7:0] _T_1361; // @[CSR.scala 278:45:@5715.8]
  wire [39:0] _T_1362; // @[Cat.scala 30:58:@5716.8]
  wire [40:0] _GEN_65; // @[CSR.scala 278:29:@5714.6]
  wire [31:0] _T_1364; // @[CSR.scala 277:72:@5721.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:@5722.8]
  wire [40:0] _GEN_66; // @[CSR.scala 277:29:@5719.6]
  wire [7:0] _T_1366; // @[CSR.scala 278:45:@5726.8]
  wire [39:0] _T_1367; // @[Cat.scala 30:58:@5727.8]
  wire [40:0] _GEN_67; // @[CSR.scala 278:29:@5725.6]
  wire [31:0] _T_1369; // @[CSR.scala 277:72:@5732.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:@5733.8]
  wire [40:0] _GEN_68; // @[CSR.scala 277:29:@5730.6]
  wire [7:0] _T_1371; // @[CSR.scala 278:45:@5737.8]
  wire [39:0] _T_1372; // @[Cat.scala 30:58:@5738.8]
  wire [40:0] _GEN_69; // @[CSR.scala 278:29:@5736.6]
  wire [31:0] _T_1374; // @[CSR.scala 277:72:@5743.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:@5744.8]
  wire [40:0] _GEN_70; // @[CSR.scala 277:29:@5741.6]
  wire [7:0] _T_1376; // @[CSR.scala 278:45:@5748.8]
  wire [39:0] _T_1377; // @[Cat.scala 30:58:@5749.8]
  wire [40:0] _GEN_71; // @[CSR.scala 278:29:@5747.6]
  wire [31:0] _T_1379; // @[CSR.scala 277:72:@5754.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:@5755.8]
  wire [40:0] _GEN_72; // @[CSR.scala 277:29:@5752.6]
  wire [7:0] _T_1381; // @[CSR.scala 278:45:@5759.8]
  wire [39:0] _T_1382; // @[Cat.scala 30:58:@5760.8]
  wire [40:0] _GEN_73; // @[CSR.scala 278:29:@5758.6]
  wire [31:0] _T_1384; // @[CSR.scala 277:72:@5765.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:@5766.8]
  wire [40:0] _GEN_74; // @[CSR.scala 277:29:@5763.6]
  wire [7:0] _T_1386; // @[CSR.scala 278:45:@5770.8]
  wire [39:0] _T_1387; // @[Cat.scala 30:58:@5771.8]
  wire [40:0] _GEN_75; // @[CSR.scala 278:29:@5769.6]
  wire [31:0] _T_1389; // @[CSR.scala 277:72:@5776.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:@5777.8]
  wire [40:0] _GEN_76; // @[CSR.scala 277:29:@5774.6]
  wire [7:0] _T_1391; // @[CSR.scala 278:45:@5781.8]
  wire [39:0] _T_1392; // @[Cat.scala 30:58:@5782.8]
  wire [40:0] _GEN_77; // @[CSR.scala 278:29:@5780.6]
  wire [31:0] _T_1394; // @[CSR.scala 277:72:@5787.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:@5788.8]
  wire [40:0] _GEN_78; // @[CSR.scala 277:29:@5785.6]
  wire [7:0] _T_1396; // @[CSR.scala 278:45:@5792.8]
  wire [39:0] _T_1397; // @[Cat.scala 30:58:@5793.8]
  wire [40:0] _GEN_79; // @[CSR.scala 278:29:@5791.6]
  wire [31:0] _T_1399; // @[CSR.scala 277:72:@5798.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:@5799.8]
  wire [40:0] _GEN_80; // @[CSR.scala 277:29:@5796.6]
  wire [7:0] _T_1401; // @[CSR.scala 278:45:@5803.8]
  wire [39:0] _T_1402; // @[Cat.scala 30:58:@5804.8]
  wire [40:0] _GEN_81; // @[CSR.scala 278:29:@5802.6]
  wire [31:0] _T_1404; // @[CSR.scala 277:72:@5809.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:@5810.8]
  wire [40:0] _GEN_82; // @[CSR.scala 277:29:@5807.6]
  wire [7:0] _T_1406; // @[CSR.scala 278:45:@5814.8]
  wire [39:0] _T_1407; // @[Cat.scala 30:58:@5815.8]
  wire [40:0] _GEN_83; // @[CSR.scala 278:29:@5813.6]
  wire [31:0] _T_1409; // @[CSR.scala 277:72:@5820.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:@5821.8]
  wire [40:0] _GEN_84; // @[CSR.scala 277:29:@5818.6]
  wire [7:0] _T_1411; // @[CSR.scala 278:45:@5825.8]
  wire [39:0] _T_1412; // @[Cat.scala 30:58:@5826.8]
  wire [40:0] _GEN_85; // @[CSR.scala 278:29:@5824.6]
  wire [31:0] _T_1414; // @[CSR.scala 277:72:@5831.8]
  wire [63:0] _T_1415; // @[Cat.scala 30:58:@5832.8]
  wire [57:0] _T_1416; // @[Util.scala 133:28:@5834.8]
  wire [63:0] _GEN_86; // @[CSR.scala 277:29:@5829.6]
  wire [57:0] _GEN_87; // @[CSR.scala 277:29:@5829.6]
  wire [31:0] _T_1417; // @[CSR.scala 278:45:@5838.8]
  wire [63:0] _T_1418; // @[Cat.scala 30:58:@5839.8]
  wire [57:0] _T_1419; // @[Util.scala 133:28:@5841.8]
  wire [63:0] _GEN_88; // @[CSR.scala 278:29:@5837.6]
  wire [57:0] _GEN_89; // @[CSR.scala 278:29:@5837.6]
  wire [31:0] _T_1421; // @[CSR.scala 277:72:@5846.8]
  wire [63:0] _T_1422; // @[Cat.scala 30:58:@5847.8]
  wire [57:0] _T_1423; // @[Util.scala 133:28:@5849.8]
  wire [63:0] _GEN_90; // @[CSR.scala 277:29:@5844.6]
  wire [57:0] _GEN_91; // @[CSR.scala 277:29:@5844.6]
  wire [31:0] _T_1424; // @[CSR.scala 278:45:@5853.8]
  wire [63:0] _T_1425; // @[Cat.scala 30:58:@5854.8]
  wire [57:0] _T_1426; // @[Util.scala 133:28:@5856.8]
  wire [63:0] _GEN_92; // @[CSR.scala 278:29:@5852.6]
  wire [57:0] _GEN_93; // @[CSR.scala 278:29:@5852.6]
  wire [31:0] _GEN_94; // @[CSR.scala 265:40:@5859.6]
  wire [31:0] _T_1429; // @[CSR.scala 267:78:@5864.8]
  wire [34:0] _GEN_225; // @[CSR.scala 267:86:@5865.8]
  wire [34:0] _T_1431; // @[CSR.scala 267:86:@5865.8]
  wire [34:0] _GEN_95; // @[CSR.scala 267:40:@5862.6]
  wire [31:0] _GEN_96; // @[CSR.scala 268:40:@5868.6]
  wire [31:0] _T_1433; // @[CSR.scala 269:62:@5872.8]
  wire [31:0] _GEN_97; // @[CSR.scala 269:40:@5871.6]
  wire [31:0] _GEN_98; // @[CSR.scala 270:40:@5875.6]
  wire [31:0] _GEN_99; // @[CSR.scala 271:42:@5879.6]
  wire  _GEN_100; // @[CSR.scala 242:14:@5408.4]
  wire  _GEN_101; // @[CSR.scala 242:14:@5408.4]
  wire  _GEN_102; // @[CSR.scala 242:14:@5408.4]
  wire  _GEN_103; // @[CSR.scala 242:14:@5408.4]
  wire  _GEN_104; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_105; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_106; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_107; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_108; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_109; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_110; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_111; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_112; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_113; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_114; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_115; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_116; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_117; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_118; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_119; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_120; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_121; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_122; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_123; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_124; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_125; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_126; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_127; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_128; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_129; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_130; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_131; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_132; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_133; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_134; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_135; // @[CSR.scala 242:14:@5408.4]
  wire [40:0] _GEN_136; // @[CSR.scala 242:14:@5408.4]
  wire [63:0] _GEN_137; // @[CSR.scala 242:14:@5408.4]
  wire [57:0] _GEN_138; // @[CSR.scala 242:14:@5408.4]
  wire [63:0] _GEN_139; // @[CSR.scala 242:14:@5408.4]
  wire [57:0] _GEN_140; // @[CSR.scala 242:14:@5408.4]
  wire [34:0] _GEN_142; // @[CSR.scala 242:14:@5408.4]
  assign _T_241 = _T_240 + 6'h1; // @[Util.scala 113:33:@4654.4]
  assign _T_245 = _T_241[6]; // @[Util.scala 118:20:@4657.4]
  assign _T_247 = _T_244 + 58'h1; // @[Util.scala 118:43:@4659.6]
  assign _T_248 = _T_244 + 58'h1; // @[Util.scala 118:43:@4660.6]
  assign _GEN_0 = _T_245 ? _T_248 : _T_244; // @[Util.scala 118:34:@4658.4]
  assign _T_249 = {_T_244,_T_240}; // @[Cat.scala 30:58:@4663.4]
  assign _GEN_147 = {{4'd0}, io_retire}; // @[Util.scala 113:33:@4665.4]
  assign _T_253 = _T_252 + _GEN_147; // @[Util.scala 113:33:@4665.4]
  assign _T_257 = _T_253[6]; // @[Util.scala 118:20:@4668.4]
  assign _T_259 = _T_256 + 58'h1; // @[Util.scala 118:43:@4670.6]
  assign _T_260 = _T_256 + 58'h1; // @[Util.scala 118:43:@4671.6]
  assign _GEN_1 = _T_257 ? _T_260 : _T_256; // @[Util.scala 118:34:@4669.4]
  assign _T_261 = {_T_256,_T_252}; // @[Cat.scala 30:58:@4674.4]
  assign _T_265 = {{1'd0}, _T_264}; // @[Util.scala 113:33:@4677.4]
  assign _T_268 = {{1'd0}, _T_267}; // @[Util.scala 113:33:@4680.4]
  assign _T_271 = {{1'd0}, _T_270}; // @[Util.scala 113:33:@4683.4]
  assign _T_274 = {{1'd0}, _T_273}; // @[Util.scala 113:33:@4686.4]
  assign _T_277 = {{1'd0}, _T_276}; // @[Util.scala 113:33:@4689.4]
  assign _T_280 = {{1'd0}, _T_279}; // @[Util.scala 113:33:@4692.4]
  assign _T_283 = {{1'd0}, _T_282}; // @[Util.scala 113:33:@4695.4]
  assign _T_286 = {{1'd0}, _T_285}; // @[Util.scala 113:33:@4698.4]
  assign _T_289 = {{1'd0}, _T_288}; // @[Util.scala 113:33:@4701.4]
  assign _T_292 = {{1'd0}, _T_291}; // @[Util.scala 113:33:@4704.4]
  assign _T_295 = {{1'd0}, _T_294}; // @[Util.scala 113:33:@4707.4]
  assign _T_298 = {{1'd0}, _T_297}; // @[Util.scala 113:33:@4710.4]
  assign _T_301 = {{1'd0}, _T_300}; // @[Util.scala 113:33:@4713.4]
  assign _T_304 = {{1'd0}, _T_303}; // @[Util.scala 113:33:@4716.4]
  assign _T_307 = {{1'd0}, _T_306}; // @[Util.scala 113:33:@4719.4]
  assign _T_310 = {{1'd0}, _T_309}; // @[Util.scala 113:33:@4722.4]
  assign _T_313 = {{1'd0}, _T_312}; // @[Util.scala 113:33:@4725.4]
  assign _T_316 = {{1'd0}, _T_315}; // @[Util.scala 113:33:@4728.4]
  assign _T_319 = {{1'd0}, _T_318}; // @[Util.scala 113:33:@4731.4]
  assign _T_322 = {{1'd0}, _T_321}; // @[Util.scala 113:33:@4734.4]
  assign _T_325 = {{1'd0}, _T_324}; // @[Util.scala 113:33:@4737.4]
  assign _T_328 = {{1'd0}, _T_327}; // @[Util.scala 113:33:@4740.4]
  assign _T_331 = {{1'd0}, _T_330}; // @[Util.scala 113:33:@4743.4]
  assign _T_334 = {{1'd0}, _T_333}; // @[Util.scala 113:33:@4746.4]
  assign _T_337 = {{1'd0}, _T_336}; // @[Util.scala 113:33:@4749.4]
  assign _T_340 = {{1'd0}, _T_339}; // @[Util.scala 113:33:@4752.4]
  assign _T_343 = {{1'd0}, _T_342}; // @[Util.scala 113:33:@4755.4]
  assign _T_346 = {{1'd0}, _T_345}; // @[Util.scala 113:33:@4758.4]
  assign _T_349 = {{1'd0}, _T_348}; // @[Util.scala 113:33:@4761.4]
  assign _T_352 = {{1'd0}, _T_351}; // @[Util.scala 113:33:@4764.4]
  assign _T_355 = {{1'd0}, _T_354}; // @[Util.scala 113:33:@4767.4]
  assign _T_358 = {{1'd0}, _T_357}; // @[Util.scala 113:33:@4770.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 137:31:@4861.4]
  assign _T_446 = io_rw_cmd != 3'h0; // @[CSR.scala 138:27:@4862.4]
  assign _T_448 = system_insn == 1'h0; // @[CSR.scala 138:40:@4863.4]
  assign cpu_ren = _T_446 & _T_448; // @[CSR.scala 138:37:@4864.4]
  assign read_mstatus = {io_status_prv,io_status_unimp5,io_status_mprv,io_status_unimp4,io_status_mpp,io_status_unimp3,io_status_mpie,io_status_unimp2,io_status_mie,io_status_unimp1}; // @[CSR.scala 140:32:@4873.4]
  assign _T_468 = {5'h0,3'h0,reg_mip_mtip,3'h0,reg_mip_msip,3'h0}; // @[CSR.scala 156:25:@4879.4]
  assign _T_474 = {5'h0,3'h0,reg_mie_mtip,3'h0,reg_mie_msip,3'h0}; // @[CSR.scala 157:25:@4885.4]
  assign _T_478 = io_rw_addr == 12'hb00; // @[CSR.scala 177:73:@4886.4]
  assign _T_480 = io_rw_addr == 12'hb02; // @[CSR.scala 177:73:@4887.4]
  assign _T_482 = io_rw_addr == 12'hf13; // @[CSR.scala 177:73:@4888.4]
  assign _T_488 = io_rw_addr == 12'h301; // @[CSR.scala 177:73:@4891.4]
  assign _T_490 = io_rw_addr == 12'h300; // @[CSR.scala 177:73:@4892.4]
  assign _T_492 = io_rw_addr == 12'h305; // @[CSR.scala 177:73:@4893.4]
  assign _T_494 = io_rw_addr == 12'h344; // @[CSR.scala 177:73:@4894.4]
  assign _T_496 = io_rw_addr == 12'h304; // @[CSR.scala 177:73:@4895.4]
  assign _T_498 = io_rw_addr == 12'h340; // @[CSR.scala 177:73:@4896.4]
  assign _T_500 = io_rw_addr == 12'h341; // @[CSR.scala 177:73:@4897.4]
  assign _T_502 = io_rw_addr == 12'h343; // @[CSR.scala 177:73:@4898.4]
  assign _T_504 = io_rw_addr == 12'h342; // @[CSR.scala 177:73:@4899.4]
  assign _T_508 = io_rw_addr == 12'h7b2; // @[CSR.scala 177:73:@4901.4]
  assign _T_510 = io_rw_addr == 12'h302; // @[CSR.scala 177:73:@4902.4]
  assign _T_512 = io_rw_addr == 12'hb03; // @[CSR.scala 177:73:@4903.4]
  assign _T_514 = io_rw_addr == 12'hb83; // @[CSR.scala 177:73:@4904.4]
  assign _T_516 = io_rw_addr == 12'hb04; // @[CSR.scala 177:73:@4905.4]
  assign _T_518 = io_rw_addr == 12'hb84; // @[CSR.scala 177:73:@4906.4]
  assign _T_520 = io_rw_addr == 12'hb05; // @[CSR.scala 177:73:@4907.4]
  assign _T_522 = io_rw_addr == 12'hb85; // @[CSR.scala 177:73:@4908.4]
  assign _T_524 = io_rw_addr == 12'hb06; // @[CSR.scala 177:73:@4909.4]
  assign _T_526 = io_rw_addr == 12'hb86; // @[CSR.scala 177:73:@4910.4]
  assign _T_528 = io_rw_addr == 12'hb07; // @[CSR.scala 177:73:@4911.4]
  assign _T_530 = io_rw_addr == 12'hb87; // @[CSR.scala 177:73:@4912.4]
  assign _T_532 = io_rw_addr == 12'hb08; // @[CSR.scala 177:73:@4913.4]
  assign _T_534 = io_rw_addr == 12'hb88; // @[CSR.scala 177:73:@4914.4]
  assign _T_536 = io_rw_addr == 12'hb09; // @[CSR.scala 177:73:@4915.4]
  assign _T_538 = io_rw_addr == 12'hb89; // @[CSR.scala 177:73:@4916.4]
  assign _T_540 = io_rw_addr == 12'hb0a; // @[CSR.scala 177:73:@4917.4]
  assign _T_542 = io_rw_addr == 12'hb8a; // @[CSR.scala 177:73:@4918.4]
  assign _T_544 = io_rw_addr == 12'hb0b; // @[CSR.scala 177:73:@4919.4]
  assign _T_546 = io_rw_addr == 12'hb8b; // @[CSR.scala 177:73:@4920.4]
  assign _T_548 = io_rw_addr == 12'hb0c; // @[CSR.scala 177:73:@4921.4]
  assign _T_550 = io_rw_addr == 12'hb8c; // @[CSR.scala 177:73:@4922.4]
  assign _T_552 = io_rw_addr == 12'hb0d; // @[CSR.scala 177:73:@4923.4]
  assign _T_554 = io_rw_addr == 12'hb8d; // @[CSR.scala 177:73:@4924.4]
  assign _T_556 = io_rw_addr == 12'hb0e; // @[CSR.scala 177:73:@4925.4]
  assign _T_558 = io_rw_addr == 12'hb8e; // @[CSR.scala 177:73:@4926.4]
  assign _T_560 = io_rw_addr == 12'hb0f; // @[CSR.scala 177:73:@4927.4]
  assign _T_562 = io_rw_addr == 12'hb8f; // @[CSR.scala 177:73:@4928.4]
  assign _T_564 = io_rw_addr == 12'hb10; // @[CSR.scala 177:73:@4929.4]
  assign _T_566 = io_rw_addr == 12'hb90; // @[CSR.scala 177:73:@4930.4]
  assign _T_568 = io_rw_addr == 12'hb11; // @[CSR.scala 177:73:@4931.4]
  assign _T_570 = io_rw_addr == 12'hb91; // @[CSR.scala 177:73:@4932.4]
  assign _T_572 = io_rw_addr == 12'hb12; // @[CSR.scala 177:73:@4933.4]
  assign _T_574 = io_rw_addr == 12'hb92; // @[CSR.scala 177:73:@4934.4]
  assign _T_576 = io_rw_addr == 12'hb13; // @[CSR.scala 177:73:@4935.4]
  assign _T_578 = io_rw_addr == 12'hb93; // @[CSR.scala 177:73:@4936.4]
  assign _T_580 = io_rw_addr == 12'hb14; // @[CSR.scala 177:73:@4937.4]
  assign _T_582 = io_rw_addr == 12'hb94; // @[CSR.scala 177:73:@4938.4]
  assign _T_584 = io_rw_addr == 12'hb15; // @[CSR.scala 177:73:@4939.4]
  assign _T_586 = io_rw_addr == 12'hb95; // @[CSR.scala 177:73:@4940.4]
  assign _T_588 = io_rw_addr == 12'hb16; // @[CSR.scala 177:73:@4941.4]
  assign _T_590 = io_rw_addr == 12'hb96; // @[CSR.scala 177:73:@4942.4]
  assign _T_592 = io_rw_addr == 12'hb17; // @[CSR.scala 177:73:@4943.4]
  assign _T_594 = io_rw_addr == 12'hb97; // @[CSR.scala 177:73:@4944.4]
  assign _T_596 = io_rw_addr == 12'hb18; // @[CSR.scala 177:73:@4945.4]
  assign _T_598 = io_rw_addr == 12'hb98; // @[CSR.scala 177:73:@4946.4]
  assign _T_600 = io_rw_addr == 12'hb19; // @[CSR.scala 177:73:@4947.4]
  assign _T_602 = io_rw_addr == 12'hb99; // @[CSR.scala 177:73:@4948.4]
  assign _T_604 = io_rw_addr == 12'hb1a; // @[CSR.scala 177:73:@4949.4]
  assign _T_606 = io_rw_addr == 12'hb9a; // @[CSR.scala 177:73:@4950.4]
  assign _T_608 = io_rw_addr == 12'hb1b; // @[CSR.scala 177:73:@4951.4]
  assign _T_610 = io_rw_addr == 12'hb9b; // @[CSR.scala 177:73:@4952.4]
  assign _T_612 = io_rw_addr == 12'hb1c; // @[CSR.scala 177:73:@4953.4]
  assign _T_614 = io_rw_addr == 12'hb9c; // @[CSR.scala 177:73:@4954.4]
  assign _T_616 = io_rw_addr == 12'hb1d; // @[CSR.scala 177:73:@4955.4]
  assign _T_618 = io_rw_addr == 12'hb9d; // @[CSR.scala 177:73:@4956.4]
  assign _T_620 = io_rw_addr == 12'hb1e; // @[CSR.scala 177:73:@4957.4]
  assign _T_622 = io_rw_addr == 12'hb9e; // @[CSR.scala 177:73:@4958.4]
  assign _T_624 = io_rw_addr == 12'hb1f; // @[CSR.scala 177:73:@4959.4]
  assign _T_626 = io_rw_addr == 12'hb9f; // @[CSR.scala 177:73:@4960.4]
  assign _T_628 = io_rw_addr == 12'hb20; // @[CSR.scala 177:73:@4961.4]
  assign _T_630 = io_rw_addr == 12'hba0; // @[CSR.scala 177:73:@4962.4]
  assign _T_632 = io_rw_addr == 12'hb21; // @[CSR.scala 177:73:@4963.4]
  assign _T_634 = io_rw_addr == 12'hba1; // @[CSR.scala 177:73:@4964.4]
  assign _T_636 = io_rw_addr == 12'hb22; // @[CSR.scala 177:73:@4965.4]
  assign _T_638 = io_rw_addr == 12'hba2; // @[CSR.scala 177:73:@4966.4]
  assign _T_640 = io_rw_addr == 12'hb80; // @[CSR.scala 177:73:@4967.4]
  assign _T_642 = io_rw_addr == 12'hb82; // @[CSR.scala 177:73:@4968.4]
  assign _T_643 = io_rw_addr[9:8]; // @[CSR.scala 179:54:@4969.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_643; // @[CSR.scala 179:41:@4970.4]
  assign _T_644 = io_rw_addr[11:10]; // @[CSR.scala 180:29:@4971.4]
  assign _T_645 = ~ _T_644; // @[CSR.scala 180:37:@4972.4]
  assign read_only = _T_645 == 2'h0; // @[CSR.scala 180:37:@4973.4]
  assign _T_647 = io_rw_cmd != 3'h5; // @[CSR.scala 181:38:@4974.4]
  assign _T_648 = cpu_ren & _T_647; // @[CSR.scala 181:25:@4975.4]
  assign cpu_wen = _T_648 & priv_sufficient; // @[CSR.scala 181:48:@4976.4]
  assign _T_650 = read_only == 1'h0; // @[CSR.scala 182:24:@4977.4]
  assign wen = cpu_wen & _T_650; // @[CSR.scala 182:21:@4978.4]
  assign _T_651 = io_rw_cmd == 3'h2; // @[Util.scala 23:47:@4979.4]
  assign _T_652 = io_rw_cmd == 3'h3; // @[Util.scala 23:47:@4980.4]
  assign _T_653 = _T_651 | _T_652; // @[Util.scala 23:62:@4981.4]
  assign _T_655 = _T_653 ? io_rw_rdata : 32'h0; // @[CSR.scala 281:9:@4982.4]
  assign _T_656 = _T_655 | io_rw_wdata; // @[CSR.scala 281:49:@4983.4]
  assign _T_659 = _T_652 ? io_rw_wdata : 32'h0; // @[CSR.scala 281:64:@4985.4]
  assign _T_660 = ~ _T_659; // @[CSR.scala 281:60:@4986.4]
  assign wdata = _T_656 & _T_660; // @[CSR.scala 281:58:@4987.4]
  assign _T_662 = io_rw_addr[2:0]; // @[CSR.scala 185:33:@4988.4]
  assign opcode = 8'h1 << _T_662; // @[CSR.scala 185:20:@4989.4]
  assign _T_663 = opcode[0]; // @[CSR.scala 186:40:@4990.4]
  assign insn_call = system_insn & _T_663; // @[CSR.scala 186:31:@4991.4]
  assign _T_664 = opcode[1]; // @[CSR.scala 187:41:@4992.4]
  assign insn_break = system_insn & _T_664; // @[CSR.scala 187:32:@4993.4]
  assign _T_665 = opcode[2]; // @[CSR.scala 188:39:@4994.4]
  assign _T_666 = system_insn & _T_665; // @[CSR.scala 188:30:@4995.4]
  assign insn_ret = _T_666 & priv_sufficient; // @[CSR.scala 188:43:@4996.4]
  assign _T_940 = insn_call | insn_break; // @[CSR.scala 199:24:@5195.4]
  assign _T_942 = {{1'd0}, insn_ret}; // @[Bitwise.scala 48:55:@5198.4]
  assign _T_944 = _T_942 <= 2'h1; // @[CSR.scala 201:50:@5199.4]
  assign _T_946 = _T_944 | reset; // @[CSR.scala 201:9:@5201.4]
  assign _T_948 = _T_946 == 1'h0; // @[CSR.scala 201:9:@5202.4]
  assign _T_951 = io_rw_addr[10]; // @[CSR.scala 208:32:@5211.4]
  assign _T_953 = _T_951 == 1'h0; // @[CSR.scala 208:21:@5212.4]
  assign _T_954 = insn_ret & _T_953; // @[CSR.scala 208:18:@5213.4]
  assign _GEN_3 = _T_954 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 208:38:@5214.4]
  assign _GEN_4 = _T_954 ? 1'h1 : reg_mstatus_mpie; // @[CSR.scala 208:38:@5214.4]
  assign new_prv = _T_954 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 208:38:@5214.4]
  assign _GEN_148 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 218:35:@5222.6]
  assign _T_958 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@5222.6]
  assign _T_959 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@5223.6]
  assign _GEN_7 = insn_call ? 32'h80000004 : reg_mepc; // @[CSR.scala 216:18:@5220.4]
  assign _GEN_8 = insn_call ? {{28'd0}, _T_959} : reg_mcause; // @[CSR.scala 216:18:@5220.4]
  assign _GEN_9 = insn_call ? io_pc : reg_mepc; // @[CSR.scala 216:18:@5220.4]
  assign _GEN_10 = insn_break ? 32'h80000004 : _GEN_7; // @[CSR.scala 223:19:@5227.4]
  assign _GEN_11 = insn_break ? 32'h3 : _GEN_8; // @[CSR.scala 223:19:@5227.4]
  assign _GEN_12 = insn_break ? io_pc : _GEN_9; // @[CSR.scala 223:19:@5227.4]
  assign _GEN_14 = io_xcpt ? io_cause : _GEN_11; // @[CSR.scala 229:17:@5232.4]
  assign _GEN_15 = io_xcpt ? io_pc : _GEN_12; // @[CSR.scala 229:17:@5232.4]
  assign _GEN_16 = io_xcpt ? io_tval : reg_mtval; // @[CSR.scala 229:17:@5232.4]
  assign _T_965 = _T_478 ? _T_249 : 64'h0; // @[Mux.scala 19:72:@5240.4]
  assign _T_967 = _T_480 ? _T_261 : 64'h0; // @[Mux.scala 19:72:@5241.4]
  assign _T_969 = _T_482 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:@5242.4]
  assign _T_975 = _T_488 ? 31'h40000100 : 31'h0; // @[Mux.scala 19:72:@5245.4]
  assign _T_977 = _T_490 ? read_mstatus : 32'h0; // @[Mux.scala 19:72:@5246.4]
  assign _T_979 = _T_492 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:@5247.4]
  assign _T_981 = _T_494 ? _T_468 : 16'h0; // @[Mux.scala 19:72:@5248.4]
  assign _T_983 = _T_496 ? _T_474 : 16'h0; // @[Mux.scala 19:72:@5249.4]
  assign _T_985 = _T_498 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:@5250.4]
  assign _T_987 = _T_500 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:@5251.4]
  assign _T_989 = _T_502 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:@5252.4]
  assign _T_991 = _T_504 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:@5253.4]
  assign _T_995 = _T_508 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:@5255.4]
  assign _T_997 = _T_510 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:@5256.4]
  assign _T_999 = _T_512 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@5257.4]
  assign _T_1001 = _T_514 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@5258.4]
  assign _T_1003 = _T_516 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@5259.4]
  assign _T_1005 = _T_518 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@5260.4]
  assign _T_1007 = _T_520 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@5261.4]
  assign _T_1009 = _T_522 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@5262.4]
  assign _T_1011 = _T_524 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@5263.4]
  assign _T_1013 = _T_526 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@5264.4]
  assign _T_1015 = _T_528 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@5265.4]
  assign _T_1017 = _T_530 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@5266.4]
  assign _T_1019 = _T_532 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@5267.4]
  assign _T_1021 = _T_534 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@5268.4]
  assign _T_1023 = _T_536 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@5269.4]
  assign _T_1025 = _T_538 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@5270.4]
  assign _T_1027 = _T_540 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@5271.4]
  assign _T_1029 = _T_542 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@5272.4]
  assign _T_1031 = _T_544 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@5273.4]
  assign _T_1033 = _T_546 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@5274.4]
  assign _T_1035 = _T_548 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@5275.4]
  assign _T_1037 = _T_550 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@5276.4]
  assign _T_1039 = _T_552 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@5277.4]
  assign _T_1041 = _T_554 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@5278.4]
  assign _T_1043 = _T_556 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@5279.4]
  assign _T_1045 = _T_558 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@5280.4]
  assign _T_1047 = _T_560 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@5281.4]
  assign _T_1049 = _T_562 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@5282.4]
  assign _T_1051 = _T_564 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@5283.4]
  assign _T_1053 = _T_566 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@5284.4]
  assign _T_1055 = _T_568 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@5285.4]
  assign _T_1057 = _T_570 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@5286.4]
  assign _T_1059 = _T_572 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@5287.4]
  assign _T_1061 = _T_574 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@5288.4]
  assign _T_1063 = _T_576 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@5289.4]
  assign _T_1065 = _T_578 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@5290.4]
  assign _T_1067 = _T_580 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@5291.4]
  assign _T_1069 = _T_582 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@5292.4]
  assign _T_1071 = _T_584 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@5293.4]
  assign _T_1073 = _T_586 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@5294.4]
  assign _T_1075 = _T_588 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@5295.4]
  assign _T_1077 = _T_590 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@5296.4]
  assign _T_1079 = _T_592 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@5297.4]
  assign _T_1081 = _T_594 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@5298.4]
  assign _T_1083 = _T_596 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@5299.4]
  assign _T_1085 = _T_598 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@5300.4]
  assign _T_1087 = _T_600 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@5301.4]
  assign _T_1089 = _T_602 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@5302.4]
  assign _T_1091 = _T_604 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@5303.4]
  assign _T_1093 = _T_606 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@5304.4]
  assign _T_1095 = _T_608 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@5305.4]
  assign _T_1097 = _T_610 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@5306.4]
  assign _T_1099 = _T_612 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@5307.4]
  assign _T_1101 = _T_614 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@5308.4]
  assign _T_1103 = _T_616 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@5309.4]
  assign _T_1105 = _T_618 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@5310.4]
  assign _T_1107 = _T_620 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@5311.4]
  assign _T_1109 = _T_622 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@5312.4]
  assign _T_1111 = _T_624 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@5313.4]
  assign _T_1113 = _T_626 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@5314.4]
  assign _T_1115 = _T_628 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@5315.4]
  assign _T_1117 = _T_630 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@5316.4]
  assign _T_1119 = _T_632 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@5317.4]
  assign _T_1121 = _T_634 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@5318.4]
  assign _T_1123 = _T_636 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@5319.4]
  assign _T_1125 = _T_638 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@5320.4]
  assign _T_1130 = _T_965 | _T_967; // @[Mux.scala 19:72:@5323.4]
  assign _GEN_149 = {{48'd0}, _T_969}; // @[Mux.scala 19:72:@5324.4]
  assign _T_1131 = _T_1130 | _GEN_149; // @[Mux.scala 19:72:@5324.4]
  assign _GEN_150 = {{33'd0}, _T_975}; // @[Mux.scala 19:72:@5327.4]
  assign _T_1134 = _T_1131 | _GEN_150; // @[Mux.scala 19:72:@5327.4]
  assign _GEN_151 = {{32'd0}, _T_977}; // @[Mux.scala 19:72:@5328.4]
  assign _T_1135 = _T_1134 | _GEN_151; // @[Mux.scala 19:72:@5328.4]
  assign _GEN_152 = {{55'd0}, _T_979}; // @[Mux.scala 19:72:@5329.4]
  assign _T_1136 = _T_1135 | _GEN_152; // @[Mux.scala 19:72:@5329.4]
  assign _GEN_153 = {{48'd0}, _T_981}; // @[Mux.scala 19:72:@5330.4]
  assign _T_1137 = _T_1136 | _GEN_153; // @[Mux.scala 19:72:@5330.4]
  assign _GEN_154 = {{48'd0}, _T_983}; // @[Mux.scala 19:72:@5331.4]
  assign _T_1138 = _T_1137 | _GEN_154; // @[Mux.scala 19:72:@5331.4]
  assign _GEN_155 = {{32'd0}, _T_985}; // @[Mux.scala 19:72:@5332.4]
  assign _T_1139 = _T_1138 | _GEN_155; // @[Mux.scala 19:72:@5332.4]
  assign _GEN_156 = {{32'd0}, _T_987}; // @[Mux.scala 19:72:@5333.4]
  assign _T_1140 = _T_1139 | _GEN_156; // @[Mux.scala 19:72:@5333.4]
  assign _GEN_157 = {{32'd0}, _T_989}; // @[Mux.scala 19:72:@5334.4]
  assign _T_1141 = _T_1140 | _GEN_157; // @[Mux.scala 19:72:@5334.4]
  assign _GEN_158 = {{32'd0}, _T_991}; // @[Mux.scala 19:72:@5335.4]
  assign _T_1142 = _T_1141 | _GEN_158; // @[Mux.scala 19:72:@5335.4]
  assign _GEN_159 = {{32'd0}, _T_995}; // @[Mux.scala 19:72:@5337.4]
  assign _T_1144 = _T_1142 | _GEN_159; // @[Mux.scala 19:72:@5337.4]
  assign _GEN_160 = {{32'd0}, _T_997}; // @[Mux.scala 19:72:@5338.4]
  assign _T_1145 = _T_1144 | _GEN_160; // @[Mux.scala 19:72:@5338.4]
  assign _GEN_161 = {{24'd0}, _T_999}; // @[Mux.scala 19:72:@5339.4]
  assign _T_1146 = _T_1145 | _GEN_161; // @[Mux.scala 19:72:@5339.4]
  assign _GEN_162 = {{24'd0}, _T_1001}; // @[Mux.scala 19:72:@5340.4]
  assign _T_1147 = _T_1146 | _GEN_162; // @[Mux.scala 19:72:@5340.4]
  assign _GEN_163 = {{24'd0}, _T_1003}; // @[Mux.scala 19:72:@5341.4]
  assign _T_1148 = _T_1147 | _GEN_163; // @[Mux.scala 19:72:@5341.4]
  assign _GEN_164 = {{24'd0}, _T_1005}; // @[Mux.scala 19:72:@5342.4]
  assign _T_1149 = _T_1148 | _GEN_164; // @[Mux.scala 19:72:@5342.4]
  assign _GEN_165 = {{24'd0}, _T_1007}; // @[Mux.scala 19:72:@5343.4]
  assign _T_1150 = _T_1149 | _GEN_165; // @[Mux.scala 19:72:@5343.4]
  assign _GEN_166 = {{24'd0}, _T_1009}; // @[Mux.scala 19:72:@5344.4]
  assign _T_1151 = _T_1150 | _GEN_166; // @[Mux.scala 19:72:@5344.4]
  assign _GEN_167 = {{24'd0}, _T_1011}; // @[Mux.scala 19:72:@5345.4]
  assign _T_1152 = _T_1151 | _GEN_167; // @[Mux.scala 19:72:@5345.4]
  assign _GEN_168 = {{24'd0}, _T_1013}; // @[Mux.scala 19:72:@5346.4]
  assign _T_1153 = _T_1152 | _GEN_168; // @[Mux.scala 19:72:@5346.4]
  assign _GEN_169 = {{24'd0}, _T_1015}; // @[Mux.scala 19:72:@5347.4]
  assign _T_1154 = _T_1153 | _GEN_169; // @[Mux.scala 19:72:@5347.4]
  assign _GEN_170 = {{24'd0}, _T_1017}; // @[Mux.scala 19:72:@5348.4]
  assign _T_1155 = _T_1154 | _GEN_170; // @[Mux.scala 19:72:@5348.4]
  assign _GEN_171 = {{24'd0}, _T_1019}; // @[Mux.scala 19:72:@5349.4]
  assign _T_1156 = _T_1155 | _GEN_171; // @[Mux.scala 19:72:@5349.4]
  assign _GEN_172 = {{24'd0}, _T_1021}; // @[Mux.scala 19:72:@5350.4]
  assign _T_1157 = _T_1156 | _GEN_172; // @[Mux.scala 19:72:@5350.4]
  assign _GEN_173 = {{24'd0}, _T_1023}; // @[Mux.scala 19:72:@5351.4]
  assign _T_1158 = _T_1157 | _GEN_173; // @[Mux.scala 19:72:@5351.4]
  assign _GEN_174 = {{24'd0}, _T_1025}; // @[Mux.scala 19:72:@5352.4]
  assign _T_1159 = _T_1158 | _GEN_174; // @[Mux.scala 19:72:@5352.4]
  assign _GEN_175 = {{24'd0}, _T_1027}; // @[Mux.scala 19:72:@5353.4]
  assign _T_1160 = _T_1159 | _GEN_175; // @[Mux.scala 19:72:@5353.4]
  assign _GEN_176 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:@5354.4]
  assign _T_1161 = _T_1160 | _GEN_176; // @[Mux.scala 19:72:@5354.4]
  assign _GEN_177 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:@5355.4]
  assign _T_1162 = _T_1161 | _GEN_177; // @[Mux.scala 19:72:@5355.4]
  assign _GEN_178 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:@5356.4]
  assign _T_1163 = _T_1162 | _GEN_178; // @[Mux.scala 19:72:@5356.4]
  assign _GEN_179 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:@5357.4]
  assign _T_1164 = _T_1163 | _GEN_179; // @[Mux.scala 19:72:@5357.4]
  assign _GEN_180 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:@5358.4]
  assign _T_1165 = _T_1164 | _GEN_180; // @[Mux.scala 19:72:@5358.4]
  assign _GEN_181 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:@5359.4]
  assign _T_1166 = _T_1165 | _GEN_181; // @[Mux.scala 19:72:@5359.4]
  assign _GEN_182 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:@5360.4]
  assign _T_1167 = _T_1166 | _GEN_182; // @[Mux.scala 19:72:@5360.4]
  assign _GEN_183 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:@5361.4]
  assign _T_1168 = _T_1167 | _GEN_183; // @[Mux.scala 19:72:@5361.4]
  assign _GEN_184 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:@5362.4]
  assign _T_1169 = _T_1168 | _GEN_184; // @[Mux.scala 19:72:@5362.4]
  assign _GEN_185 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:@5363.4]
  assign _T_1170 = _T_1169 | _GEN_185; // @[Mux.scala 19:72:@5363.4]
  assign _GEN_186 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:@5364.4]
  assign _T_1171 = _T_1170 | _GEN_186; // @[Mux.scala 19:72:@5364.4]
  assign _GEN_187 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:@5365.4]
  assign _T_1172 = _T_1171 | _GEN_187; // @[Mux.scala 19:72:@5365.4]
  assign _GEN_188 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:@5366.4]
  assign _T_1173 = _T_1172 | _GEN_188; // @[Mux.scala 19:72:@5366.4]
  assign _GEN_189 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:@5367.4]
  assign _T_1174 = _T_1173 | _GEN_189; // @[Mux.scala 19:72:@5367.4]
  assign _GEN_190 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:@5368.4]
  assign _T_1175 = _T_1174 | _GEN_190; // @[Mux.scala 19:72:@5368.4]
  assign _GEN_191 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:@5369.4]
  assign _T_1176 = _T_1175 | _GEN_191; // @[Mux.scala 19:72:@5369.4]
  assign _GEN_192 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:@5370.4]
  assign _T_1177 = _T_1176 | _GEN_192; // @[Mux.scala 19:72:@5370.4]
  assign _GEN_193 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:@5371.4]
  assign _T_1178 = _T_1177 | _GEN_193; // @[Mux.scala 19:72:@5371.4]
  assign _GEN_194 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:@5372.4]
  assign _T_1179 = _T_1178 | _GEN_194; // @[Mux.scala 19:72:@5372.4]
  assign _GEN_195 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:@5373.4]
  assign _T_1180 = _T_1179 | _GEN_195; // @[Mux.scala 19:72:@5373.4]
  assign _GEN_196 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:@5374.4]
  assign _T_1181 = _T_1180 | _GEN_196; // @[Mux.scala 19:72:@5374.4]
  assign _GEN_197 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:@5375.4]
  assign _T_1182 = _T_1181 | _GEN_197; // @[Mux.scala 19:72:@5375.4]
  assign _GEN_198 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:@5376.4]
  assign _T_1183 = _T_1182 | _GEN_198; // @[Mux.scala 19:72:@5376.4]
  assign _GEN_199 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:@5377.4]
  assign _T_1184 = _T_1183 | _GEN_199; // @[Mux.scala 19:72:@5377.4]
  assign _GEN_200 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:@5378.4]
  assign _T_1185 = _T_1184 | _GEN_200; // @[Mux.scala 19:72:@5378.4]
  assign _GEN_201 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:@5379.4]
  assign _T_1186 = _T_1185 | _GEN_201; // @[Mux.scala 19:72:@5379.4]
  assign _GEN_202 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:@5380.4]
  assign _T_1187 = _T_1186 | _GEN_202; // @[Mux.scala 19:72:@5380.4]
  assign _GEN_203 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:@5381.4]
  assign _T_1188 = _T_1187 | _GEN_203; // @[Mux.scala 19:72:@5381.4]
  assign _GEN_204 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:@5382.4]
  assign _T_1189 = _T_1188 | _GEN_204; // @[Mux.scala 19:72:@5382.4]
  assign _GEN_205 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:@5383.4]
  assign _T_1190 = _T_1189 | _GEN_205; // @[Mux.scala 19:72:@5383.4]
  assign _GEN_206 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:@5384.4]
  assign _T_1191 = _T_1190 | _GEN_206; // @[Mux.scala 19:72:@5384.4]
  assign _GEN_207 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:@5385.4]
  assign _T_1192 = _T_1191 | _GEN_207; // @[Mux.scala 19:72:@5385.4]
  assign _GEN_208 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:@5386.4]
  assign _T_1193 = _T_1192 | _GEN_208; // @[Mux.scala 19:72:@5386.4]
  assign _GEN_209 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:@5387.4]
  assign _T_1194 = _T_1193 | _GEN_209; // @[Mux.scala 19:72:@5387.4]
  assign _GEN_210 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:@5388.4]
  assign _T_1195 = _T_1194 | _GEN_210; // @[Mux.scala 19:72:@5388.4]
  assign _GEN_211 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:@5389.4]
  assign _T_1196 = _T_1195 | _GEN_211; // @[Mux.scala 19:72:@5389.4]
  assign _GEN_212 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:@5390.4]
  assign _T_1197 = _T_1196 | _GEN_212; // @[Mux.scala 19:72:@5390.4]
  assign _GEN_213 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:@5391.4]
  assign _T_1198 = _T_1197 | _GEN_213; // @[Mux.scala 19:72:@5391.4]
  assign _GEN_214 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:@5392.4]
  assign _T_1199 = _T_1198 | _GEN_214; // @[Mux.scala 19:72:@5392.4]
  assign _GEN_215 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:@5393.4]
  assign _T_1200 = _T_1199 | _GEN_215; // @[Mux.scala 19:72:@5393.4]
  assign _GEN_216 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:@5394.4]
  assign _T_1201 = _T_1200 | _GEN_216; // @[Mux.scala 19:72:@5394.4]
  assign _GEN_217 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:@5395.4]
  assign _T_1202 = _T_1201 | _GEN_217; // @[Mux.scala 19:72:@5395.4]
  assign _GEN_218 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:@5396.4]
  assign _T_1203 = _T_1202 | _GEN_218; // @[Mux.scala 19:72:@5396.4]
  assign _GEN_219 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:@5397.4]
  assign _T_1204 = _T_1203 | _GEN_219; // @[Mux.scala 19:72:@5397.4]
  assign _GEN_220 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:@5398.4]
  assign _T_1205 = _T_1204 | _GEN_220; // @[Mux.scala 19:72:@5398.4]
  assign _GEN_221 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:@5399.4]
  assign _T_1206 = _T_1205 | _GEN_221; // @[Mux.scala 19:72:@5399.4]
  assign _GEN_222 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:@5400.4]
  assign _T_1207 = _T_1206 | _GEN_222; // @[Mux.scala 19:72:@5400.4]
  assign _GEN_223 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:@5401.4]
  assign _T_1208 = _T_1207 | _GEN_223; // @[Mux.scala 19:72:@5401.4]
  assign _GEN_224 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:@5402.4]
  assign _T_1209 = _T_1208 | _GEN_224; // @[Mux.scala 19:72:@5402.4]
  assign _T_1220 = wdata[3]; // @[CSR.scala 245:39:@5415.8]
  assign _T_1222 = wdata[7]; // @[CSR.scala 245:39:@5419.8]
  assign _GEN_17 = _T_490 ? _T_1220 : _GEN_3; // @[CSR.scala 244:39:@5409.6]
  assign _GEN_18 = _T_490 ? _T_1222 : _GEN_4; // @[CSR.scala 244:39:@5409.6]
  assign _T_1233 = wdata[15:0]; // @[:@5438.8 :@5439.8]
  assign _T_1235 = _T_1233[3]; // @[CSR.scala 250:35:@5442.8]
  assign _T_1237 = _T_1233[7]; // @[CSR.scala 250:35:@5446.8]
  assign _GEN_19 = _T_494 ? _T_1235 : reg_mip_msip; // @[CSR.scala 249:35:@5436.6]
  assign _GEN_20 = _T_496 ? _T_1235 : reg_mie_msip; // @[CSR.scala 253:35:@5456.6]
  assign _GEN_21 = _T_496 ? _T_1237 : reg_mie_mtip; // @[CSR.scala 253:35:@5456.6]
  assign _T_1253 = wdata[7:0]; // @[CSR.scala 277:47:@5478.8]
  assign _T_1254 = _T_264[31:0]; // @[CSR.scala 277:72:@5479.8]
  assign _T_1255 = {_T_1253,_T_1254}; // @[Cat.scala 30:58:@5480.8]
  assign _GEN_22 = _T_514 ? {{1'd0}, _T_1255} : _T_265; // @[CSR.scala 277:29:@5477.6]
  assign _T_1256 = _T_264[39:32]; // @[CSR.scala 278:45:@5484.8]
  assign _T_1257 = {_T_1256,wdata}; // @[Cat.scala 30:58:@5485.8]
  assign _GEN_23 = _T_512 ? {{1'd0}, _T_1257} : _GEN_22; // @[CSR.scala 278:29:@5483.6]
  assign _T_1259 = _T_267[31:0]; // @[CSR.scala 277:72:@5490.8]
  assign _T_1260 = {_T_1253,_T_1259}; // @[Cat.scala 30:58:@5491.8]
  assign _GEN_24 = _T_518 ? {{1'd0}, _T_1260} : _T_268; // @[CSR.scala 277:29:@5488.6]
  assign _T_1261 = _T_267[39:32]; // @[CSR.scala 278:45:@5495.8]
  assign _T_1262 = {_T_1261,wdata}; // @[Cat.scala 30:58:@5496.8]
  assign _GEN_25 = _T_516 ? {{1'd0}, _T_1262} : _GEN_24; // @[CSR.scala 278:29:@5494.6]
  assign _T_1264 = _T_270[31:0]; // @[CSR.scala 277:72:@5501.8]
  assign _T_1265 = {_T_1253,_T_1264}; // @[Cat.scala 30:58:@5502.8]
  assign _GEN_26 = _T_522 ? {{1'd0}, _T_1265} : _T_271; // @[CSR.scala 277:29:@5499.6]
  assign _T_1266 = _T_270[39:32]; // @[CSR.scala 278:45:@5506.8]
  assign _T_1267 = {_T_1266,wdata}; // @[Cat.scala 30:58:@5507.8]
  assign _GEN_27 = _T_520 ? {{1'd0}, _T_1267} : _GEN_26; // @[CSR.scala 278:29:@5505.6]
  assign _T_1269 = _T_273[31:0]; // @[CSR.scala 277:72:@5512.8]
  assign _T_1270 = {_T_1253,_T_1269}; // @[Cat.scala 30:58:@5513.8]
  assign _GEN_28 = _T_526 ? {{1'd0}, _T_1270} : _T_274; // @[CSR.scala 277:29:@5510.6]
  assign _T_1271 = _T_273[39:32]; // @[CSR.scala 278:45:@5517.8]
  assign _T_1272 = {_T_1271,wdata}; // @[Cat.scala 30:58:@5518.8]
  assign _GEN_29 = _T_524 ? {{1'd0}, _T_1272} : _GEN_28; // @[CSR.scala 278:29:@5516.6]
  assign _T_1274 = _T_276[31:0]; // @[CSR.scala 277:72:@5523.8]
  assign _T_1275 = {_T_1253,_T_1274}; // @[Cat.scala 30:58:@5524.8]
  assign _GEN_30 = _T_530 ? {{1'd0}, _T_1275} : _T_277; // @[CSR.scala 277:29:@5521.6]
  assign _T_1276 = _T_276[39:32]; // @[CSR.scala 278:45:@5528.8]
  assign _T_1277 = {_T_1276,wdata}; // @[Cat.scala 30:58:@5529.8]
  assign _GEN_31 = _T_528 ? {{1'd0}, _T_1277} : _GEN_30; // @[CSR.scala 278:29:@5527.6]
  assign _T_1279 = _T_279[31:0]; // @[CSR.scala 277:72:@5534.8]
  assign _T_1280 = {_T_1253,_T_1279}; // @[Cat.scala 30:58:@5535.8]
  assign _GEN_32 = _T_534 ? {{1'd0}, _T_1280} : _T_280; // @[CSR.scala 277:29:@5532.6]
  assign _T_1281 = _T_279[39:32]; // @[CSR.scala 278:45:@5539.8]
  assign _T_1282 = {_T_1281,wdata}; // @[Cat.scala 30:58:@5540.8]
  assign _GEN_33 = _T_532 ? {{1'd0}, _T_1282} : _GEN_32; // @[CSR.scala 278:29:@5538.6]
  assign _T_1284 = _T_282[31:0]; // @[CSR.scala 277:72:@5545.8]
  assign _T_1285 = {_T_1253,_T_1284}; // @[Cat.scala 30:58:@5546.8]
  assign _GEN_34 = _T_538 ? {{1'd0}, _T_1285} : _T_283; // @[CSR.scala 277:29:@5543.6]
  assign _T_1286 = _T_282[39:32]; // @[CSR.scala 278:45:@5550.8]
  assign _T_1287 = {_T_1286,wdata}; // @[Cat.scala 30:58:@5551.8]
  assign _GEN_35 = _T_536 ? {{1'd0}, _T_1287} : _GEN_34; // @[CSR.scala 278:29:@5549.6]
  assign _T_1289 = _T_285[31:0]; // @[CSR.scala 277:72:@5556.8]
  assign _T_1290 = {_T_1253,_T_1289}; // @[Cat.scala 30:58:@5557.8]
  assign _GEN_36 = _T_542 ? {{1'd0}, _T_1290} : _T_286; // @[CSR.scala 277:29:@5554.6]
  assign _T_1291 = _T_285[39:32]; // @[CSR.scala 278:45:@5561.8]
  assign _T_1292 = {_T_1291,wdata}; // @[Cat.scala 30:58:@5562.8]
  assign _GEN_37 = _T_540 ? {{1'd0}, _T_1292} : _GEN_36; // @[CSR.scala 278:29:@5560.6]
  assign _T_1294 = _T_288[31:0]; // @[CSR.scala 277:72:@5567.8]
  assign _T_1295 = {_T_1253,_T_1294}; // @[Cat.scala 30:58:@5568.8]
  assign _GEN_38 = _T_546 ? {{1'd0}, _T_1295} : _T_289; // @[CSR.scala 277:29:@5565.6]
  assign _T_1296 = _T_288[39:32]; // @[CSR.scala 278:45:@5572.8]
  assign _T_1297 = {_T_1296,wdata}; // @[Cat.scala 30:58:@5573.8]
  assign _GEN_39 = _T_544 ? {{1'd0}, _T_1297} : _GEN_38; // @[CSR.scala 278:29:@5571.6]
  assign _T_1299 = _T_291[31:0]; // @[CSR.scala 277:72:@5578.8]
  assign _T_1300 = {_T_1253,_T_1299}; // @[Cat.scala 30:58:@5579.8]
  assign _GEN_40 = _T_550 ? {{1'd0}, _T_1300} : _T_292; // @[CSR.scala 277:29:@5576.6]
  assign _T_1301 = _T_291[39:32]; // @[CSR.scala 278:45:@5583.8]
  assign _T_1302 = {_T_1301,wdata}; // @[Cat.scala 30:58:@5584.8]
  assign _GEN_41 = _T_548 ? {{1'd0}, _T_1302} : _GEN_40; // @[CSR.scala 278:29:@5582.6]
  assign _T_1304 = _T_294[31:0]; // @[CSR.scala 277:72:@5589.8]
  assign _T_1305 = {_T_1253,_T_1304}; // @[Cat.scala 30:58:@5590.8]
  assign _GEN_42 = _T_554 ? {{1'd0}, _T_1305} : _T_295; // @[CSR.scala 277:29:@5587.6]
  assign _T_1306 = _T_294[39:32]; // @[CSR.scala 278:45:@5594.8]
  assign _T_1307 = {_T_1306,wdata}; // @[Cat.scala 30:58:@5595.8]
  assign _GEN_43 = _T_552 ? {{1'd0}, _T_1307} : _GEN_42; // @[CSR.scala 278:29:@5593.6]
  assign _T_1309 = _T_297[31:0]; // @[CSR.scala 277:72:@5600.8]
  assign _T_1310 = {_T_1253,_T_1309}; // @[Cat.scala 30:58:@5601.8]
  assign _GEN_44 = _T_558 ? {{1'd0}, _T_1310} : _T_298; // @[CSR.scala 277:29:@5598.6]
  assign _T_1311 = _T_297[39:32]; // @[CSR.scala 278:45:@5605.8]
  assign _T_1312 = {_T_1311,wdata}; // @[Cat.scala 30:58:@5606.8]
  assign _GEN_45 = _T_556 ? {{1'd0}, _T_1312} : _GEN_44; // @[CSR.scala 278:29:@5604.6]
  assign _T_1314 = _T_300[31:0]; // @[CSR.scala 277:72:@5611.8]
  assign _T_1315 = {_T_1253,_T_1314}; // @[Cat.scala 30:58:@5612.8]
  assign _GEN_46 = _T_562 ? {{1'd0}, _T_1315} : _T_301; // @[CSR.scala 277:29:@5609.6]
  assign _T_1316 = _T_300[39:32]; // @[CSR.scala 278:45:@5616.8]
  assign _T_1317 = {_T_1316,wdata}; // @[Cat.scala 30:58:@5617.8]
  assign _GEN_47 = _T_560 ? {{1'd0}, _T_1317} : _GEN_46; // @[CSR.scala 278:29:@5615.6]
  assign _T_1319 = _T_303[31:0]; // @[CSR.scala 277:72:@5622.8]
  assign _T_1320 = {_T_1253,_T_1319}; // @[Cat.scala 30:58:@5623.8]
  assign _GEN_48 = _T_566 ? {{1'd0}, _T_1320} : _T_304; // @[CSR.scala 277:29:@5620.6]
  assign _T_1321 = _T_303[39:32]; // @[CSR.scala 278:45:@5627.8]
  assign _T_1322 = {_T_1321,wdata}; // @[Cat.scala 30:58:@5628.8]
  assign _GEN_49 = _T_564 ? {{1'd0}, _T_1322} : _GEN_48; // @[CSR.scala 278:29:@5626.6]
  assign _T_1324 = _T_306[31:0]; // @[CSR.scala 277:72:@5633.8]
  assign _T_1325 = {_T_1253,_T_1324}; // @[Cat.scala 30:58:@5634.8]
  assign _GEN_50 = _T_570 ? {{1'd0}, _T_1325} : _T_307; // @[CSR.scala 277:29:@5631.6]
  assign _T_1326 = _T_306[39:32]; // @[CSR.scala 278:45:@5638.8]
  assign _T_1327 = {_T_1326,wdata}; // @[Cat.scala 30:58:@5639.8]
  assign _GEN_51 = _T_568 ? {{1'd0}, _T_1327} : _GEN_50; // @[CSR.scala 278:29:@5637.6]
  assign _T_1329 = _T_309[31:0]; // @[CSR.scala 277:72:@5644.8]
  assign _T_1330 = {_T_1253,_T_1329}; // @[Cat.scala 30:58:@5645.8]
  assign _GEN_52 = _T_574 ? {{1'd0}, _T_1330} : _T_310; // @[CSR.scala 277:29:@5642.6]
  assign _T_1331 = _T_309[39:32]; // @[CSR.scala 278:45:@5649.8]
  assign _T_1332 = {_T_1331,wdata}; // @[Cat.scala 30:58:@5650.8]
  assign _GEN_53 = _T_572 ? {{1'd0}, _T_1332} : _GEN_52; // @[CSR.scala 278:29:@5648.6]
  assign _T_1334 = _T_312[31:0]; // @[CSR.scala 277:72:@5655.8]
  assign _T_1335 = {_T_1253,_T_1334}; // @[Cat.scala 30:58:@5656.8]
  assign _GEN_54 = _T_578 ? {{1'd0}, _T_1335} : _T_313; // @[CSR.scala 277:29:@5653.6]
  assign _T_1336 = _T_312[39:32]; // @[CSR.scala 278:45:@5660.8]
  assign _T_1337 = {_T_1336,wdata}; // @[Cat.scala 30:58:@5661.8]
  assign _GEN_55 = _T_576 ? {{1'd0}, _T_1337} : _GEN_54; // @[CSR.scala 278:29:@5659.6]
  assign _T_1339 = _T_315[31:0]; // @[CSR.scala 277:72:@5666.8]
  assign _T_1340 = {_T_1253,_T_1339}; // @[Cat.scala 30:58:@5667.8]
  assign _GEN_56 = _T_582 ? {{1'd0}, _T_1340} : _T_316; // @[CSR.scala 277:29:@5664.6]
  assign _T_1341 = _T_315[39:32]; // @[CSR.scala 278:45:@5671.8]
  assign _T_1342 = {_T_1341,wdata}; // @[Cat.scala 30:58:@5672.8]
  assign _GEN_57 = _T_580 ? {{1'd0}, _T_1342} : _GEN_56; // @[CSR.scala 278:29:@5670.6]
  assign _T_1344 = _T_318[31:0]; // @[CSR.scala 277:72:@5677.8]
  assign _T_1345 = {_T_1253,_T_1344}; // @[Cat.scala 30:58:@5678.8]
  assign _GEN_58 = _T_586 ? {{1'd0}, _T_1345} : _T_319; // @[CSR.scala 277:29:@5675.6]
  assign _T_1346 = _T_318[39:32]; // @[CSR.scala 278:45:@5682.8]
  assign _T_1347 = {_T_1346,wdata}; // @[Cat.scala 30:58:@5683.8]
  assign _GEN_59 = _T_584 ? {{1'd0}, _T_1347} : _GEN_58; // @[CSR.scala 278:29:@5681.6]
  assign _T_1349 = _T_321[31:0]; // @[CSR.scala 277:72:@5688.8]
  assign _T_1350 = {_T_1253,_T_1349}; // @[Cat.scala 30:58:@5689.8]
  assign _GEN_60 = _T_590 ? {{1'd0}, _T_1350} : _T_322; // @[CSR.scala 277:29:@5686.6]
  assign _T_1351 = _T_321[39:32]; // @[CSR.scala 278:45:@5693.8]
  assign _T_1352 = {_T_1351,wdata}; // @[Cat.scala 30:58:@5694.8]
  assign _GEN_61 = _T_588 ? {{1'd0}, _T_1352} : _GEN_60; // @[CSR.scala 278:29:@5692.6]
  assign _T_1354 = _T_324[31:0]; // @[CSR.scala 277:72:@5699.8]
  assign _T_1355 = {_T_1253,_T_1354}; // @[Cat.scala 30:58:@5700.8]
  assign _GEN_62 = _T_594 ? {{1'd0}, _T_1355} : _T_325; // @[CSR.scala 277:29:@5697.6]
  assign _T_1356 = _T_324[39:32]; // @[CSR.scala 278:45:@5704.8]
  assign _T_1357 = {_T_1356,wdata}; // @[Cat.scala 30:58:@5705.8]
  assign _GEN_63 = _T_592 ? {{1'd0}, _T_1357} : _GEN_62; // @[CSR.scala 278:29:@5703.6]
  assign _T_1359 = _T_327[31:0]; // @[CSR.scala 277:72:@5710.8]
  assign _T_1360 = {_T_1253,_T_1359}; // @[Cat.scala 30:58:@5711.8]
  assign _GEN_64 = _T_598 ? {{1'd0}, _T_1360} : _T_328; // @[CSR.scala 277:29:@5708.6]
  assign _T_1361 = _T_327[39:32]; // @[CSR.scala 278:45:@5715.8]
  assign _T_1362 = {_T_1361,wdata}; // @[Cat.scala 30:58:@5716.8]
  assign _GEN_65 = _T_596 ? {{1'd0}, _T_1362} : _GEN_64; // @[CSR.scala 278:29:@5714.6]
  assign _T_1364 = _T_330[31:0]; // @[CSR.scala 277:72:@5721.8]
  assign _T_1365 = {_T_1253,_T_1364}; // @[Cat.scala 30:58:@5722.8]
  assign _GEN_66 = _T_602 ? {{1'd0}, _T_1365} : _T_331; // @[CSR.scala 277:29:@5719.6]
  assign _T_1366 = _T_330[39:32]; // @[CSR.scala 278:45:@5726.8]
  assign _T_1367 = {_T_1366,wdata}; // @[Cat.scala 30:58:@5727.8]
  assign _GEN_67 = _T_600 ? {{1'd0}, _T_1367} : _GEN_66; // @[CSR.scala 278:29:@5725.6]
  assign _T_1369 = _T_333[31:0]; // @[CSR.scala 277:72:@5732.8]
  assign _T_1370 = {_T_1253,_T_1369}; // @[Cat.scala 30:58:@5733.8]
  assign _GEN_68 = _T_606 ? {{1'd0}, _T_1370} : _T_334; // @[CSR.scala 277:29:@5730.6]
  assign _T_1371 = _T_333[39:32]; // @[CSR.scala 278:45:@5737.8]
  assign _T_1372 = {_T_1371,wdata}; // @[Cat.scala 30:58:@5738.8]
  assign _GEN_69 = _T_604 ? {{1'd0}, _T_1372} : _GEN_68; // @[CSR.scala 278:29:@5736.6]
  assign _T_1374 = _T_336[31:0]; // @[CSR.scala 277:72:@5743.8]
  assign _T_1375 = {_T_1253,_T_1374}; // @[Cat.scala 30:58:@5744.8]
  assign _GEN_70 = _T_610 ? {{1'd0}, _T_1375} : _T_337; // @[CSR.scala 277:29:@5741.6]
  assign _T_1376 = _T_336[39:32]; // @[CSR.scala 278:45:@5748.8]
  assign _T_1377 = {_T_1376,wdata}; // @[Cat.scala 30:58:@5749.8]
  assign _GEN_71 = _T_608 ? {{1'd0}, _T_1377} : _GEN_70; // @[CSR.scala 278:29:@5747.6]
  assign _T_1379 = _T_339[31:0]; // @[CSR.scala 277:72:@5754.8]
  assign _T_1380 = {_T_1253,_T_1379}; // @[Cat.scala 30:58:@5755.8]
  assign _GEN_72 = _T_614 ? {{1'd0}, _T_1380} : _T_340; // @[CSR.scala 277:29:@5752.6]
  assign _T_1381 = _T_339[39:32]; // @[CSR.scala 278:45:@5759.8]
  assign _T_1382 = {_T_1381,wdata}; // @[Cat.scala 30:58:@5760.8]
  assign _GEN_73 = _T_612 ? {{1'd0}, _T_1382} : _GEN_72; // @[CSR.scala 278:29:@5758.6]
  assign _T_1384 = _T_342[31:0]; // @[CSR.scala 277:72:@5765.8]
  assign _T_1385 = {_T_1253,_T_1384}; // @[Cat.scala 30:58:@5766.8]
  assign _GEN_74 = _T_618 ? {{1'd0}, _T_1385} : _T_343; // @[CSR.scala 277:29:@5763.6]
  assign _T_1386 = _T_342[39:32]; // @[CSR.scala 278:45:@5770.8]
  assign _T_1387 = {_T_1386,wdata}; // @[Cat.scala 30:58:@5771.8]
  assign _GEN_75 = _T_616 ? {{1'd0}, _T_1387} : _GEN_74; // @[CSR.scala 278:29:@5769.6]
  assign _T_1389 = _T_345[31:0]; // @[CSR.scala 277:72:@5776.8]
  assign _T_1390 = {_T_1253,_T_1389}; // @[Cat.scala 30:58:@5777.8]
  assign _GEN_76 = _T_622 ? {{1'd0}, _T_1390} : _T_346; // @[CSR.scala 277:29:@5774.6]
  assign _T_1391 = _T_345[39:32]; // @[CSR.scala 278:45:@5781.8]
  assign _T_1392 = {_T_1391,wdata}; // @[Cat.scala 30:58:@5782.8]
  assign _GEN_77 = _T_620 ? {{1'd0}, _T_1392} : _GEN_76; // @[CSR.scala 278:29:@5780.6]
  assign _T_1394 = _T_348[31:0]; // @[CSR.scala 277:72:@5787.8]
  assign _T_1395 = {_T_1253,_T_1394}; // @[Cat.scala 30:58:@5788.8]
  assign _GEN_78 = _T_626 ? {{1'd0}, _T_1395} : _T_349; // @[CSR.scala 277:29:@5785.6]
  assign _T_1396 = _T_348[39:32]; // @[CSR.scala 278:45:@5792.8]
  assign _T_1397 = {_T_1396,wdata}; // @[Cat.scala 30:58:@5793.8]
  assign _GEN_79 = _T_624 ? {{1'd0}, _T_1397} : _GEN_78; // @[CSR.scala 278:29:@5791.6]
  assign _T_1399 = _T_351[31:0]; // @[CSR.scala 277:72:@5798.8]
  assign _T_1400 = {_T_1253,_T_1399}; // @[Cat.scala 30:58:@5799.8]
  assign _GEN_80 = _T_630 ? {{1'd0}, _T_1400} : _T_352; // @[CSR.scala 277:29:@5796.6]
  assign _T_1401 = _T_351[39:32]; // @[CSR.scala 278:45:@5803.8]
  assign _T_1402 = {_T_1401,wdata}; // @[Cat.scala 30:58:@5804.8]
  assign _GEN_81 = _T_628 ? {{1'd0}, _T_1402} : _GEN_80; // @[CSR.scala 278:29:@5802.6]
  assign _T_1404 = _T_354[31:0]; // @[CSR.scala 277:72:@5809.8]
  assign _T_1405 = {_T_1253,_T_1404}; // @[Cat.scala 30:58:@5810.8]
  assign _GEN_82 = _T_634 ? {{1'd0}, _T_1405} : _T_355; // @[CSR.scala 277:29:@5807.6]
  assign _T_1406 = _T_354[39:32]; // @[CSR.scala 278:45:@5814.8]
  assign _T_1407 = {_T_1406,wdata}; // @[Cat.scala 30:58:@5815.8]
  assign _GEN_83 = _T_632 ? {{1'd0}, _T_1407} : _GEN_82; // @[CSR.scala 278:29:@5813.6]
  assign _T_1409 = _T_357[31:0]; // @[CSR.scala 277:72:@5820.8]
  assign _T_1410 = {_T_1253,_T_1409}; // @[Cat.scala 30:58:@5821.8]
  assign _GEN_84 = _T_638 ? {{1'd0}, _T_1410} : _T_358; // @[CSR.scala 277:29:@5818.6]
  assign _T_1411 = _T_357[39:32]; // @[CSR.scala 278:45:@5825.8]
  assign _T_1412 = {_T_1411,wdata}; // @[Cat.scala 30:58:@5826.8]
  assign _GEN_85 = _T_636 ? {{1'd0}, _T_1412} : _GEN_84; // @[CSR.scala 278:29:@5824.6]
  assign _T_1414 = _T_249[31:0]; // @[CSR.scala 277:72:@5831.8]
  assign _T_1415 = {wdata,_T_1414}; // @[Cat.scala 30:58:@5832.8]
  assign _T_1416 = _T_1415[63:6]; // @[Util.scala 133:28:@5834.8]
  assign _GEN_86 = _T_640 ? _T_1415 : {{57'd0}, _T_241}; // @[CSR.scala 277:29:@5829.6]
  assign _GEN_87 = _T_640 ? _T_1416 : _GEN_0; // @[CSR.scala 277:29:@5829.6]
  assign _T_1417 = _T_249[63:32]; // @[CSR.scala 278:45:@5838.8]
  assign _T_1418 = {_T_1417,wdata}; // @[Cat.scala 30:58:@5839.8]
  assign _T_1419 = _T_1418[63:6]; // @[Util.scala 133:28:@5841.8]
  assign _GEN_88 = _T_478 ? _T_1418 : _GEN_86; // @[CSR.scala 278:29:@5837.6]
  assign _GEN_89 = _T_478 ? _T_1419 : _GEN_87; // @[CSR.scala 278:29:@5837.6]
  assign _T_1421 = _T_261[31:0]; // @[CSR.scala 277:72:@5846.8]
  assign _T_1422 = {wdata,_T_1421}; // @[Cat.scala 30:58:@5847.8]
  assign _T_1423 = _T_1422[63:6]; // @[Util.scala 133:28:@5849.8]
  assign _GEN_90 = _T_642 ? _T_1422 : {{57'd0}, _T_253}; // @[CSR.scala 277:29:@5844.6]
  assign _GEN_91 = _T_642 ? _T_1423 : _GEN_1; // @[CSR.scala 277:29:@5844.6]
  assign _T_1424 = _T_261[63:32]; // @[CSR.scala 278:45:@5853.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:@5854.8]
  assign _T_1426 = _T_1425[63:6]; // @[Util.scala 133:28:@5856.8]
  assign _GEN_92 = _T_480 ? _T_1425 : _GEN_90; // @[CSR.scala 278:29:@5852.6]
  assign _GEN_93 = _T_480 ? _T_1426 : _GEN_91; // @[CSR.scala 278:29:@5852.6]
  assign _GEN_94 = _T_508 ? wdata : reg_dscratch; // @[CSR.scala 265:40:@5859.6]
  assign _T_1429 = wdata >> 2'h2; // @[CSR.scala 267:78:@5864.8]
  assign _GEN_225 = {{3'd0}, _T_1429}; // @[CSR.scala 267:86:@5865.8]
  assign _T_1431 = _GEN_225 << 2'h2; // @[CSR.scala 267:86:@5865.8]
  assign _GEN_95 = _T_500 ? _T_1431 : {{3'd0}, _GEN_15}; // @[CSR.scala 267:40:@5862.6]
  assign _GEN_96 = _T_498 ? wdata : reg_mscratch; // @[CSR.scala 268:40:@5868.6]
  assign _T_1433 = wdata & 32'h8000001f; // @[CSR.scala 269:62:@5872.8]
  assign _GEN_97 = _T_504 ? _T_1433 : _GEN_14; // @[CSR.scala 269:40:@5871.6]
  assign _GEN_98 = _T_502 ? wdata : _GEN_16; // @[CSR.scala 270:40:@5875.6]
  assign _GEN_99 = _T_510 ? wdata : reg_medeleg; // @[CSR.scala 271:42:@5879.6]
  assign _GEN_100 = wen ? _GEN_17 : _GEN_3; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_101 = wen ? _GEN_18 : _GEN_4; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_102 = wen ? _GEN_19 : reg_mip_msip; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_103 = wen ? _GEN_20 : reg_mie_msip; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_104 = wen ? _GEN_21 : reg_mie_mtip; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_105 = wen ? _GEN_23 : _T_265; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_106 = wen ? _GEN_25 : _T_268; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_107 = wen ? _GEN_27 : _T_271; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_108 = wen ? _GEN_29 : _T_274; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_109 = wen ? _GEN_31 : _T_277; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_110 = wen ? _GEN_33 : _T_280; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_111 = wen ? _GEN_35 : _T_283; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_112 = wen ? _GEN_37 : _T_286; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_113 = wen ? _GEN_39 : _T_289; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_114 = wen ? _GEN_41 : _T_292; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_115 = wen ? _GEN_43 : _T_295; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_116 = wen ? _GEN_45 : _T_298; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_117 = wen ? _GEN_47 : _T_301; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_118 = wen ? _GEN_49 : _T_304; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_119 = wen ? _GEN_51 : _T_307; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_120 = wen ? _GEN_53 : _T_310; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_121 = wen ? _GEN_55 : _T_313; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_122 = wen ? _GEN_57 : _T_316; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_123 = wen ? _GEN_59 : _T_319; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_124 = wen ? _GEN_61 : _T_322; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_125 = wen ? _GEN_63 : _T_325; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_126 = wen ? _GEN_65 : _T_328; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_127 = wen ? _GEN_67 : _T_331; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_128 = wen ? _GEN_69 : _T_334; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_129 = wen ? _GEN_71 : _T_337; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_130 = wen ? _GEN_73 : _T_340; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_131 = wen ? _GEN_75 : _T_343; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_132 = wen ? _GEN_77 : _T_346; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_133 = wen ? _GEN_79 : _T_349; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_134 = wen ? _GEN_81 : _T_352; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_135 = wen ? _GEN_83 : _T_355; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_136 = wen ? _GEN_85 : _T_358; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_137 = wen ? _GEN_88 : {{57'd0}, _T_241}; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_138 = wen ? _GEN_89 : _GEN_0; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_139 = wen ? _GEN_92 : {{57'd0}, _T_253}; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_140 = wen ? _GEN_93 : _GEN_1; // @[CSR.scala 242:14:@5408.4]
  assign _GEN_142 = wen ? _GEN_95 : {{3'd0}, _GEN_15}; // @[CSR.scala 242:14:@5408.4]
  assign io_rw_rdata = _T_1209[31:0]; // @[CSR.scala 240:15:@5407.4]
  assign io_eret = _T_940 | insn_ret; // @[CSR.scala 199:11:@5197.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 197:13:@5194.4]
  assign io_status_unimp5 = 14'h0; // @[CSR.scala 197:13:@5193.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 197:13:@5192.4]
  assign io_status_unimp4 = 2'h0; // @[CSR.scala 197:13:@5191.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 197:13:@5190.4]
  assign io_status_unimp3 = 3'h0; // @[CSR.scala 197:13:@5189.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 197:13:@5188.4]
  assign io_status_unimp2 = 3'h0; // @[CSR.scala 197:13:@5187.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 197:13:@5186.4]
  assign io_status_unimp1 = 3'h0; // @[CSR.scala 197:13:@5185.4]
  assign io_evec = io_xcpt ? 32'h80000004 : _GEN_10; // @[CSR.scala 212:13:@5218.6 CSR.scala 217:13:@5221.6 CSR.scala 224:13:@5228.6 CSR.scala 230:13:@5233.6]
  assign io_time = _T_249[31:0]; // @[CSR.scala 236:11:@5238.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_240 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_244 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_252 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_256 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_264 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_267 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_270 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_273 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_276 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_279 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_282 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_285 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_288 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_291 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_294 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_297 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_300 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_303 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_306 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_309 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_312 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_315 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_318 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_321 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_324 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_327 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_330 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_333 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_336 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_339 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_342 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_345 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_348 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_351 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_354 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_357 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_954) begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mpie <= _T_1222;
        end else begin
          if (_T_954) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mpie <= 1'h1;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mie <= _T_1220;
        end else begin
          if (_T_954) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end
    end
    reg_mepc <= _GEN_142[31:0];
    if (wen) begin
      if (_T_504) begin
        reg_mcause <= _T_1433;
      end else begin
        if (io_xcpt) begin
          reg_mcause <= io_cause;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_959};
            end
          end
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mcause <= io_cause;
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_959};
          end
        end
      end
    end
    if (wen) begin
      if (_T_502) begin
        reg_mtval <= wdata;
      end else begin
        if (io_xcpt) begin
          reg_mtval <= io_tval;
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mtval <= io_tval;
      end
    end
    if (wen) begin
      if (_T_498) begin
        reg_mscratch <= wdata;
      end
    end
    if (wen) begin
      if (_T_510) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (reset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_494) begin
          reg_mip_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_mtip <= _T_1237;
        end
      end
    end
    if (reset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      _T_240 <= 6'h0;
    end else begin
      _T_240 <= _GEN_137[5:0];
    end
    if (reset) begin
      _T_244 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_478) begin
          _T_244 <= _T_1419;
        end else begin
          if (_T_640) begin
            _T_244 <= _T_1416;
          end else begin
            if (_T_245) begin
              _T_244 <= _T_248;
            end
          end
        end
      end else begin
        if (_T_245) begin
          _T_244 <= _T_248;
        end
      end
    end
    if (reset) begin
      _T_252 <= 6'h0;
    end else begin
      _T_252 <= _GEN_139[5:0];
    end
    if (reset) begin
      _T_256 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_480) begin
          _T_256 <= _T_1426;
        end else begin
          if (_T_642) begin
            _T_256 <= _T_1423;
          end else begin
            if (_T_257) begin
              _T_256 <= _T_260;
            end
          end
        end
      end else begin
        if (_T_257) begin
          _T_256 <= _T_260;
        end
      end
    end
    _T_264 <= _GEN_105[39:0];
    _T_267 <= _GEN_106[39:0];
    _T_270 <= _GEN_107[39:0];
    _T_273 <= _GEN_108[39:0];
    _T_276 <= _GEN_109[39:0];
    _T_279 <= _GEN_110[39:0];
    _T_282 <= _GEN_111[39:0];
    _T_285 <= _GEN_112[39:0];
    _T_288 <= _GEN_113[39:0];
    _T_291 <= _GEN_114[39:0];
    _T_294 <= _GEN_115[39:0];
    _T_297 <= _GEN_116[39:0];
    _T_300 <= _GEN_117[39:0];
    _T_303 <= _GEN_118[39:0];
    _T_306 <= _GEN_119[39:0];
    _T_309 <= _GEN_120[39:0];
    _T_312 <= _GEN_121[39:0];
    _T_315 <= _GEN_122[39:0];
    _T_318 <= _GEN_123[39:0];
    _T_321 <= _GEN_124[39:0];
    _T_324 <= _GEN_125[39:0];
    _T_327 <= _GEN_126[39:0];
    _T_330 <= _GEN_127[39:0];
    _T_333 <= _GEN_128[39:0];
    _T_336 <= _GEN_129[39:0];
    _T_339 <= _GEN_130[39:0];
    _T_342 <= _GEN_131[39:0];
    _T_345 <= _GEN_132[39:0];
    _T_348 <= _GEN_133[39:0];
    _T_351 <= _GEN_134[39:0];
    _T_354 <= _GEN_135[39:0];
    _T_357 <= _GEN_136[39:0];
    if (wen) begin
      if (_T_508) begin
        reg_dscratch <= wdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:201 assert(PopCount(insn_ret :: io.illegal :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 201:9:@5204.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[CSR.scala 201:9:@5205.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module Regfile( // @[:@5885.2]
  input         clock, // @[:@5886.4]
  input  [4:0]  io_rs1_addr_0, // @[:@5888.4]
  input  [4:0]  io_rs1_addr_1, // @[:@5888.4]
  output [31:0] io_rs1_data_0, // @[:@5888.4]
  output [31:0] io_rs1_data_1, // @[:@5888.4]
  input  [4:0]  io_rs2_addr_0, // @[:@5888.4]
  input  [4:0]  io_rs2_addr_1, // @[:@5888.4]
  output [31:0] io_rs2_data_0, // @[:@5888.4]
  output [31:0] io_rs2_data_1, // @[:@5888.4]
  input  [4:0]  io_waddr_0, // @[:@5888.4]
  input  [4:0]  io_waddr_1, // @[:@5888.4]
  input  [31:0] io_wdata_0, // @[:@5888.4]
  input  [31:0] io_wdata_1, // @[:@5888.4]
  input         io_wen_0, // @[:@5888.4]
  input         io_wen_1 // @[:@5888.4]
);
  reg [31:0] regfile [0:31]; // @[Regfile.scala 23:20:@5890.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_109_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_109_addr; // @[Regfile.scala 23:20:@5890.4]
  wire [31:0] regfile__T_114_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_114_addr; // @[Regfile.scala 23:20:@5890.4]
  wire [31:0] regfile__T_119_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_119_addr; // @[Regfile.scala 23:20:@5890.4]
  wire [31:0] regfile__T_124_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_124_addr; // @[Regfile.scala 23:20:@5890.4]
  wire [31:0] regfile__T_105_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_105_addr; // @[Regfile.scala 23:20:@5890.4]
  wire  regfile__T_105_mask; // @[Regfile.scala 23:20:@5890.4]
  wire  regfile__T_105_en; // @[Regfile.scala 23:20:@5890.4]
  wire [31:0] regfile__T_106_data; // @[Regfile.scala 23:20:@5890.4]
  wire [4:0] regfile__T_106_addr; // @[Regfile.scala 23:20:@5890.4]
  wire  regfile__T_106_mask; // @[Regfile.scala 23:20:@5890.4]
  wire  regfile__T_106_en; // @[Regfile.scala 23:20:@5890.4]
  wire  _T_108; // @[Regfile.scala 28:42:@5899.4]
  wire  _T_113; // @[Regfile.scala 29:42:@5903.4]
  wire  _T_118; // @[Regfile.scala 28:42:@5907.4]
  wire  _T_123; // @[Regfile.scala 29:42:@5911.4]
  assign regfile__T_109_addr = io_rs1_addr_0;
  assign regfile__T_109_data = regfile[regfile__T_109_addr]; // @[Regfile.scala 23:20:@5890.4]
  assign regfile__T_114_addr = io_rs2_addr_0;
  assign regfile__T_114_data = regfile[regfile__T_114_addr]; // @[Regfile.scala 23:20:@5890.4]
  assign regfile__T_119_addr = io_rs1_addr_1;
  assign regfile__T_119_data = regfile[regfile__T_119_addr]; // @[Regfile.scala 23:20:@5890.4]
  assign regfile__T_124_addr = io_rs2_addr_1;
  assign regfile__T_124_data = regfile[regfile__T_124_addr]; // @[Regfile.scala 23:20:@5890.4]
  assign regfile__T_105_data = io_wdata_0;
  assign regfile__T_105_addr = io_waddr_0;
  assign regfile__T_105_mask = 1'h1;
  assign regfile__T_105_en = io_wen_0;
  assign regfile__T_106_data = io_wdata_1;
  assign regfile__T_106_addr = io_waddr_1;
  assign regfile__T_106_mask = 1'h1;
  assign regfile__T_106_en = io_wen_1;
  assign _T_108 = io_rs1_addr_0 != 5'h0; // @[Regfile.scala 28:42:@5899.4]
  assign _T_113 = io_rs2_addr_0 != 5'h0; // @[Regfile.scala 29:42:@5903.4]
  assign _T_118 = io_rs1_addr_1 != 5'h0; // @[Regfile.scala 28:42:@5907.4]
  assign _T_123 = io_rs2_addr_1 != 5'h0; // @[Regfile.scala 29:42:@5911.4]
  assign io_rs1_data_0 = _T_108 ? regfile__T_109_data : 32'h0; // @[Regfile.scala 28:20:@5902.4]
  assign io_rs1_data_1 = _T_118 ? regfile__T_119_data : 32'h0; // @[Regfile.scala 28:20:@5910.4]
  assign io_rs2_data_0 = _T_113 ? regfile__T_114_data : 32'h0; // @[Regfile.scala 29:20:@5906.4]
  assign io_rs2_data_1 = _T_123 ? regfile__T_124_data : 32'h0; // @[Regfile.scala 29:20:@5914.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(regfile__T_105_en & regfile__T_105_mask) begin
      regfile[regfile__T_105_addr] <= regfile__T_105_data; // @[Regfile.scala 23:20:@5890.4]
    end
    if(regfile__T_106_en & regfile__T_106_mask) begin
      regfile[regfile__T_106_addr] <= regfile__T_106_data; // @[Regfile.scala 23:20:@5890.4]
    end
  end
endmodule
module ALU( // @[:@5916.2]
  input  [31:0] io_op1, // @[:@5919.4]
  input  [31:0] io_op2, // @[:@5919.4]
  input  [31:0] io_pc, // @[:@5919.4]
  input  [3:0]  io_ctrl_fun, // @[:@5919.4]
  input  [3:0]  io_ctrl_br_type, // @[:@5919.4]
  input  [1:0]  io_ctrl_wb_sel, // @[:@5919.4]
  output [1:0]  io_ctrl_pc_sel, // @[:@5919.4]
  input  [31:0] io_rs2_data, // @[:@5919.4]
  output [31:0] io_result, // @[:@5919.4]
  output [31:0] io_target_brjmp, // @[:@5919.4]
  output [31:0] io_target_jpreg, // @[:@5919.4]
  output [31:0] io_target_conti // @[:@5919.4]
);
  wire [4:0] alu_shamt; // @[ALU.scala 32:32:@5921.4]
  wire [32:0] _T_25; // @[ALU.scala 33:34:@5922.4]
  wire [31:0] add_result; // @[ALU.scala 33:34:@5923.4]
  wire  _T_29; // @[ALU.scala 38:18:@5926.4]
  wire  _T_30; // @[ALU.scala 39:18:@5927.4]
  wire [32:0] _T_31; // @[ALU.scala 39:44:@5928.4]
  wire [32:0] _T_32; // @[ALU.scala 39:44:@5929.4]
  wire [31:0] _T_33; // @[ALU.scala 39:44:@5930.4]
  wire  _T_34; // @[ALU.scala 40:18:@5931.4]
  wire [31:0] _T_35; // @[ALU.scala 40:44:@5932.4]
  wire  _T_36; // @[ALU.scala 41:18:@5933.4]
  wire [31:0] _T_37; // @[ALU.scala 41:44:@5934.4]
  wire  _T_38; // @[ALU.scala 42:18:@5935.4]
  wire [31:0] _T_39; // @[ALU.scala 42:44:@5936.4]
  wire  _T_40; // @[ALU.scala 43:18:@5937.4]
  wire [31:0] _T_41; // @[ALU.scala 43:44:@5938.4]
  wire [31:0] _T_42; // @[ALU.scala 43:60:@5939.4]
  wire  _T_43; // @[ALU.scala 43:51:@5940.4]
  wire  _T_44; // @[ALU.scala 44:18:@5941.4]
  wire  _T_45; // @[ALU.scala 44:44:@5942.4]
  wire  _T_46; // @[ALU.scala 45:18:@5943.4]
  wire [62:0] _GEN_0; // @[ALU.scala 45:44:@5944.4]
  wire [62:0] _T_47; // @[ALU.scala 45:44:@5944.4]
  wire [31:0] _T_48; // @[ALU.scala 45:57:@5945.4]
  wire  _T_49; // @[ALU.scala 46:18:@5946.4]
  wire [31:0] _T_51; // @[ALU.scala 46:51:@5948.4]
  wire [31:0] _T_52; // @[ALU.scala 46:65:@5949.4]
  wire  _T_53; // @[ALU.scala 47:18:@5950.4]
  wire [31:0] _T_54; // @[ALU.scala 47:44:@5951.4]
  wire  _T_55; // @[ALU.scala 48:18:@5952.4]
  wire  _T_56; // @[ALU.scala 49:18:@5953.4]
  wire [31:0] _T_57; // @[Mux.scala 61:16:@5954.4]
  wire [31:0] _T_58; // @[Mux.scala 61:16:@5955.4]
  wire [31:0] _T_59; // @[Mux.scala 61:16:@5956.4]
  wire [31:0] _T_60; // @[Mux.scala 61:16:@5957.4]
  wire [31:0] _T_61; // @[Mux.scala 61:16:@5958.4]
  wire [31:0] _T_62; // @[Mux.scala 61:16:@5959.4]
  wire [31:0] _T_63; // @[Mux.scala 61:16:@5960.4]
  wire [31:0] _T_64; // @[Mux.scala 61:16:@5961.4]
  wire [31:0] _T_65; // @[Mux.scala 61:16:@5962.4]
  wire [31:0] _T_66; // @[Mux.scala 61:16:@5963.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@5964.4]
  wire [31:0] result; // @[Mux.scala 61:16:@5965.4]
  wire [32:0] _T_69; // @[ALU.scala 52:31:@5967.4]
  wire [30:0] _T_71; // @[ALU.scala 53:39:@5970.4]
  wire [32:0] _T_75; // @[ALU.scala 54:31:@5973.4]
  wire  _T_77; // @[ALU.scala 55:35:@5976.4]
  wire  br_eq; // @[ALU.scala 57:29:@5979.4]
  wire [31:0] _T_80; // @[ALU.scala 58:50:@5981.4]
  wire  br_lt; // @[ALU.scala 58:36:@5982.4]
  wire  br_ltu; // @[ALU.scala 59:36:@5983.4]
  wire  _T_81; // @[ALU.scala 63:25:@5984.4]
  wire  _T_82; // @[ALU.scala 64:25:@5985.4]
  wire  _T_84; // @[ALU.scala 64:41:@5986.4]
  wire [1:0] _T_85; // @[ALU.scala 64:40:@5987.4]
  wire  _T_86; // @[ALU.scala 65:25:@5988.4]
  wire [1:0] _T_87; // @[ALU.scala 65:40:@5989.4]
  wire  _T_88; // @[ALU.scala 66:25:@5990.4]
  wire  _T_90; // @[ALU.scala 66:41:@5991.4]
  wire [1:0] _T_91; // @[ALU.scala 66:40:@5992.4]
  wire  _T_92; // @[ALU.scala 67:25:@5993.4]
  wire  _T_94; // @[ALU.scala 67:41:@5994.4]
  wire [1:0] _T_95; // @[ALU.scala 67:40:@5995.4]
  wire  _T_96; // @[ALU.scala 68:25:@5996.4]
  wire [1:0] _T_97; // @[ALU.scala 68:40:@5997.4]
  wire  _T_98; // @[ALU.scala 69:25:@5998.4]
  wire [1:0] _T_99; // @[ALU.scala 69:40:@5999.4]
  wire  _T_100; // @[ALU.scala 70:25:@6000.4]
  wire  _T_101; // @[ALU.scala 71:25:@6001.4]
  wire [1:0] _T_102; // @[ALU.scala 71:8:@6002.4]
  wire [1:0] _T_103; // @[ALU.scala 70:8:@6003.4]
  wire [1:0] _T_104; // @[ALU.scala 69:8:@6004.4]
  wire [1:0] _T_105; // @[ALU.scala 68:8:@6005.4]
  wire [1:0] _T_106; // @[ALU.scala 67:8:@6006.4]
  wire [1:0] _T_107; // @[ALU.scala 66:8:@6007.4]
  wire [1:0] _T_108; // @[ALU.scala 65:8:@6008.4]
  wire [1:0] _T_109; // @[ALU.scala 64:8:@6009.4]
  assign alu_shamt = io_op2[4:0]; // @[ALU.scala 32:32:@5921.4]
  assign _T_25 = io_op1 + io_op2; // @[ALU.scala 33:34:@5922.4]
  assign add_result = io_op1 + io_op2; // @[ALU.scala 33:34:@5923.4]
  assign _T_29 = io_ctrl_fun == 4'h0; // @[ALU.scala 38:18:@5926.4]
  assign _T_30 = io_ctrl_fun == 4'h1; // @[ALU.scala 39:18:@5927.4]
  assign _T_31 = io_op1 - io_op2; // @[ALU.scala 39:44:@5928.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 39:44:@5929.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 39:44:@5930.4]
  assign _T_34 = io_ctrl_fun == 4'h5; // @[ALU.scala 40:18:@5931.4]
  assign _T_35 = io_op1 & io_op2; // @[ALU.scala 40:44:@5932.4]
  assign _T_36 = io_ctrl_fun == 4'h6; // @[ALU.scala 41:18:@5933.4]
  assign _T_37 = io_op1 | io_op2; // @[ALU.scala 41:44:@5934.4]
  assign _T_38 = io_ctrl_fun == 4'h7; // @[ALU.scala 42:18:@5935.4]
  assign _T_39 = io_op1 ^ io_op2; // @[ALU.scala 42:44:@5936.4]
  assign _T_40 = io_ctrl_fun == 4'h8; // @[ALU.scala 43:18:@5937.4]
  assign _T_41 = $signed(io_op1); // @[ALU.scala 43:44:@5938.4]
  assign _T_42 = $signed(io_op2); // @[ALU.scala 43:60:@5939.4]
  assign _T_43 = $signed(_T_41) < $signed(_T_42); // @[ALU.scala 43:51:@5940.4]
  assign _T_44 = io_ctrl_fun == 4'h9; // @[ALU.scala 44:18:@5941.4]
  assign _T_45 = io_op1 < io_op2; // @[ALU.scala 44:44:@5942.4]
  assign _T_46 = io_ctrl_fun == 4'h2; // @[ALU.scala 45:18:@5943.4]
  assign _GEN_0 = {{31'd0}, io_op1}; // @[ALU.scala 45:44:@5944.4]
  assign _T_47 = _GEN_0 << alu_shamt; // @[ALU.scala 45:44:@5944.4]
  assign _T_48 = _T_47[31:0]; // @[ALU.scala 45:57:@5945.4]
  assign _T_49 = io_ctrl_fun == 4'h4; // @[ALU.scala 46:18:@5946.4]
  assign _T_51 = $signed(_T_41) >>> alu_shamt; // @[ALU.scala 46:51:@5948.4]
  assign _T_52 = $unsigned(_T_51); // @[ALU.scala 46:65:@5949.4]
  assign _T_53 = io_ctrl_fun == 4'h3; // @[ALU.scala 47:18:@5950.4]
  assign _T_54 = io_op1 >> alu_shamt; // @[ALU.scala 47:44:@5951.4]
  assign _T_55 = io_ctrl_fun == 4'ha; // @[ALU.scala 48:18:@5952.4]
  assign _T_56 = io_ctrl_fun == 4'hb; // @[ALU.scala 49:18:@5953.4]
  assign _T_57 = _T_56 ? io_op2 : 32'h0; // @[Mux.scala 61:16:@5954.4]
  assign _T_58 = _T_55 ? io_op1 : _T_57; // @[Mux.scala 61:16:@5955.4]
  assign _T_59 = _T_53 ? _T_54 : _T_58; // @[Mux.scala 61:16:@5956.4]
  assign _T_60 = _T_49 ? _T_52 : _T_59; // @[Mux.scala 61:16:@5957.4]
  assign _T_61 = _T_46 ? _T_48 : _T_60; // @[Mux.scala 61:16:@5958.4]
  assign _T_62 = _T_44 ? {{31'd0}, _T_45} : _T_61; // @[Mux.scala 61:16:@5959.4]
  assign _T_63 = _T_40 ? {{31'd0}, _T_43} : _T_62; // @[Mux.scala 61:16:@5960.4]
  assign _T_64 = _T_38 ? _T_39 : _T_63; // @[Mux.scala 61:16:@5961.4]
  assign _T_65 = _T_36 ? _T_37 : _T_64; // @[Mux.scala 61:16:@5962.4]
  assign _T_66 = _T_34 ? _T_35 : _T_65; // @[Mux.scala 61:16:@5963.4]
  assign _T_67 = _T_30 ? _T_33 : _T_66; // @[Mux.scala 61:16:@5964.4]
  assign result = _T_29 ? add_result : _T_67; // @[Mux.scala 61:16:@5965.4]
  assign _T_69 = io_pc + io_op2; // @[ALU.scala 52:31:@5967.4]
  assign _T_71 = add_result[31:1]; // @[ALU.scala 53:39:@5970.4]
  assign _T_75 = io_pc + 32'h4; // @[ALU.scala 54:31:@5973.4]
  assign _T_77 = io_ctrl_wb_sel == 2'h2; // @[ALU.scala 55:35:@5976.4]
  assign br_eq = io_op1 == io_rs2_data; // @[ALU.scala 57:29:@5979.4]
  assign _T_80 = $signed(io_rs2_data); // @[ALU.scala 58:50:@5981.4]
  assign br_lt = $signed(_T_41) < $signed(_T_80); // @[ALU.scala 58:36:@5982.4]
  assign br_ltu = io_op1 < io_rs2_data; // @[ALU.scala 59:36:@5983.4]
  assign _T_81 = io_ctrl_br_type == 4'h0; // @[ALU.scala 63:25:@5984.4]
  assign _T_82 = io_ctrl_br_type == 4'h1; // @[ALU.scala 64:25:@5985.4]
  assign _T_84 = br_eq == 1'h0; // @[ALU.scala 64:41:@5986.4]
  assign _T_85 = _T_84 ? 2'h1 : 2'h0; // @[ALU.scala 64:40:@5987.4]
  assign _T_86 = io_ctrl_br_type == 4'h2; // @[ALU.scala 65:25:@5988.4]
  assign _T_87 = br_eq ? 2'h1 : 2'h0; // @[ALU.scala 65:40:@5989.4]
  assign _T_88 = io_ctrl_br_type == 4'h3; // @[ALU.scala 66:25:@5990.4]
  assign _T_90 = br_lt == 1'h0; // @[ALU.scala 66:41:@5991.4]
  assign _T_91 = _T_90 ? 2'h1 : 2'h0; // @[ALU.scala 66:40:@5992.4]
  assign _T_92 = io_ctrl_br_type == 4'h4; // @[ALU.scala 67:25:@5993.4]
  assign _T_94 = br_ltu == 1'h0; // @[ALU.scala 67:41:@5994.4]
  assign _T_95 = _T_94 ? 2'h1 : 2'h0; // @[ALU.scala 67:40:@5995.4]
  assign _T_96 = io_ctrl_br_type == 4'h5; // @[ALU.scala 68:25:@5996.4]
  assign _T_97 = br_lt ? 2'h1 : 2'h0; // @[ALU.scala 68:40:@5997.4]
  assign _T_98 = io_ctrl_br_type == 4'h6; // @[ALU.scala 69:25:@5998.4]
  assign _T_99 = br_ltu ? 2'h1 : 2'h0; // @[ALU.scala 69:40:@5999.4]
  assign _T_100 = io_ctrl_br_type == 4'h7; // @[ALU.scala 70:25:@6000.4]
  assign _T_101 = io_ctrl_br_type == 4'h8; // @[ALU.scala 71:25:@6001.4]
  assign _T_102 = _T_101 ? 2'h2 : 2'h0; // @[ALU.scala 71:8:@6002.4]
  assign _T_103 = _T_100 ? 2'h1 : _T_102; // @[ALU.scala 70:8:@6003.4]
  assign _T_104 = _T_98 ? _T_99 : _T_103; // @[ALU.scala 69:8:@6004.4]
  assign _T_105 = _T_96 ? _T_97 : _T_104; // @[ALU.scala 68:8:@6005.4]
  assign _T_106 = _T_92 ? _T_95 : _T_105; // @[ALU.scala 67:8:@6006.4]
  assign _T_107 = _T_88 ? _T_91 : _T_106; // @[ALU.scala 66:8:@6007.4]
  assign _T_108 = _T_86 ? _T_87 : _T_107; // @[ALU.scala 65:8:@6008.4]
  assign _T_109 = _T_82 ? _T_85 : _T_108; // @[ALU.scala 64:8:@6009.4]
  assign io_ctrl_pc_sel = _T_81 ? 2'h0 : _T_109; // @[ALU.scala 62:18:@6011.4]
  assign io_result = _T_77 ? io_target_conti : result; // @[ALU.scala 55:13:@5978.4]
  assign io_target_brjmp = io_pc + io_op2; // @[ALU.scala 52:22:@5969.4]
  assign io_target_jpreg = {_T_71,1'h0}; // @[ALU.scala 53:22:@5972.4]
  assign io_target_conti = io_pc + 32'h4; // @[ALU.scala 54:22:@5975.4]
endmodule
module InstDecoder( // @[:@6110.2]
  input  [31:0] io_inst, // @[:@6113.4]
  output [3:0]  io_cinfo_br_type, // @[:@6113.4]
  output [1:0]  io_cinfo_op1_sel, // @[:@6113.4]
  output [2:0]  io_cinfo_op2_sel, // @[:@6113.4]
  output        io_cinfo_rs1_oen, // @[:@6113.4]
  output        io_cinfo_rs2_oen, // @[:@6113.4]
  output [3:0]  io_cinfo_alu_fun, // @[:@6113.4]
  output [1:0]  io_cinfo_wb_sel, // @[:@6113.4]
  output        io_cinfo_rf_wen, // @[:@6113.4]
  output        io_cinfo_mem_en, // @[:@6113.4]
  output        io_cinfo_mem_fcn, // @[:@6113.4]
  output [2:0]  io_cinfo_mem_typ, // @[:@6113.4]
  output [2:0]  io_cinfo_csr_cmd, // @[:@6113.4]
  output        io_cinfo_illegal, // @[:@6113.4]
  output        io_cinfo_fencei, // @[:@6113.4]
  output        io_cinfo_branch, // @[:@6113.4]
  output        io_cinfo_push, // @[:@6113.4]
  output        io_cinfo_pop, // @[:@6113.4]
  output        io_cinfo_isBJ, // @[:@6113.4]
  output [4:0]  io_cinfo_rs1_addr, // @[:@6113.4]
  output [4:0]  io_cinfo_rs2_addr, // @[:@6113.4]
  output [4:0]  io_cinfo_wbaddr, // @[:@6113.4]
  output [31:0] io_dinfo_imm_i, // @[:@6113.4]
  output [31:0] io_dinfo_imm_s, // @[:@6113.4]
  output [31:0] io_dinfo_imm_sb, // @[:@6113.4]
  output [31:0] io_dinfo_imm_u, // @[:@6113.4]
  output [31:0] io_dinfo_imm_uj, // @[:@6113.4]
  output [31:0] io_dinfo_imm_z // @[:@6113.4]
);
  wire [31:0] _T_13; // @[Lookup.scala 9:38:@6115.4]
  wire  _T_14; // @[Lookup.scala 9:38:@6116.4]
  wire  _T_18; // @[Lookup.scala 9:38:@6118.4]
  wire  _T_22; // @[Lookup.scala 9:38:@6120.4]
  wire  _T_26; // @[Lookup.scala 9:38:@6122.4]
  wire  _T_30; // @[Lookup.scala 9:38:@6124.4]
  wire  _T_34; // @[Lookup.scala 9:38:@6126.4]
  wire  _T_38; // @[Lookup.scala 9:38:@6128.4]
  wire  _T_42; // @[Lookup.scala 9:38:@6130.4]
  wire [31:0] _T_45; // @[Lookup.scala 9:38:@6131.4]
  wire  _T_46; // @[Lookup.scala 9:38:@6132.4]
  wire  _T_50; // @[Lookup.scala 9:38:@6134.4]
  wire  _T_54; // @[Lookup.scala 9:38:@6136.4]
  wire  _T_58; // @[Lookup.scala 9:38:@6138.4]
  wire  _T_62; // @[Lookup.scala 9:38:@6140.4]
  wire  _T_66; // @[Lookup.scala 9:38:@6142.4]
  wire  _T_70; // @[Lookup.scala 9:38:@6144.4]
  wire  _T_74; // @[Lookup.scala 9:38:@6146.4]
  wire [31:0] _T_77; // @[Lookup.scala 9:38:@6147.4]
  wire  _T_78; // @[Lookup.scala 9:38:@6148.4]
  wire  _T_82; // @[Lookup.scala 9:38:@6150.4]
  wire  _T_86; // @[Lookup.scala 9:38:@6152.4]
  wire [31:0] _T_89; // @[Lookup.scala 9:38:@6153.4]
  wire  _T_90; // @[Lookup.scala 9:38:@6154.4]
  wire  _T_94; // @[Lookup.scala 9:38:@6156.4]
  wire  _T_98; // @[Lookup.scala 9:38:@6158.4]
  wire  _T_102; // @[Lookup.scala 9:38:@6160.4]
  wire  _T_106; // @[Lookup.scala 9:38:@6162.4]
  wire  _T_110; // @[Lookup.scala 9:38:@6164.4]
  wire  _T_114; // @[Lookup.scala 9:38:@6166.4]
  wire  _T_118; // @[Lookup.scala 9:38:@6168.4]
  wire  _T_122; // @[Lookup.scala 9:38:@6170.4]
  wire  _T_126; // @[Lookup.scala 9:38:@6172.4]
  wire  _T_130; // @[Lookup.scala 9:38:@6174.4]
  wire  _T_134; // @[Lookup.scala 9:38:@6176.4]
  wire  _T_138; // @[Lookup.scala 9:38:@6178.4]
  wire  _T_142; // @[Lookup.scala 9:38:@6180.4]
  wire  _T_146; // @[Lookup.scala 9:38:@6182.4]
  wire  _T_150; // @[Lookup.scala 9:38:@6184.4]
  wire  _T_154; // @[Lookup.scala 9:38:@6186.4]
  wire  _T_158; // @[Lookup.scala 9:38:@6188.4]
  wire  _T_162; // @[Lookup.scala 9:38:@6190.4]
  wire  _T_166; // @[Lookup.scala 9:38:@6192.4]
  wire  _T_170; // @[Lookup.scala 9:38:@6194.4]
  wire  _T_174; // @[Lookup.scala 9:38:@6196.4]
  wire  _T_178; // @[Lookup.scala 9:38:@6198.4]
  wire  _T_182; // @[Lookup.scala 9:38:@6200.4]
  wire  _T_186; // @[Lookup.scala 9:38:@6202.4]
  wire  _T_190; // @[Lookup.scala 9:38:@6204.4]
  wire  _T_194; // @[Lookup.scala 9:38:@6206.4]
  wire  _T_198; // @[Lookup.scala 9:38:@6208.4]
  wire  _T_202; // @[Lookup.scala 9:38:@6210.4]
  wire  _T_206; // @[Lookup.scala 9:38:@6212.4]
  wire  _T_210; // @[Lookup.scala 9:38:@6214.4]
  wire  _T_212; // @[Lookup.scala 11:37:@6216.4]
  wire  _T_213; // @[Lookup.scala 11:37:@6217.4]
  wire  _T_214; // @[Lookup.scala 11:37:@6218.4]
  wire  _T_215; // @[Lookup.scala 11:37:@6219.4]
  wire  _T_216; // @[Lookup.scala 11:37:@6220.4]
  wire  _T_217; // @[Lookup.scala 11:37:@6221.4]
  wire  _T_218; // @[Lookup.scala 11:37:@6222.4]
  wire  _T_219; // @[Lookup.scala 11:37:@6223.4]
  wire  _T_220; // @[Lookup.scala 11:37:@6224.4]
  wire  _T_221; // @[Lookup.scala 11:37:@6225.4]
  wire  _T_222; // @[Lookup.scala 11:37:@6226.4]
  wire  _T_223; // @[Lookup.scala 11:37:@6227.4]
  wire  _T_224; // @[Lookup.scala 11:37:@6228.4]
  wire  _T_225; // @[Lookup.scala 11:37:@6229.4]
  wire  _T_226; // @[Lookup.scala 11:37:@6230.4]
  wire  _T_227; // @[Lookup.scala 11:37:@6231.4]
  wire  _T_228; // @[Lookup.scala 11:37:@6232.4]
  wire  _T_229; // @[Lookup.scala 11:37:@6233.4]
  wire  _T_230; // @[Lookup.scala 11:37:@6234.4]
  wire  _T_231; // @[Lookup.scala 11:37:@6235.4]
  wire  _T_232; // @[Lookup.scala 11:37:@6236.4]
  wire  _T_233; // @[Lookup.scala 11:37:@6237.4]
  wire  _T_234; // @[Lookup.scala 11:37:@6238.4]
  wire  _T_235; // @[Lookup.scala 11:37:@6239.4]
  wire  _T_236; // @[Lookup.scala 11:37:@6240.4]
  wire  _T_237; // @[Lookup.scala 11:37:@6241.4]
  wire  _T_238; // @[Lookup.scala 11:37:@6242.4]
  wire  _T_239; // @[Lookup.scala 11:37:@6243.4]
  wire  _T_240; // @[Lookup.scala 11:37:@6244.4]
  wire  _T_241; // @[Lookup.scala 11:37:@6245.4]
  wire  _T_242; // @[Lookup.scala 11:37:@6246.4]
  wire  _T_243; // @[Lookup.scala 11:37:@6247.4]
  wire  _T_244; // @[Lookup.scala 11:37:@6248.4]
  wire  _T_245; // @[Lookup.scala 11:37:@6249.4]
  wire  _T_246; // @[Lookup.scala 11:37:@6250.4]
  wire  _T_247; // @[Lookup.scala 11:37:@6251.4]
  wire  _T_248; // @[Lookup.scala 11:37:@6252.4]
  wire  _T_249; // @[Lookup.scala 11:37:@6253.4]
  wire  _T_250; // @[Lookup.scala 11:37:@6254.4]
  wire  _T_251; // @[Lookup.scala 11:37:@6255.4]
  wire  _T_252; // @[Lookup.scala 11:37:@6256.4]
  wire  _T_253; // @[Lookup.scala 11:37:@6257.4]
  wire  _T_254; // @[Lookup.scala 11:37:@6258.4]
  wire  _T_255; // @[Lookup.scala 11:37:@6259.4]
  wire  _T_256; // @[Lookup.scala 11:37:@6260.4]
  wire  _T_257; // @[Lookup.scala 11:37:@6261.4]
  wire  _T_258; // @[Lookup.scala 11:37:@6262.4]
  wire  _T_259; // @[Lookup.scala 11:37:@6263.4]
  wire  signals_0; // @[Lookup.scala 11:37:@6264.4]
  wire [3:0] _T_273; // @[Lookup.scala 11:37:@6278.4]
  wire [3:0] _T_274; // @[Lookup.scala 11:37:@6279.4]
  wire [3:0] _T_275; // @[Lookup.scala 11:37:@6280.4]
  wire [3:0] _T_276; // @[Lookup.scala 11:37:@6281.4]
  wire [3:0] _T_277; // @[Lookup.scala 11:37:@6282.4]
  wire [3:0] _T_278; // @[Lookup.scala 11:37:@6283.4]
  wire [3:0] _T_279; // @[Lookup.scala 11:37:@6284.4]
  wire [3:0] _T_280; // @[Lookup.scala 11:37:@6285.4]
  wire [3:0] _T_281; // @[Lookup.scala 11:37:@6286.4]
  wire [3:0] _T_282; // @[Lookup.scala 11:37:@6287.4]
  wire [3:0] _T_283; // @[Lookup.scala 11:37:@6288.4]
  wire [3:0] _T_284; // @[Lookup.scala 11:37:@6289.4]
  wire [3:0] _T_285; // @[Lookup.scala 11:37:@6290.4]
  wire [3:0] _T_286; // @[Lookup.scala 11:37:@6291.4]
  wire [3:0] _T_287; // @[Lookup.scala 11:37:@6292.4]
  wire [3:0] _T_288; // @[Lookup.scala 11:37:@6293.4]
  wire [3:0] _T_289; // @[Lookup.scala 11:37:@6294.4]
  wire [3:0] _T_290; // @[Lookup.scala 11:37:@6295.4]
  wire [3:0] _T_291; // @[Lookup.scala 11:37:@6296.4]
  wire [3:0] _T_292; // @[Lookup.scala 11:37:@6297.4]
  wire [3:0] _T_293; // @[Lookup.scala 11:37:@6298.4]
  wire [3:0] _T_294; // @[Lookup.scala 11:37:@6299.4]
  wire [3:0] _T_295; // @[Lookup.scala 11:37:@6300.4]
  wire [3:0] _T_296; // @[Lookup.scala 11:37:@6301.4]
  wire [3:0] _T_297; // @[Lookup.scala 11:37:@6302.4]
  wire [3:0] _T_298; // @[Lookup.scala 11:37:@6303.4]
  wire [3:0] _T_299; // @[Lookup.scala 11:37:@6304.4]
  wire [3:0] _T_300; // @[Lookup.scala 11:37:@6305.4]
  wire [3:0] _T_301; // @[Lookup.scala 11:37:@6306.4]
  wire [3:0] _T_302; // @[Lookup.scala 11:37:@6307.4]
  wire [3:0] _T_303; // @[Lookup.scala 11:37:@6308.4]
  wire [3:0] _T_304; // @[Lookup.scala 11:37:@6309.4]
  wire [3:0] _T_305; // @[Lookup.scala 11:37:@6310.4]
  wire [3:0] _T_306; // @[Lookup.scala 11:37:@6311.4]
  wire [3:0] _T_307; // @[Lookup.scala 11:37:@6312.4]
  wire [3:0] _T_308; // @[Lookup.scala 11:37:@6313.4]
  wire [1:0] _T_316; // @[Lookup.scala 11:37:@6322.4]
  wire [1:0] _T_317; // @[Lookup.scala 11:37:@6323.4]
  wire [1:0] _T_318; // @[Lookup.scala 11:37:@6324.4]
  wire [1:0] _T_319; // @[Lookup.scala 11:37:@6325.4]
  wire [1:0] _T_320; // @[Lookup.scala 11:37:@6326.4]
  wire [1:0] _T_321; // @[Lookup.scala 11:37:@6327.4]
  wire [1:0] _T_322; // @[Lookup.scala 11:37:@6328.4]
  wire [1:0] _T_323; // @[Lookup.scala 11:37:@6329.4]
  wire [1:0] _T_324; // @[Lookup.scala 11:37:@6330.4]
  wire [1:0] _T_325; // @[Lookup.scala 11:37:@6331.4]
  wire [1:0] _T_326; // @[Lookup.scala 11:37:@6332.4]
  wire [1:0] _T_327; // @[Lookup.scala 11:37:@6333.4]
  wire [1:0] _T_328; // @[Lookup.scala 11:37:@6334.4]
  wire [1:0] _T_329; // @[Lookup.scala 11:37:@6335.4]
  wire [1:0] _T_330; // @[Lookup.scala 11:37:@6336.4]
  wire [1:0] _T_331; // @[Lookup.scala 11:37:@6337.4]
  wire [1:0] _T_332; // @[Lookup.scala 11:37:@6338.4]
  wire [1:0] _T_333; // @[Lookup.scala 11:37:@6339.4]
  wire [1:0] _T_334; // @[Lookup.scala 11:37:@6340.4]
  wire [1:0] _T_335; // @[Lookup.scala 11:37:@6341.4]
  wire [1:0] _T_336; // @[Lookup.scala 11:37:@6342.4]
  wire [1:0] _T_337; // @[Lookup.scala 11:37:@6343.4]
  wire [1:0] _T_338; // @[Lookup.scala 11:37:@6344.4]
  wire [1:0] _T_339; // @[Lookup.scala 11:37:@6345.4]
  wire [1:0] _T_340; // @[Lookup.scala 11:37:@6346.4]
  wire [1:0] _T_341; // @[Lookup.scala 11:37:@6347.4]
  wire [1:0] _T_342; // @[Lookup.scala 11:37:@6348.4]
  wire [1:0] _T_343; // @[Lookup.scala 11:37:@6349.4]
  wire [1:0] _T_344; // @[Lookup.scala 11:37:@6350.4]
  wire [1:0] _T_345; // @[Lookup.scala 11:37:@6351.4]
  wire [1:0] _T_346; // @[Lookup.scala 11:37:@6352.4]
  wire [1:0] _T_347; // @[Lookup.scala 11:37:@6353.4]
  wire [1:0] _T_348; // @[Lookup.scala 11:37:@6354.4]
  wire [1:0] _T_349; // @[Lookup.scala 11:37:@6355.4]
  wire [1:0] _T_350; // @[Lookup.scala 11:37:@6356.4]
  wire [1:0] _T_351; // @[Lookup.scala 11:37:@6357.4]
  wire [1:0] _T_352; // @[Lookup.scala 11:37:@6358.4]
  wire [1:0] _T_353; // @[Lookup.scala 11:37:@6359.4]
  wire [1:0] _T_354; // @[Lookup.scala 11:37:@6360.4]
  wire [1:0] _T_355; // @[Lookup.scala 11:37:@6361.4]
  wire [1:0] _T_356; // @[Lookup.scala 11:37:@6362.4]
  wire [1:0] _T_357; // @[Lookup.scala 11:37:@6363.4]
  wire [2:0] _T_371; // @[Lookup.scala 11:37:@6378.4]
  wire [2:0] _T_372; // @[Lookup.scala 11:37:@6379.4]
  wire [2:0] _T_373; // @[Lookup.scala 11:37:@6380.4]
  wire [2:0] _T_374; // @[Lookup.scala 11:37:@6381.4]
  wire [2:0] _T_375; // @[Lookup.scala 11:37:@6382.4]
  wire [2:0] _T_376; // @[Lookup.scala 11:37:@6383.4]
  wire [2:0] _T_377; // @[Lookup.scala 11:37:@6384.4]
  wire [2:0] _T_378; // @[Lookup.scala 11:37:@6385.4]
  wire [2:0] _T_379; // @[Lookup.scala 11:37:@6386.4]
  wire [2:0] _T_380; // @[Lookup.scala 11:37:@6387.4]
  wire [2:0] _T_381; // @[Lookup.scala 11:37:@6388.4]
  wire [2:0] _T_382; // @[Lookup.scala 11:37:@6389.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@6390.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@6391.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@6392.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@6393.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@6394.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@6395.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@6396.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@6397.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@6398.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@6399.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@6400.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@6401.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@6402.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@6403.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@6404.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@6405.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@6406.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@6407.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@6408.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@6409.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@6410.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@6411.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@6412.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@6413.4]
  wire  _T_415; // @[Lookup.scala 11:37:@6423.4]
  wire  _T_416; // @[Lookup.scala 11:37:@6424.4]
  wire  _T_417; // @[Lookup.scala 11:37:@6425.4]
  wire  _T_418; // @[Lookup.scala 11:37:@6426.4]
  wire  _T_419; // @[Lookup.scala 11:37:@6427.4]
  wire  _T_420; // @[Lookup.scala 11:37:@6428.4]
  wire  _T_421; // @[Lookup.scala 11:37:@6429.4]
  wire  _T_422; // @[Lookup.scala 11:37:@6430.4]
  wire  _T_423; // @[Lookup.scala 11:37:@6431.4]
  wire  _T_424; // @[Lookup.scala 11:37:@6432.4]
  wire  _T_425; // @[Lookup.scala 11:37:@6433.4]
  wire  _T_426; // @[Lookup.scala 11:37:@6434.4]
  wire  _T_427; // @[Lookup.scala 11:37:@6435.4]
  wire  _T_428; // @[Lookup.scala 11:37:@6436.4]
  wire  _T_429; // @[Lookup.scala 11:37:@6437.4]
  wire  _T_430; // @[Lookup.scala 11:37:@6438.4]
  wire  _T_431; // @[Lookup.scala 11:37:@6439.4]
  wire  _T_432; // @[Lookup.scala 11:37:@6440.4]
  wire  _T_433; // @[Lookup.scala 11:37:@6441.4]
  wire  _T_434; // @[Lookup.scala 11:37:@6442.4]
  wire  _T_435; // @[Lookup.scala 11:37:@6443.4]
  wire  _T_436; // @[Lookup.scala 11:37:@6444.4]
  wire  _T_437; // @[Lookup.scala 11:37:@6445.4]
  wire  _T_438; // @[Lookup.scala 11:37:@6446.4]
  wire  _T_439; // @[Lookup.scala 11:37:@6447.4]
  wire  _T_440; // @[Lookup.scala 11:37:@6448.4]
  wire  _T_441; // @[Lookup.scala 11:37:@6449.4]
  wire  _T_442; // @[Lookup.scala 11:37:@6450.4]
  wire  _T_443; // @[Lookup.scala 11:37:@6451.4]
  wire  _T_444; // @[Lookup.scala 11:37:@6452.4]
  wire  _T_445; // @[Lookup.scala 11:37:@6453.4]
  wire  _T_446; // @[Lookup.scala 11:37:@6454.4]
  wire  _T_447; // @[Lookup.scala 11:37:@6455.4]
  wire  _T_448; // @[Lookup.scala 11:37:@6456.4]
  wire  _T_449; // @[Lookup.scala 11:37:@6457.4]
  wire  _T_450; // @[Lookup.scala 11:37:@6458.4]
  wire  _T_451; // @[Lookup.scala 11:37:@6459.4]
  wire  _T_452; // @[Lookup.scala 11:37:@6460.4]
  wire  _T_453; // @[Lookup.scala 11:37:@6461.4]
  wire  _T_454; // @[Lookup.scala 11:37:@6462.4]
  wire  _T_455; // @[Lookup.scala 11:37:@6463.4]
  wire  _T_475; // @[Lookup.scala 11:37:@6484.4]
  wire  _T_476; // @[Lookup.scala 11:37:@6485.4]
  wire  _T_477; // @[Lookup.scala 11:37:@6486.4]
  wire  _T_478; // @[Lookup.scala 11:37:@6487.4]
  wire  _T_479; // @[Lookup.scala 11:37:@6488.4]
  wire  _T_480; // @[Lookup.scala 11:37:@6489.4]
  wire  _T_481; // @[Lookup.scala 11:37:@6490.4]
  wire  _T_482; // @[Lookup.scala 11:37:@6491.4]
  wire  _T_483; // @[Lookup.scala 11:37:@6492.4]
  wire  _T_484; // @[Lookup.scala 11:37:@6493.4]
  wire  _T_485; // @[Lookup.scala 11:37:@6494.4]
  wire  _T_486; // @[Lookup.scala 11:37:@6495.4]
  wire  _T_487; // @[Lookup.scala 11:37:@6496.4]
  wire  _T_488; // @[Lookup.scala 11:37:@6497.4]
  wire  _T_489; // @[Lookup.scala 11:37:@6498.4]
  wire  _T_490; // @[Lookup.scala 11:37:@6499.4]
  wire  _T_491; // @[Lookup.scala 11:37:@6500.4]
  wire  _T_492; // @[Lookup.scala 11:37:@6501.4]
  wire  _T_493; // @[Lookup.scala 11:37:@6502.4]
  wire  _T_494; // @[Lookup.scala 11:37:@6503.4]
  wire  _T_495; // @[Lookup.scala 11:37:@6504.4]
  wire  _T_496; // @[Lookup.scala 11:37:@6505.4]
  wire  _T_497; // @[Lookup.scala 11:37:@6506.4]
  wire  _T_498; // @[Lookup.scala 11:37:@6507.4]
  wire  _T_499; // @[Lookup.scala 11:37:@6508.4]
  wire  _T_500; // @[Lookup.scala 11:37:@6509.4]
  wire  _T_501; // @[Lookup.scala 11:37:@6510.4]
  wire  _T_502; // @[Lookup.scala 11:37:@6511.4]
  wire  _T_503; // @[Lookup.scala 11:37:@6512.4]
  wire  _T_504; // @[Lookup.scala 11:37:@6513.4]
  wire [3:0] _T_512; // @[Lookup.scala 11:37:@6522.4]
  wire [3:0] _T_513; // @[Lookup.scala 11:37:@6523.4]
  wire [3:0] _T_514; // @[Lookup.scala 11:37:@6524.4]
  wire [3:0] _T_515; // @[Lookup.scala 11:37:@6525.4]
  wire [3:0] _T_516; // @[Lookup.scala 11:37:@6526.4]
  wire [3:0] _T_517; // @[Lookup.scala 11:37:@6527.4]
  wire [3:0] _T_518; // @[Lookup.scala 11:37:@6528.4]
  wire [3:0] _T_519; // @[Lookup.scala 11:37:@6529.4]
  wire [3:0] _T_520; // @[Lookup.scala 11:37:@6530.4]
  wire [3:0] _T_521; // @[Lookup.scala 11:37:@6531.4]
  wire [3:0] _T_522; // @[Lookup.scala 11:37:@6532.4]
  wire [3:0] _T_523; // @[Lookup.scala 11:37:@6533.4]
  wire [3:0] _T_524; // @[Lookup.scala 11:37:@6534.4]
  wire [3:0] _T_525; // @[Lookup.scala 11:37:@6535.4]
  wire [3:0] _T_526; // @[Lookup.scala 11:37:@6536.4]
  wire [3:0] _T_527; // @[Lookup.scala 11:37:@6537.4]
  wire [3:0] _T_528; // @[Lookup.scala 11:37:@6538.4]
  wire [3:0] _T_529; // @[Lookup.scala 11:37:@6539.4]
  wire [3:0] _T_530; // @[Lookup.scala 11:37:@6540.4]
  wire [3:0] _T_531; // @[Lookup.scala 11:37:@6541.4]
  wire [3:0] _T_532; // @[Lookup.scala 11:37:@6542.4]
  wire [3:0] _T_533; // @[Lookup.scala 11:37:@6543.4]
  wire [3:0] _T_534; // @[Lookup.scala 11:37:@6544.4]
  wire [3:0] _T_535; // @[Lookup.scala 11:37:@6545.4]
  wire [3:0] _T_536; // @[Lookup.scala 11:37:@6546.4]
  wire [3:0] _T_537; // @[Lookup.scala 11:37:@6547.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:@6548.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:@6549.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:@6550.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:@6551.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:@6552.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:@6553.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:@6554.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:@6555.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:@6556.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:@6557.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:@6558.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:@6559.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:@6560.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:@6561.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:@6562.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:@6563.4]
  wire [1:0] _T_561; // @[Lookup.scala 11:37:@6572.4]
  wire [1:0] _T_562; // @[Lookup.scala 11:37:@6573.4]
  wire [1:0] _T_563; // @[Lookup.scala 11:37:@6574.4]
  wire [1:0] _T_564; // @[Lookup.scala 11:37:@6575.4]
  wire [1:0] _T_565; // @[Lookup.scala 11:37:@6576.4]
  wire [1:0] _T_566; // @[Lookup.scala 11:37:@6577.4]
  wire [1:0] _T_567; // @[Lookup.scala 11:37:@6578.4]
  wire [1:0] _T_568; // @[Lookup.scala 11:37:@6579.4]
  wire [1:0] _T_569; // @[Lookup.scala 11:37:@6580.4]
  wire [1:0] _T_570; // @[Lookup.scala 11:37:@6581.4]
  wire [1:0] _T_571; // @[Lookup.scala 11:37:@6582.4]
  wire [1:0] _T_572; // @[Lookup.scala 11:37:@6583.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@6584.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@6585.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@6586.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@6587.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@6588.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@6589.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@6590.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@6591.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@6592.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@6593.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@6594.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@6595.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@6596.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@6597.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@6598.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@6599.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@6600.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@6601.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@6602.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@6603.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@6604.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@6605.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@6606.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@6607.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@6608.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@6609.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@6610.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@6611.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@6612.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@6613.4]
  wire  _T_616; // @[Lookup.scala 11:37:@6628.4]
  wire  _T_617; // @[Lookup.scala 11:37:@6629.4]
  wire  _T_618; // @[Lookup.scala 11:37:@6630.4]
  wire  _T_619; // @[Lookup.scala 11:37:@6631.4]
  wire  _T_620; // @[Lookup.scala 11:37:@6632.4]
  wire  _T_621; // @[Lookup.scala 11:37:@6633.4]
  wire  _T_622; // @[Lookup.scala 11:37:@6634.4]
  wire  _T_623; // @[Lookup.scala 11:37:@6635.4]
  wire  _T_624; // @[Lookup.scala 11:37:@6636.4]
  wire  _T_625; // @[Lookup.scala 11:37:@6637.4]
  wire  _T_626; // @[Lookup.scala 11:37:@6638.4]
  wire  _T_627; // @[Lookup.scala 11:37:@6639.4]
  wire  _T_628; // @[Lookup.scala 11:37:@6640.4]
  wire  _T_629; // @[Lookup.scala 11:37:@6641.4]
  wire  _T_630; // @[Lookup.scala 11:37:@6642.4]
  wire  _T_631; // @[Lookup.scala 11:37:@6643.4]
  wire  _T_632; // @[Lookup.scala 11:37:@6644.4]
  wire  _T_633; // @[Lookup.scala 11:37:@6645.4]
  wire  _T_634; // @[Lookup.scala 11:37:@6646.4]
  wire  _T_635; // @[Lookup.scala 11:37:@6647.4]
  wire  _T_636; // @[Lookup.scala 11:37:@6648.4]
  wire  _T_637; // @[Lookup.scala 11:37:@6649.4]
  wire  _T_638; // @[Lookup.scala 11:37:@6650.4]
  wire  _T_639; // @[Lookup.scala 11:37:@6651.4]
  wire  _T_640; // @[Lookup.scala 11:37:@6652.4]
  wire  _T_641; // @[Lookup.scala 11:37:@6653.4]
  wire  _T_642; // @[Lookup.scala 11:37:@6654.4]
  wire  _T_643; // @[Lookup.scala 11:37:@6655.4]
  wire  _T_644; // @[Lookup.scala 11:37:@6656.4]
  wire  _T_645; // @[Lookup.scala 11:37:@6657.4]
  wire  _T_646; // @[Lookup.scala 11:37:@6658.4]
  wire  _T_647; // @[Lookup.scala 11:37:@6659.4]
  wire  _T_648; // @[Lookup.scala 11:37:@6660.4]
  wire  _T_649; // @[Lookup.scala 11:37:@6661.4]
  wire  _T_650; // @[Lookup.scala 11:37:@6662.4]
  wire  _T_651; // @[Lookup.scala 11:37:@6663.4]
  wire  _T_653; // @[Lookup.scala 11:37:@6666.4]
  wire  _T_654; // @[Lookup.scala 11:37:@6667.4]
  wire  _T_655; // @[Lookup.scala 11:37:@6668.4]
  wire  _T_656; // @[Lookup.scala 11:37:@6669.4]
  wire  _T_657; // @[Lookup.scala 11:37:@6670.4]
  wire  _T_658; // @[Lookup.scala 11:37:@6671.4]
  wire  _T_659; // @[Lookup.scala 11:37:@6672.4]
  wire  _T_660; // @[Lookup.scala 11:37:@6673.4]
  wire  _T_661; // @[Lookup.scala 11:37:@6674.4]
  wire  _T_662; // @[Lookup.scala 11:37:@6675.4]
  wire  _T_663; // @[Lookup.scala 11:37:@6676.4]
  wire  _T_664; // @[Lookup.scala 11:37:@6677.4]
  wire  _T_665; // @[Lookup.scala 11:37:@6678.4]
  wire  _T_666; // @[Lookup.scala 11:37:@6679.4]
  wire  _T_667; // @[Lookup.scala 11:37:@6680.4]
  wire  _T_668; // @[Lookup.scala 11:37:@6681.4]
  wire  _T_669; // @[Lookup.scala 11:37:@6682.4]
  wire  _T_670; // @[Lookup.scala 11:37:@6683.4]
  wire  _T_671; // @[Lookup.scala 11:37:@6684.4]
  wire  _T_672; // @[Lookup.scala 11:37:@6685.4]
  wire  _T_673; // @[Lookup.scala 11:37:@6686.4]
  wire  _T_674; // @[Lookup.scala 11:37:@6687.4]
  wire  _T_675; // @[Lookup.scala 11:37:@6688.4]
  wire  _T_676; // @[Lookup.scala 11:37:@6689.4]
  wire  _T_677; // @[Lookup.scala 11:37:@6690.4]
  wire  _T_678; // @[Lookup.scala 11:37:@6691.4]
  wire  _T_679; // @[Lookup.scala 11:37:@6692.4]
  wire  _T_680; // @[Lookup.scala 11:37:@6693.4]
  wire  _T_681; // @[Lookup.scala 11:37:@6694.4]
  wire  _T_682; // @[Lookup.scala 11:37:@6695.4]
  wire  _T_683; // @[Lookup.scala 11:37:@6696.4]
  wire  _T_684; // @[Lookup.scala 11:37:@6697.4]
  wire  _T_685; // @[Lookup.scala 11:37:@6698.4]
  wire  _T_686; // @[Lookup.scala 11:37:@6699.4]
  wire  _T_687; // @[Lookup.scala 11:37:@6700.4]
  wire  _T_688; // @[Lookup.scala 11:37:@6701.4]
  wire  _T_689; // @[Lookup.scala 11:37:@6702.4]
  wire  _T_690; // @[Lookup.scala 11:37:@6703.4]
  wire  _T_691; // @[Lookup.scala 11:37:@6704.4]
  wire  _T_692; // @[Lookup.scala 11:37:@6705.4]
  wire  _T_693; // @[Lookup.scala 11:37:@6706.4]
  wire  _T_694; // @[Lookup.scala 11:37:@6707.4]
  wire  _T_695; // @[Lookup.scala 11:37:@6708.4]
  wire  _T_696; // @[Lookup.scala 11:37:@6709.4]
  wire  _T_697; // @[Lookup.scala 11:37:@6710.4]
  wire  _T_698; // @[Lookup.scala 11:37:@6711.4]
  wire  _T_699; // @[Lookup.scala 11:37:@6712.4]
  wire  _T_700; // @[Lookup.scala 11:37:@6713.4]
  wire  _T_744; // @[Lookup.scala 11:37:@6758.4]
  wire  _T_745; // @[Lookup.scala 11:37:@6759.4]
  wire  _T_746; // @[Lookup.scala 11:37:@6760.4]
  wire  _T_747; // @[Lookup.scala 11:37:@6761.4]
  wire  _T_748; // @[Lookup.scala 11:37:@6762.4]
  wire  _T_749; // @[Lookup.scala 11:37:@6763.4]
  wire [2:0] _T_792; // @[Lookup.scala 11:37:@6807.4]
  wire [2:0] _T_793; // @[Lookup.scala 11:37:@6808.4]
  wire [2:0] _T_794; // @[Lookup.scala 11:37:@6809.4]
  wire [2:0] _T_795; // @[Lookup.scala 11:37:@6810.4]
  wire [2:0] _T_796; // @[Lookup.scala 11:37:@6811.4]
  wire [2:0] _T_797; // @[Lookup.scala 11:37:@6812.4]
  wire [2:0] _T_798; // @[Lookup.scala 11:37:@6813.4]
  wire [2:0] _T_802; // @[Lookup.scala 11:37:@6818.4]
  wire [2:0] _T_803; // @[Lookup.scala 11:37:@6819.4]
  wire [2:0] _T_804; // @[Lookup.scala 11:37:@6820.4]
  wire [2:0] _T_805; // @[Lookup.scala 11:37:@6821.4]
  wire [2:0] _T_806; // @[Lookup.scala 11:37:@6822.4]
  wire [2:0] _T_807; // @[Lookup.scala 11:37:@6823.4]
  wire [2:0] _T_808; // @[Lookup.scala 11:37:@6824.4]
  wire [2:0] _T_809; // @[Lookup.scala 11:37:@6825.4]
  wire [2:0] _T_810; // @[Lookup.scala 11:37:@6826.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@6827.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@6828.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@6829.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@6830.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@6831.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@6832.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@6833.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@6834.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@6835.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@6836.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@6837.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@6838.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@6839.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@6840.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@6841.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@6842.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@6843.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@6844.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@6845.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@6846.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@6847.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@6848.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@6849.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@6850.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@6851.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@6852.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@6853.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@6854.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@6855.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@6856.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@6857.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@6858.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@6859.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@6860.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@6861.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@6862.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@6863.4]
  wire  _T_850; // @[Lookup.scala 11:37:@6867.4]
  wire  _T_851; // @[Lookup.scala 11:37:@6868.4]
  wire  _T_852; // @[Lookup.scala 11:37:@6869.4]
  wire  _T_853; // @[Lookup.scala 11:37:@6870.4]
  wire  _T_854; // @[Lookup.scala 11:37:@6871.4]
  wire  _T_855; // @[Lookup.scala 11:37:@6872.4]
  wire  _T_856; // @[Lookup.scala 11:37:@6873.4]
  wire  _T_857; // @[Lookup.scala 11:37:@6874.4]
  wire  _T_858; // @[Lookup.scala 11:37:@6875.4]
  wire  _T_859; // @[Lookup.scala 11:37:@6876.4]
  wire  _T_860; // @[Lookup.scala 11:37:@6877.4]
  wire  _T_861; // @[Lookup.scala 11:37:@6878.4]
  wire  _T_862; // @[Lookup.scala 11:37:@6879.4]
  wire  _T_863; // @[Lookup.scala 11:37:@6880.4]
  wire  _T_864; // @[Lookup.scala 11:37:@6881.4]
  wire  _T_865; // @[Lookup.scala 11:37:@6882.4]
  wire  _T_866; // @[Lookup.scala 11:37:@6883.4]
  wire  _T_867; // @[Lookup.scala 11:37:@6884.4]
  wire  _T_868; // @[Lookup.scala 11:37:@6885.4]
  wire  _T_869; // @[Lookup.scala 11:37:@6886.4]
  wire  _T_870; // @[Lookup.scala 11:37:@6887.4]
  wire  _T_871; // @[Lookup.scala 11:37:@6888.4]
  wire  _T_872; // @[Lookup.scala 11:37:@6889.4]
  wire  _T_873; // @[Lookup.scala 11:37:@6890.4]
  wire  _T_874; // @[Lookup.scala 11:37:@6891.4]
  wire  _T_875; // @[Lookup.scala 11:37:@6892.4]
  wire  _T_876; // @[Lookup.scala 11:37:@6893.4]
  wire  _T_877; // @[Lookup.scala 11:37:@6894.4]
  wire  _T_878; // @[Lookup.scala 11:37:@6895.4]
  wire  _T_879; // @[Lookup.scala 11:37:@6896.4]
  wire  _T_880; // @[Lookup.scala 11:37:@6897.4]
  wire  _T_881; // @[Lookup.scala 11:37:@6898.4]
  wire  _T_882; // @[Lookup.scala 11:37:@6899.4]
  wire  _T_883; // @[Lookup.scala 11:37:@6900.4]
  wire  _T_884; // @[Lookup.scala 11:37:@6901.4]
  wire  _T_885; // @[Lookup.scala 11:37:@6902.4]
  wire  _T_886; // @[Lookup.scala 11:37:@6903.4]
  wire  _T_887; // @[Lookup.scala 11:37:@6904.4]
  wire  _T_888; // @[Lookup.scala 11:37:@6905.4]
  wire  _T_889; // @[Lookup.scala 11:37:@6906.4]
  wire  _T_890; // @[Lookup.scala 11:37:@6907.4]
  wire  _T_891; // @[Lookup.scala 11:37:@6908.4]
  wire  _T_892; // @[Lookup.scala 11:37:@6909.4]
  wire  _T_893; // @[Lookup.scala 11:37:@6910.4]
  wire  _T_894; // @[Lookup.scala 11:37:@6911.4]
  wire  _T_895; // @[Lookup.scala 11:37:@6912.4]
  wire  _T_896; // @[Lookup.scala 11:37:@6913.4]
  wire [4:0] _T_899; // @[InstDecoder.scala 131:31:@6930.4]
  wire [4:0] _T_901; // @[InstDecoder.scala 133:31:@6934.4]
  wire [4:0] func; // @[InstDecoder.scala 135:21:@6936.4]
  wire  _T_903; // @[InstDecoder.scala 139:37:@6937.4]
  wire  _T_905; // @[InstDecoder.scala 137:38:@6938.4]
  wire  _T_906; // @[InstDecoder.scala 140:33:@6939.4]
  wire  _T_915; // @[InstDecoder.scala 138:39:@6946.4]
  wire  _T_916; // @[InstDecoder.scala 142:34:@6947.4]
  wire  _T_918; // @[InstDecoder.scala 136:37:@6948.4]
  wire  _T_920; // @[InstDecoder.scala 136:53:@6949.4]
  wire  _T_921; // @[InstDecoder.scala 136:45:@6950.4]
  wire [4:0] _GEN_0; // @[InstDecoder.scala 143:27:@6954.4]
  wire  _T_925; // @[InstDecoder.scala 143:27:@6954.4]
  wire  _T_927; // @[InstDecoder.scala 136:37:@6955.4]
  wire  _T_929; // @[InstDecoder.scala 136:53:@6956.4]
  wire  _T_930; // @[InstDecoder.scala 136:45:@6957.4]
  wire  _T_931; // @[InstDecoder.scala 143:44:@6958.4]
  wire  _T_938; // @[InstDecoder.scala 144:6:@6962.4]
  wire  _T_939; // @[InstDecoder.scala 144:50:@6963.4]
  wire  _T_940; // @[InstDecoder.scala 144:29:@6964.4]
  wire [11:0] imm_itype; // @[InstDecoder.scala 147:27:@6967.4]
  wire [6:0] _T_942; // @[InstDecoder.scala 148:31:@6968.4]
  wire [11:0] imm_stype; // @[Cat.scala 30:58:@6970.4]
  wire  _T_944; // @[InstDecoder.scala 149:31:@6971.4]
  wire  _T_945; // @[InstDecoder.scala 149:44:@6972.4]
  wire [5:0] _T_946; // @[InstDecoder.scala 149:56:@6973.4]
  wire [3:0] _T_947; // @[InstDecoder.scala 149:73:@6974.4]
  wire [11:0] imm_sbtype; // @[Cat.scala 30:58:@6977.4]
  wire [19:0] imm_utype; // @[InstDecoder.scala 150:27:@6978.4]
  wire [7:0] _T_951; // @[InstDecoder.scala 151:44:@6980.4]
  wire  _T_952; // @[InstDecoder.scala 151:60:@6981.4]
  wire [9:0] _T_953; // @[InstDecoder.scala 151:73:@6982.4]
  wire [19:0] imm_ujtype; // @[Cat.scala 30:58:@6985.4]
  wire  _T_956; // @[InstDecoder.scala 154:43:@6986.4]
  wire [19:0] _T_960; // @[Bitwise.scala 72:12:@6988.4]
  wire  _T_962; // @[InstDecoder.scala 155:43:@6991.4]
  wire [19:0] _T_966; // @[Bitwise.scala 72:12:@6993.4]
  wire  _T_968; // @[InstDecoder.scala 156:44:@6996.4]
  wire [18:0] _T_972; // @[Bitwise.scala 72:12:@6998.4]
  wire [30:0] _T_974; // @[Cat.scala 30:58:@6999.4]
  wire  _T_982; // @[InstDecoder.scala 158:44:@7005.4]
  wire [10:0] _T_986; // @[Bitwise.scala 72:12:@7007.4]
  wire [30:0] _T_988; // @[Cat.scala 30:58:@7008.4]
  assign _T_13 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@6115.4]
  assign _T_14 = 32'h2003 == _T_13; // @[Lookup.scala 9:38:@6116.4]
  assign _T_18 = 32'h3 == _T_13; // @[Lookup.scala 9:38:@6118.4]
  assign _T_22 = 32'h4003 == _T_13; // @[Lookup.scala 9:38:@6120.4]
  assign _T_26 = 32'h1003 == _T_13; // @[Lookup.scala 9:38:@6122.4]
  assign _T_30 = 32'h5003 == _T_13; // @[Lookup.scala 9:38:@6124.4]
  assign _T_34 = 32'h2023 == _T_13; // @[Lookup.scala 9:38:@6126.4]
  assign _T_38 = 32'h23 == _T_13; // @[Lookup.scala 9:38:@6128.4]
  assign _T_42 = 32'h1023 == _T_13; // @[Lookup.scala 9:38:@6130.4]
  assign _T_45 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@6131.4]
  assign _T_46 = 32'h17 == _T_45; // @[Lookup.scala 9:38:@6132.4]
  assign _T_50 = 32'h37 == _T_45; // @[Lookup.scala 9:38:@6134.4]
  assign _T_54 = 32'h13 == _T_13; // @[Lookup.scala 9:38:@6136.4]
  assign _T_58 = 32'h7013 == _T_13; // @[Lookup.scala 9:38:@6138.4]
  assign _T_62 = 32'h6013 == _T_13; // @[Lookup.scala 9:38:@6140.4]
  assign _T_66 = 32'h4013 == _T_13; // @[Lookup.scala 9:38:@6142.4]
  assign _T_70 = 32'h2013 == _T_13; // @[Lookup.scala 9:38:@6144.4]
  assign _T_74 = 32'h3013 == _T_13; // @[Lookup.scala 9:38:@6146.4]
  assign _T_77 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@6147.4]
  assign _T_78 = 32'h1013 == _T_77; // @[Lookup.scala 9:38:@6148.4]
  assign _T_82 = 32'h40005013 == _T_77; // @[Lookup.scala 9:38:@6150.4]
  assign _T_86 = 32'h5013 == _T_77; // @[Lookup.scala 9:38:@6152.4]
  assign _T_89 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@6153.4]
  assign _T_90 = 32'h1033 == _T_89; // @[Lookup.scala 9:38:@6154.4]
  assign _T_94 = 32'h33 == _T_89; // @[Lookup.scala 9:38:@6156.4]
  assign _T_98 = 32'h40000033 == _T_89; // @[Lookup.scala 9:38:@6158.4]
  assign _T_102 = 32'h2033 == _T_89; // @[Lookup.scala 9:38:@6160.4]
  assign _T_106 = 32'h3033 == _T_89; // @[Lookup.scala 9:38:@6162.4]
  assign _T_110 = 32'h7033 == _T_89; // @[Lookup.scala 9:38:@6164.4]
  assign _T_114 = 32'h6033 == _T_89; // @[Lookup.scala 9:38:@6166.4]
  assign _T_118 = 32'h4033 == _T_89; // @[Lookup.scala 9:38:@6168.4]
  assign _T_122 = 32'h40005033 == _T_89; // @[Lookup.scala 9:38:@6170.4]
  assign _T_126 = 32'h5033 == _T_89; // @[Lookup.scala 9:38:@6172.4]
  assign _T_130 = 32'h6f == _T_45; // @[Lookup.scala 9:38:@6174.4]
  assign _T_134 = 32'h67 == _T_13; // @[Lookup.scala 9:38:@6176.4]
  assign _T_138 = 32'h63 == _T_13; // @[Lookup.scala 9:38:@6178.4]
  assign _T_142 = 32'h1063 == _T_13; // @[Lookup.scala 9:38:@6180.4]
  assign _T_146 = 32'h5063 == _T_13; // @[Lookup.scala 9:38:@6182.4]
  assign _T_150 = 32'h7063 == _T_13; // @[Lookup.scala 9:38:@6184.4]
  assign _T_154 = 32'h4063 == _T_13; // @[Lookup.scala 9:38:@6186.4]
  assign _T_158 = 32'h6063 == _T_13; // @[Lookup.scala 9:38:@6188.4]
  assign _T_162 = 32'h5073 == _T_13; // @[Lookup.scala 9:38:@6190.4]
  assign _T_166 = 32'h6073 == _T_13; // @[Lookup.scala 9:38:@6192.4]
  assign _T_170 = 32'h1073 == _T_13; // @[Lookup.scala 9:38:@6194.4]
  assign _T_174 = 32'h2073 == _T_13; // @[Lookup.scala 9:38:@6196.4]
  assign _T_178 = 32'h3073 == _T_13; // @[Lookup.scala 9:38:@6198.4]
  assign _T_182 = 32'h7073 == _T_13; // @[Lookup.scala 9:38:@6200.4]
  assign _T_186 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@6202.4]
  assign _T_190 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@6204.4]
  assign _T_194 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@6206.4]
  assign _T_198 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@6208.4]
  assign _T_202 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@6210.4]
  assign _T_206 = 32'h100f == _T_13; // @[Lookup.scala 9:38:@6212.4]
  assign _T_210 = 32'hf == _T_13; // @[Lookup.scala 9:38:@6214.4]
  assign _T_212 = _T_206 ? 1'h1 : _T_210; // @[Lookup.scala 11:37:@6216.4]
  assign _T_213 = _T_202 ? 1'h1 : _T_212; // @[Lookup.scala 11:37:@6217.4]
  assign _T_214 = _T_198 ? 1'h1 : _T_213; // @[Lookup.scala 11:37:@6218.4]
  assign _T_215 = _T_194 ? 1'h1 : _T_214; // @[Lookup.scala 11:37:@6219.4]
  assign _T_216 = _T_190 ? 1'h1 : _T_215; // @[Lookup.scala 11:37:@6220.4]
  assign _T_217 = _T_186 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@6221.4]
  assign _T_218 = _T_182 ? 1'h1 : _T_217; // @[Lookup.scala 11:37:@6222.4]
  assign _T_219 = _T_178 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@6223.4]
  assign _T_220 = _T_174 ? 1'h1 : _T_219; // @[Lookup.scala 11:37:@6224.4]
  assign _T_221 = _T_170 ? 1'h1 : _T_220; // @[Lookup.scala 11:37:@6225.4]
  assign _T_222 = _T_166 ? 1'h1 : _T_221; // @[Lookup.scala 11:37:@6226.4]
  assign _T_223 = _T_162 ? 1'h1 : _T_222; // @[Lookup.scala 11:37:@6227.4]
  assign _T_224 = _T_158 ? 1'h1 : _T_223; // @[Lookup.scala 11:37:@6228.4]
  assign _T_225 = _T_154 ? 1'h1 : _T_224; // @[Lookup.scala 11:37:@6229.4]
  assign _T_226 = _T_150 ? 1'h1 : _T_225; // @[Lookup.scala 11:37:@6230.4]
  assign _T_227 = _T_146 ? 1'h1 : _T_226; // @[Lookup.scala 11:37:@6231.4]
  assign _T_228 = _T_142 ? 1'h1 : _T_227; // @[Lookup.scala 11:37:@6232.4]
  assign _T_229 = _T_138 ? 1'h1 : _T_228; // @[Lookup.scala 11:37:@6233.4]
  assign _T_230 = _T_134 ? 1'h1 : _T_229; // @[Lookup.scala 11:37:@6234.4]
  assign _T_231 = _T_130 ? 1'h1 : _T_230; // @[Lookup.scala 11:37:@6235.4]
  assign _T_232 = _T_126 ? 1'h1 : _T_231; // @[Lookup.scala 11:37:@6236.4]
  assign _T_233 = _T_122 ? 1'h1 : _T_232; // @[Lookup.scala 11:37:@6237.4]
  assign _T_234 = _T_118 ? 1'h1 : _T_233; // @[Lookup.scala 11:37:@6238.4]
  assign _T_235 = _T_114 ? 1'h1 : _T_234; // @[Lookup.scala 11:37:@6239.4]
  assign _T_236 = _T_110 ? 1'h1 : _T_235; // @[Lookup.scala 11:37:@6240.4]
  assign _T_237 = _T_106 ? 1'h1 : _T_236; // @[Lookup.scala 11:37:@6241.4]
  assign _T_238 = _T_102 ? 1'h1 : _T_237; // @[Lookup.scala 11:37:@6242.4]
  assign _T_239 = _T_98 ? 1'h1 : _T_238; // @[Lookup.scala 11:37:@6243.4]
  assign _T_240 = _T_94 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@6244.4]
  assign _T_241 = _T_90 ? 1'h1 : _T_240; // @[Lookup.scala 11:37:@6245.4]
  assign _T_242 = _T_86 ? 1'h1 : _T_241; // @[Lookup.scala 11:37:@6246.4]
  assign _T_243 = _T_82 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@6247.4]
  assign _T_244 = _T_78 ? 1'h1 : _T_243; // @[Lookup.scala 11:37:@6248.4]
  assign _T_245 = _T_74 ? 1'h1 : _T_244; // @[Lookup.scala 11:37:@6249.4]
  assign _T_246 = _T_70 ? 1'h1 : _T_245; // @[Lookup.scala 11:37:@6250.4]
  assign _T_247 = _T_66 ? 1'h1 : _T_246; // @[Lookup.scala 11:37:@6251.4]
  assign _T_248 = _T_62 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@6252.4]
  assign _T_249 = _T_58 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@6253.4]
  assign _T_250 = _T_54 ? 1'h1 : _T_249; // @[Lookup.scala 11:37:@6254.4]
  assign _T_251 = _T_50 ? 1'h1 : _T_250; // @[Lookup.scala 11:37:@6255.4]
  assign _T_252 = _T_46 ? 1'h1 : _T_251; // @[Lookup.scala 11:37:@6256.4]
  assign _T_253 = _T_42 ? 1'h1 : _T_252; // @[Lookup.scala 11:37:@6257.4]
  assign _T_254 = _T_38 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@6258.4]
  assign _T_255 = _T_34 ? 1'h1 : _T_254; // @[Lookup.scala 11:37:@6259.4]
  assign _T_256 = _T_30 ? 1'h1 : _T_255; // @[Lookup.scala 11:37:@6260.4]
  assign _T_257 = _T_26 ? 1'h1 : _T_256; // @[Lookup.scala 11:37:@6261.4]
  assign _T_258 = _T_22 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:@6262.4]
  assign _T_259 = _T_18 ? 1'h1 : _T_258; // @[Lookup.scala 11:37:@6263.4]
  assign signals_0 = _T_14 ? 1'h1 : _T_259; // @[Lookup.scala 11:37:@6264.4]
  assign _T_273 = _T_158 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@6278.4]
  assign _T_274 = _T_154 ? 4'h5 : _T_273; // @[Lookup.scala 11:37:@6279.4]
  assign _T_275 = _T_150 ? 4'h4 : _T_274; // @[Lookup.scala 11:37:@6280.4]
  assign _T_276 = _T_146 ? 4'h3 : _T_275; // @[Lookup.scala 11:37:@6281.4]
  assign _T_277 = _T_142 ? 4'h1 : _T_276; // @[Lookup.scala 11:37:@6282.4]
  assign _T_278 = _T_138 ? 4'h2 : _T_277; // @[Lookup.scala 11:37:@6283.4]
  assign _T_279 = _T_134 ? 4'h8 : _T_278; // @[Lookup.scala 11:37:@6284.4]
  assign _T_280 = _T_130 ? 4'h7 : _T_279; // @[Lookup.scala 11:37:@6285.4]
  assign _T_281 = _T_126 ? 4'h0 : _T_280; // @[Lookup.scala 11:37:@6286.4]
  assign _T_282 = _T_122 ? 4'h0 : _T_281; // @[Lookup.scala 11:37:@6287.4]
  assign _T_283 = _T_118 ? 4'h0 : _T_282; // @[Lookup.scala 11:37:@6288.4]
  assign _T_284 = _T_114 ? 4'h0 : _T_283; // @[Lookup.scala 11:37:@6289.4]
  assign _T_285 = _T_110 ? 4'h0 : _T_284; // @[Lookup.scala 11:37:@6290.4]
  assign _T_286 = _T_106 ? 4'h0 : _T_285; // @[Lookup.scala 11:37:@6291.4]
  assign _T_287 = _T_102 ? 4'h0 : _T_286; // @[Lookup.scala 11:37:@6292.4]
  assign _T_288 = _T_98 ? 4'h0 : _T_287; // @[Lookup.scala 11:37:@6293.4]
  assign _T_289 = _T_94 ? 4'h0 : _T_288; // @[Lookup.scala 11:37:@6294.4]
  assign _T_290 = _T_90 ? 4'h0 : _T_289; // @[Lookup.scala 11:37:@6295.4]
  assign _T_291 = _T_86 ? 4'h0 : _T_290; // @[Lookup.scala 11:37:@6296.4]
  assign _T_292 = _T_82 ? 4'h0 : _T_291; // @[Lookup.scala 11:37:@6297.4]
  assign _T_293 = _T_78 ? 4'h0 : _T_292; // @[Lookup.scala 11:37:@6298.4]
  assign _T_294 = _T_74 ? 4'h0 : _T_293; // @[Lookup.scala 11:37:@6299.4]
  assign _T_295 = _T_70 ? 4'h0 : _T_294; // @[Lookup.scala 11:37:@6300.4]
  assign _T_296 = _T_66 ? 4'h0 : _T_295; // @[Lookup.scala 11:37:@6301.4]
  assign _T_297 = _T_62 ? 4'h0 : _T_296; // @[Lookup.scala 11:37:@6302.4]
  assign _T_298 = _T_58 ? 4'h0 : _T_297; // @[Lookup.scala 11:37:@6303.4]
  assign _T_299 = _T_54 ? 4'h0 : _T_298; // @[Lookup.scala 11:37:@6304.4]
  assign _T_300 = _T_50 ? 4'h0 : _T_299; // @[Lookup.scala 11:37:@6305.4]
  assign _T_301 = _T_46 ? 4'h0 : _T_300; // @[Lookup.scala 11:37:@6306.4]
  assign _T_302 = _T_42 ? 4'h0 : _T_301; // @[Lookup.scala 11:37:@6307.4]
  assign _T_303 = _T_38 ? 4'h0 : _T_302; // @[Lookup.scala 11:37:@6308.4]
  assign _T_304 = _T_34 ? 4'h0 : _T_303; // @[Lookup.scala 11:37:@6309.4]
  assign _T_305 = _T_30 ? 4'h0 : _T_304; // @[Lookup.scala 11:37:@6310.4]
  assign _T_306 = _T_26 ? 4'h0 : _T_305; // @[Lookup.scala 11:37:@6311.4]
  assign _T_307 = _T_22 ? 4'h0 : _T_306; // @[Lookup.scala 11:37:@6312.4]
  assign _T_308 = _T_18 ? 4'h0 : _T_307; // @[Lookup.scala 11:37:@6313.4]
  assign _T_316 = _T_182 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@6322.4]
  assign _T_317 = _T_178 ? 2'h0 : _T_316; // @[Lookup.scala 11:37:@6323.4]
  assign _T_318 = _T_174 ? 2'h0 : _T_317; // @[Lookup.scala 11:37:@6324.4]
  assign _T_319 = _T_170 ? 2'h0 : _T_318; // @[Lookup.scala 11:37:@6325.4]
  assign _T_320 = _T_166 ? 2'h2 : _T_319; // @[Lookup.scala 11:37:@6326.4]
  assign _T_321 = _T_162 ? 2'h2 : _T_320; // @[Lookup.scala 11:37:@6327.4]
  assign _T_322 = _T_158 ? 2'h0 : _T_321; // @[Lookup.scala 11:37:@6328.4]
  assign _T_323 = _T_154 ? 2'h0 : _T_322; // @[Lookup.scala 11:37:@6329.4]
  assign _T_324 = _T_150 ? 2'h0 : _T_323; // @[Lookup.scala 11:37:@6330.4]
  assign _T_325 = _T_146 ? 2'h0 : _T_324; // @[Lookup.scala 11:37:@6331.4]
  assign _T_326 = _T_142 ? 2'h0 : _T_325; // @[Lookup.scala 11:37:@6332.4]
  assign _T_327 = _T_138 ? 2'h0 : _T_326; // @[Lookup.scala 11:37:@6333.4]
  assign _T_328 = _T_134 ? 2'h0 : _T_327; // @[Lookup.scala 11:37:@6334.4]
  assign _T_329 = _T_130 ? 2'h0 : _T_328; // @[Lookup.scala 11:37:@6335.4]
  assign _T_330 = _T_126 ? 2'h0 : _T_329; // @[Lookup.scala 11:37:@6336.4]
  assign _T_331 = _T_122 ? 2'h0 : _T_330; // @[Lookup.scala 11:37:@6337.4]
  assign _T_332 = _T_118 ? 2'h0 : _T_331; // @[Lookup.scala 11:37:@6338.4]
  assign _T_333 = _T_114 ? 2'h0 : _T_332; // @[Lookup.scala 11:37:@6339.4]
  assign _T_334 = _T_110 ? 2'h0 : _T_333; // @[Lookup.scala 11:37:@6340.4]
  assign _T_335 = _T_106 ? 2'h0 : _T_334; // @[Lookup.scala 11:37:@6341.4]
  assign _T_336 = _T_102 ? 2'h0 : _T_335; // @[Lookup.scala 11:37:@6342.4]
  assign _T_337 = _T_98 ? 2'h0 : _T_336; // @[Lookup.scala 11:37:@6343.4]
  assign _T_338 = _T_94 ? 2'h0 : _T_337; // @[Lookup.scala 11:37:@6344.4]
  assign _T_339 = _T_90 ? 2'h0 : _T_338; // @[Lookup.scala 11:37:@6345.4]
  assign _T_340 = _T_86 ? 2'h0 : _T_339; // @[Lookup.scala 11:37:@6346.4]
  assign _T_341 = _T_82 ? 2'h0 : _T_340; // @[Lookup.scala 11:37:@6347.4]
  assign _T_342 = _T_78 ? 2'h0 : _T_341; // @[Lookup.scala 11:37:@6348.4]
  assign _T_343 = _T_74 ? 2'h0 : _T_342; // @[Lookup.scala 11:37:@6349.4]
  assign _T_344 = _T_70 ? 2'h0 : _T_343; // @[Lookup.scala 11:37:@6350.4]
  assign _T_345 = _T_66 ? 2'h0 : _T_344; // @[Lookup.scala 11:37:@6351.4]
  assign _T_346 = _T_62 ? 2'h0 : _T_345; // @[Lookup.scala 11:37:@6352.4]
  assign _T_347 = _T_58 ? 2'h0 : _T_346; // @[Lookup.scala 11:37:@6353.4]
  assign _T_348 = _T_54 ? 2'h0 : _T_347; // @[Lookup.scala 11:37:@6354.4]
  assign _T_349 = _T_50 ? 2'h0 : _T_348; // @[Lookup.scala 11:37:@6355.4]
  assign _T_350 = _T_46 ? 2'h1 : _T_349; // @[Lookup.scala 11:37:@6356.4]
  assign _T_351 = _T_42 ? 2'h0 : _T_350; // @[Lookup.scala 11:37:@6357.4]
  assign _T_352 = _T_38 ? 2'h0 : _T_351; // @[Lookup.scala 11:37:@6358.4]
  assign _T_353 = _T_34 ? 2'h0 : _T_352; // @[Lookup.scala 11:37:@6359.4]
  assign _T_354 = _T_30 ? 2'h0 : _T_353; // @[Lookup.scala 11:37:@6360.4]
  assign _T_355 = _T_26 ? 2'h0 : _T_354; // @[Lookup.scala 11:37:@6361.4]
  assign _T_356 = _T_22 ? 2'h0 : _T_355; // @[Lookup.scala 11:37:@6362.4]
  assign _T_357 = _T_18 ? 2'h0 : _T_356; // @[Lookup.scala 11:37:@6363.4]
  assign _T_371 = _T_158 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37:@6378.4]
  assign _T_372 = _T_154 ? 3'h3 : _T_371; // @[Lookup.scala 11:37:@6379.4]
  assign _T_373 = _T_150 ? 3'h3 : _T_372; // @[Lookup.scala 11:37:@6380.4]
  assign _T_374 = _T_146 ? 3'h3 : _T_373; // @[Lookup.scala 11:37:@6381.4]
  assign _T_375 = _T_142 ? 3'h3 : _T_374; // @[Lookup.scala 11:37:@6382.4]
  assign _T_376 = _T_138 ? 3'h3 : _T_375; // @[Lookup.scala 11:37:@6383.4]
  assign _T_377 = _T_134 ? 3'h1 : _T_376; // @[Lookup.scala 11:37:@6384.4]
  assign _T_378 = _T_130 ? 3'h5 : _T_377; // @[Lookup.scala 11:37:@6385.4]
  assign _T_379 = _T_126 ? 3'h0 : _T_378; // @[Lookup.scala 11:37:@6386.4]
  assign _T_380 = _T_122 ? 3'h0 : _T_379; // @[Lookup.scala 11:37:@6387.4]
  assign _T_381 = _T_118 ? 3'h0 : _T_380; // @[Lookup.scala 11:37:@6388.4]
  assign _T_382 = _T_114 ? 3'h0 : _T_381; // @[Lookup.scala 11:37:@6389.4]
  assign _T_383 = _T_110 ? 3'h0 : _T_382; // @[Lookup.scala 11:37:@6390.4]
  assign _T_384 = _T_106 ? 3'h0 : _T_383; // @[Lookup.scala 11:37:@6391.4]
  assign _T_385 = _T_102 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@6392.4]
  assign _T_386 = _T_98 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@6393.4]
  assign _T_387 = _T_94 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@6394.4]
  assign _T_388 = _T_90 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@6395.4]
  assign _T_389 = _T_86 ? 3'h1 : _T_388; // @[Lookup.scala 11:37:@6396.4]
  assign _T_390 = _T_82 ? 3'h1 : _T_389; // @[Lookup.scala 11:37:@6397.4]
  assign _T_391 = _T_78 ? 3'h1 : _T_390; // @[Lookup.scala 11:37:@6398.4]
  assign _T_392 = _T_74 ? 3'h1 : _T_391; // @[Lookup.scala 11:37:@6399.4]
  assign _T_393 = _T_70 ? 3'h1 : _T_392; // @[Lookup.scala 11:37:@6400.4]
  assign _T_394 = _T_66 ? 3'h1 : _T_393; // @[Lookup.scala 11:37:@6401.4]
  assign _T_395 = _T_62 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@6402.4]
  assign _T_396 = _T_58 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@6403.4]
  assign _T_397 = _T_54 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@6404.4]
  assign _T_398 = _T_50 ? 3'h4 : _T_397; // @[Lookup.scala 11:37:@6405.4]
  assign _T_399 = _T_46 ? 3'h4 : _T_398; // @[Lookup.scala 11:37:@6406.4]
  assign _T_400 = _T_42 ? 3'h2 : _T_399; // @[Lookup.scala 11:37:@6407.4]
  assign _T_401 = _T_38 ? 3'h2 : _T_400; // @[Lookup.scala 11:37:@6408.4]
  assign _T_402 = _T_34 ? 3'h2 : _T_401; // @[Lookup.scala 11:37:@6409.4]
  assign _T_403 = _T_30 ? 3'h1 : _T_402; // @[Lookup.scala 11:37:@6410.4]
  assign _T_404 = _T_26 ? 3'h1 : _T_403; // @[Lookup.scala 11:37:@6411.4]
  assign _T_405 = _T_22 ? 3'h1 : _T_404; // @[Lookup.scala 11:37:@6412.4]
  assign _T_406 = _T_18 ? 3'h1 : _T_405; // @[Lookup.scala 11:37:@6413.4]
  assign _T_415 = _T_178 ? 1'h1 : _T_182; // @[Lookup.scala 11:37:@6423.4]
  assign _T_416 = _T_174 ? 1'h1 : _T_415; // @[Lookup.scala 11:37:@6424.4]
  assign _T_417 = _T_170 ? 1'h1 : _T_416; // @[Lookup.scala 11:37:@6425.4]
  assign _T_418 = _T_166 ? 1'h1 : _T_417; // @[Lookup.scala 11:37:@6426.4]
  assign _T_419 = _T_162 ? 1'h1 : _T_418; // @[Lookup.scala 11:37:@6427.4]
  assign _T_420 = _T_158 ? 1'h1 : _T_419; // @[Lookup.scala 11:37:@6428.4]
  assign _T_421 = _T_154 ? 1'h1 : _T_420; // @[Lookup.scala 11:37:@6429.4]
  assign _T_422 = _T_150 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@6430.4]
  assign _T_423 = _T_146 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@6431.4]
  assign _T_424 = _T_142 ? 1'h1 : _T_423; // @[Lookup.scala 11:37:@6432.4]
  assign _T_425 = _T_138 ? 1'h1 : _T_424; // @[Lookup.scala 11:37:@6433.4]
  assign _T_426 = _T_134 ? 1'h1 : _T_425; // @[Lookup.scala 11:37:@6434.4]
  assign _T_427 = _T_130 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:@6435.4]
  assign _T_428 = _T_126 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@6436.4]
  assign _T_429 = _T_122 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@6437.4]
  assign _T_430 = _T_118 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@6438.4]
  assign _T_431 = _T_114 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@6439.4]
  assign _T_432 = _T_110 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@6440.4]
  assign _T_433 = _T_106 ? 1'h1 : _T_432; // @[Lookup.scala 11:37:@6441.4]
  assign _T_434 = _T_102 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@6442.4]
  assign _T_435 = _T_98 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@6443.4]
  assign _T_436 = _T_94 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@6444.4]
  assign _T_437 = _T_90 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@6445.4]
  assign _T_438 = _T_86 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@6446.4]
  assign _T_439 = _T_82 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@6447.4]
  assign _T_440 = _T_78 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@6448.4]
  assign _T_441 = _T_74 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@6449.4]
  assign _T_442 = _T_70 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@6450.4]
  assign _T_443 = _T_66 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@6451.4]
  assign _T_444 = _T_62 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@6452.4]
  assign _T_445 = _T_58 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@6453.4]
  assign _T_446 = _T_54 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@6454.4]
  assign _T_447 = _T_50 ? 1'h0 : _T_446; // @[Lookup.scala 11:37:@6455.4]
  assign _T_448 = _T_46 ? 1'h0 : _T_447; // @[Lookup.scala 11:37:@6456.4]
  assign _T_449 = _T_42 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@6457.4]
  assign _T_450 = _T_38 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@6458.4]
  assign _T_451 = _T_34 ? 1'h1 : _T_450; // @[Lookup.scala 11:37:@6459.4]
  assign _T_452 = _T_30 ? 1'h1 : _T_451; // @[Lookup.scala 11:37:@6460.4]
  assign _T_453 = _T_26 ? 1'h1 : _T_452; // @[Lookup.scala 11:37:@6461.4]
  assign _T_454 = _T_22 ? 1'h1 : _T_453; // @[Lookup.scala 11:37:@6462.4]
  assign _T_455 = _T_18 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@6463.4]
  assign _T_475 = _T_134 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@6484.4]
  assign _T_476 = _T_130 ? 1'h0 : _T_475; // @[Lookup.scala 11:37:@6485.4]
  assign _T_477 = _T_126 ? 1'h1 : _T_476; // @[Lookup.scala 11:37:@6486.4]
  assign _T_478 = _T_122 ? 1'h1 : _T_477; // @[Lookup.scala 11:37:@6487.4]
  assign _T_479 = _T_118 ? 1'h1 : _T_478; // @[Lookup.scala 11:37:@6488.4]
  assign _T_480 = _T_114 ? 1'h1 : _T_479; // @[Lookup.scala 11:37:@6489.4]
  assign _T_481 = _T_110 ? 1'h1 : _T_480; // @[Lookup.scala 11:37:@6490.4]
  assign _T_482 = _T_106 ? 1'h1 : _T_481; // @[Lookup.scala 11:37:@6491.4]
  assign _T_483 = _T_102 ? 1'h1 : _T_482; // @[Lookup.scala 11:37:@6492.4]
  assign _T_484 = _T_98 ? 1'h1 : _T_483; // @[Lookup.scala 11:37:@6493.4]
  assign _T_485 = _T_94 ? 1'h1 : _T_484; // @[Lookup.scala 11:37:@6494.4]
  assign _T_486 = _T_90 ? 1'h1 : _T_485; // @[Lookup.scala 11:37:@6495.4]
  assign _T_487 = _T_86 ? 1'h0 : _T_486; // @[Lookup.scala 11:37:@6496.4]
  assign _T_488 = _T_82 ? 1'h0 : _T_487; // @[Lookup.scala 11:37:@6497.4]
  assign _T_489 = _T_78 ? 1'h0 : _T_488; // @[Lookup.scala 11:37:@6498.4]
  assign _T_490 = _T_74 ? 1'h0 : _T_489; // @[Lookup.scala 11:37:@6499.4]
  assign _T_491 = _T_70 ? 1'h0 : _T_490; // @[Lookup.scala 11:37:@6500.4]
  assign _T_492 = _T_66 ? 1'h0 : _T_491; // @[Lookup.scala 11:37:@6501.4]
  assign _T_493 = _T_62 ? 1'h0 : _T_492; // @[Lookup.scala 11:37:@6502.4]
  assign _T_494 = _T_58 ? 1'h0 : _T_493; // @[Lookup.scala 11:37:@6503.4]
  assign _T_495 = _T_54 ? 1'h0 : _T_494; // @[Lookup.scala 11:37:@6504.4]
  assign _T_496 = _T_50 ? 1'h0 : _T_495; // @[Lookup.scala 11:37:@6505.4]
  assign _T_497 = _T_46 ? 1'h0 : _T_496; // @[Lookup.scala 11:37:@6506.4]
  assign _T_498 = _T_42 ? 1'h1 : _T_497; // @[Lookup.scala 11:37:@6507.4]
  assign _T_499 = _T_38 ? 1'h1 : _T_498; // @[Lookup.scala 11:37:@6508.4]
  assign _T_500 = _T_34 ? 1'h1 : _T_499; // @[Lookup.scala 11:37:@6509.4]
  assign _T_501 = _T_30 ? 1'h0 : _T_500; // @[Lookup.scala 11:37:@6510.4]
  assign _T_502 = _T_26 ? 1'h0 : _T_501; // @[Lookup.scala 11:37:@6511.4]
  assign _T_503 = _T_22 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@6512.4]
  assign _T_504 = _T_18 ? 1'h0 : _T_503; // @[Lookup.scala 11:37:@6513.4]
  assign _T_512 = _T_182 ? 4'ha : 4'h0; // @[Lookup.scala 11:37:@6522.4]
  assign _T_513 = _T_178 ? 4'ha : _T_512; // @[Lookup.scala 11:37:@6523.4]
  assign _T_514 = _T_174 ? 4'ha : _T_513; // @[Lookup.scala 11:37:@6524.4]
  assign _T_515 = _T_170 ? 4'ha : _T_514; // @[Lookup.scala 11:37:@6525.4]
  assign _T_516 = _T_166 ? 4'ha : _T_515; // @[Lookup.scala 11:37:@6526.4]
  assign _T_517 = _T_162 ? 4'ha : _T_516; // @[Lookup.scala 11:37:@6527.4]
  assign _T_518 = _T_158 ? 4'h0 : _T_517; // @[Lookup.scala 11:37:@6528.4]
  assign _T_519 = _T_154 ? 4'h0 : _T_518; // @[Lookup.scala 11:37:@6529.4]
  assign _T_520 = _T_150 ? 4'h0 : _T_519; // @[Lookup.scala 11:37:@6530.4]
  assign _T_521 = _T_146 ? 4'h0 : _T_520; // @[Lookup.scala 11:37:@6531.4]
  assign _T_522 = _T_142 ? 4'h0 : _T_521; // @[Lookup.scala 11:37:@6532.4]
  assign _T_523 = _T_138 ? 4'h0 : _T_522; // @[Lookup.scala 11:37:@6533.4]
  assign _T_524 = _T_134 ? 4'h0 : _T_523; // @[Lookup.scala 11:37:@6534.4]
  assign _T_525 = _T_130 ? 4'h0 : _T_524; // @[Lookup.scala 11:37:@6535.4]
  assign _T_526 = _T_126 ? 4'h3 : _T_525; // @[Lookup.scala 11:37:@6536.4]
  assign _T_527 = _T_122 ? 4'h4 : _T_526; // @[Lookup.scala 11:37:@6537.4]
  assign _T_528 = _T_118 ? 4'h7 : _T_527; // @[Lookup.scala 11:37:@6538.4]
  assign _T_529 = _T_114 ? 4'h6 : _T_528; // @[Lookup.scala 11:37:@6539.4]
  assign _T_530 = _T_110 ? 4'h5 : _T_529; // @[Lookup.scala 11:37:@6540.4]
  assign _T_531 = _T_106 ? 4'h9 : _T_530; // @[Lookup.scala 11:37:@6541.4]
  assign _T_532 = _T_102 ? 4'h8 : _T_531; // @[Lookup.scala 11:37:@6542.4]
  assign _T_533 = _T_98 ? 4'h1 : _T_532; // @[Lookup.scala 11:37:@6543.4]
  assign _T_534 = _T_94 ? 4'h0 : _T_533; // @[Lookup.scala 11:37:@6544.4]
  assign _T_535 = _T_90 ? 4'h2 : _T_534; // @[Lookup.scala 11:37:@6545.4]
  assign _T_536 = _T_86 ? 4'h3 : _T_535; // @[Lookup.scala 11:37:@6546.4]
  assign _T_537 = _T_82 ? 4'h4 : _T_536; // @[Lookup.scala 11:37:@6547.4]
  assign _T_538 = _T_78 ? 4'h2 : _T_537; // @[Lookup.scala 11:37:@6548.4]
  assign _T_539 = _T_74 ? 4'h9 : _T_538; // @[Lookup.scala 11:37:@6549.4]
  assign _T_540 = _T_70 ? 4'h8 : _T_539; // @[Lookup.scala 11:37:@6550.4]
  assign _T_541 = _T_66 ? 4'h7 : _T_540; // @[Lookup.scala 11:37:@6551.4]
  assign _T_542 = _T_62 ? 4'h6 : _T_541; // @[Lookup.scala 11:37:@6552.4]
  assign _T_543 = _T_58 ? 4'h5 : _T_542; // @[Lookup.scala 11:37:@6553.4]
  assign _T_544 = _T_54 ? 4'h0 : _T_543; // @[Lookup.scala 11:37:@6554.4]
  assign _T_545 = _T_50 ? 4'hb : _T_544; // @[Lookup.scala 11:37:@6555.4]
  assign _T_546 = _T_46 ? 4'h0 : _T_545; // @[Lookup.scala 11:37:@6556.4]
  assign _T_547 = _T_42 ? 4'h0 : _T_546; // @[Lookup.scala 11:37:@6557.4]
  assign _T_548 = _T_38 ? 4'h0 : _T_547; // @[Lookup.scala 11:37:@6558.4]
  assign _T_549 = _T_34 ? 4'h0 : _T_548; // @[Lookup.scala 11:37:@6559.4]
  assign _T_550 = _T_30 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:@6560.4]
  assign _T_551 = _T_26 ? 4'h0 : _T_550; // @[Lookup.scala 11:37:@6561.4]
  assign _T_552 = _T_22 ? 4'h0 : _T_551; // @[Lookup.scala 11:37:@6562.4]
  assign _T_553 = _T_18 ? 4'h0 : _T_552; // @[Lookup.scala 11:37:@6563.4]
  assign _T_561 = _T_182 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@6572.4]
  assign _T_562 = _T_178 ? 2'h3 : _T_561; // @[Lookup.scala 11:37:@6573.4]
  assign _T_563 = _T_174 ? 2'h3 : _T_562; // @[Lookup.scala 11:37:@6574.4]
  assign _T_564 = _T_170 ? 2'h3 : _T_563; // @[Lookup.scala 11:37:@6575.4]
  assign _T_565 = _T_166 ? 2'h3 : _T_564; // @[Lookup.scala 11:37:@6576.4]
  assign _T_566 = _T_162 ? 2'h3 : _T_565; // @[Lookup.scala 11:37:@6577.4]
  assign _T_567 = _T_158 ? 2'h0 : _T_566; // @[Lookup.scala 11:37:@6578.4]
  assign _T_568 = _T_154 ? 2'h0 : _T_567; // @[Lookup.scala 11:37:@6579.4]
  assign _T_569 = _T_150 ? 2'h0 : _T_568; // @[Lookup.scala 11:37:@6580.4]
  assign _T_570 = _T_146 ? 2'h0 : _T_569; // @[Lookup.scala 11:37:@6581.4]
  assign _T_571 = _T_142 ? 2'h0 : _T_570; // @[Lookup.scala 11:37:@6582.4]
  assign _T_572 = _T_138 ? 2'h0 : _T_571; // @[Lookup.scala 11:37:@6583.4]
  assign _T_573 = _T_134 ? 2'h2 : _T_572; // @[Lookup.scala 11:37:@6584.4]
  assign _T_574 = _T_130 ? 2'h2 : _T_573; // @[Lookup.scala 11:37:@6585.4]
  assign _T_575 = _T_126 ? 2'h0 : _T_574; // @[Lookup.scala 11:37:@6586.4]
  assign _T_576 = _T_122 ? 2'h0 : _T_575; // @[Lookup.scala 11:37:@6587.4]
  assign _T_577 = _T_118 ? 2'h0 : _T_576; // @[Lookup.scala 11:37:@6588.4]
  assign _T_578 = _T_114 ? 2'h0 : _T_577; // @[Lookup.scala 11:37:@6589.4]
  assign _T_579 = _T_110 ? 2'h0 : _T_578; // @[Lookup.scala 11:37:@6590.4]
  assign _T_580 = _T_106 ? 2'h0 : _T_579; // @[Lookup.scala 11:37:@6591.4]
  assign _T_581 = _T_102 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@6592.4]
  assign _T_582 = _T_98 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@6593.4]
  assign _T_583 = _T_94 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@6594.4]
  assign _T_584 = _T_90 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@6595.4]
  assign _T_585 = _T_86 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@6596.4]
  assign _T_586 = _T_82 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@6597.4]
  assign _T_587 = _T_78 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@6598.4]
  assign _T_588 = _T_74 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@6599.4]
  assign _T_589 = _T_70 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@6600.4]
  assign _T_590 = _T_66 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@6601.4]
  assign _T_591 = _T_62 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@6602.4]
  assign _T_592 = _T_58 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@6603.4]
  assign _T_593 = _T_54 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@6604.4]
  assign _T_594 = _T_50 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@6605.4]
  assign _T_595 = _T_46 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@6606.4]
  assign _T_596 = _T_42 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@6607.4]
  assign _T_597 = _T_38 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@6608.4]
  assign _T_598 = _T_34 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@6609.4]
  assign _T_599 = _T_30 ? 2'h1 : _T_598; // @[Lookup.scala 11:37:@6610.4]
  assign _T_600 = _T_26 ? 2'h1 : _T_599; // @[Lookup.scala 11:37:@6611.4]
  assign _T_601 = _T_22 ? 2'h1 : _T_600; // @[Lookup.scala 11:37:@6612.4]
  assign _T_602 = _T_18 ? 2'h1 : _T_601; // @[Lookup.scala 11:37:@6613.4]
  assign _T_616 = _T_158 ? 1'h0 : _T_419; // @[Lookup.scala 11:37:@6628.4]
  assign _T_617 = _T_154 ? 1'h0 : _T_616; // @[Lookup.scala 11:37:@6629.4]
  assign _T_618 = _T_150 ? 1'h0 : _T_617; // @[Lookup.scala 11:37:@6630.4]
  assign _T_619 = _T_146 ? 1'h0 : _T_618; // @[Lookup.scala 11:37:@6631.4]
  assign _T_620 = _T_142 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@6632.4]
  assign _T_621 = _T_138 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@6633.4]
  assign _T_622 = _T_134 ? 1'h1 : _T_621; // @[Lookup.scala 11:37:@6634.4]
  assign _T_623 = _T_130 ? 1'h1 : _T_622; // @[Lookup.scala 11:37:@6635.4]
  assign _T_624 = _T_126 ? 1'h1 : _T_623; // @[Lookup.scala 11:37:@6636.4]
  assign _T_625 = _T_122 ? 1'h1 : _T_624; // @[Lookup.scala 11:37:@6637.4]
  assign _T_626 = _T_118 ? 1'h1 : _T_625; // @[Lookup.scala 11:37:@6638.4]
  assign _T_627 = _T_114 ? 1'h1 : _T_626; // @[Lookup.scala 11:37:@6639.4]
  assign _T_628 = _T_110 ? 1'h1 : _T_627; // @[Lookup.scala 11:37:@6640.4]
  assign _T_629 = _T_106 ? 1'h1 : _T_628; // @[Lookup.scala 11:37:@6641.4]
  assign _T_630 = _T_102 ? 1'h1 : _T_629; // @[Lookup.scala 11:37:@6642.4]
  assign _T_631 = _T_98 ? 1'h1 : _T_630; // @[Lookup.scala 11:37:@6643.4]
  assign _T_632 = _T_94 ? 1'h1 : _T_631; // @[Lookup.scala 11:37:@6644.4]
  assign _T_633 = _T_90 ? 1'h1 : _T_632; // @[Lookup.scala 11:37:@6645.4]
  assign _T_634 = _T_86 ? 1'h1 : _T_633; // @[Lookup.scala 11:37:@6646.4]
  assign _T_635 = _T_82 ? 1'h1 : _T_634; // @[Lookup.scala 11:37:@6647.4]
  assign _T_636 = _T_78 ? 1'h1 : _T_635; // @[Lookup.scala 11:37:@6648.4]
  assign _T_637 = _T_74 ? 1'h1 : _T_636; // @[Lookup.scala 11:37:@6649.4]
  assign _T_638 = _T_70 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:@6650.4]
  assign _T_639 = _T_66 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:@6651.4]
  assign _T_640 = _T_62 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:@6652.4]
  assign _T_641 = _T_58 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:@6653.4]
  assign _T_642 = _T_54 ? 1'h1 : _T_641; // @[Lookup.scala 11:37:@6654.4]
  assign _T_643 = _T_50 ? 1'h1 : _T_642; // @[Lookup.scala 11:37:@6655.4]
  assign _T_644 = _T_46 ? 1'h1 : _T_643; // @[Lookup.scala 11:37:@6656.4]
  assign _T_645 = _T_42 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:@6657.4]
  assign _T_646 = _T_38 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:@6658.4]
  assign _T_647 = _T_34 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:@6659.4]
  assign _T_648 = _T_30 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:@6660.4]
  assign _T_649 = _T_26 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:@6661.4]
  assign _T_650 = _T_22 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:@6662.4]
  assign _T_651 = _T_18 ? 1'h1 : _T_650; // @[Lookup.scala 11:37:@6663.4]
  assign _T_653 = _T_206 ? 1'h0 : _T_210; // @[Lookup.scala 11:37:@6666.4]
  assign _T_654 = _T_202 ? 1'h0 : _T_653; // @[Lookup.scala 11:37:@6667.4]
  assign _T_655 = _T_198 ? 1'h0 : _T_654; // @[Lookup.scala 11:37:@6668.4]
  assign _T_656 = _T_194 ? 1'h0 : _T_655; // @[Lookup.scala 11:37:@6669.4]
  assign _T_657 = _T_190 ? 1'h0 : _T_656; // @[Lookup.scala 11:37:@6670.4]
  assign _T_658 = _T_186 ? 1'h0 : _T_657; // @[Lookup.scala 11:37:@6671.4]
  assign _T_659 = _T_182 ? 1'h0 : _T_658; // @[Lookup.scala 11:37:@6672.4]
  assign _T_660 = _T_178 ? 1'h0 : _T_659; // @[Lookup.scala 11:37:@6673.4]
  assign _T_661 = _T_174 ? 1'h0 : _T_660; // @[Lookup.scala 11:37:@6674.4]
  assign _T_662 = _T_170 ? 1'h0 : _T_661; // @[Lookup.scala 11:37:@6675.4]
  assign _T_663 = _T_166 ? 1'h0 : _T_662; // @[Lookup.scala 11:37:@6676.4]
  assign _T_664 = _T_162 ? 1'h0 : _T_663; // @[Lookup.scala 11:37:@6677.4]
  assign _T_665 = _T_158 ? 1'h0 : _T_664; // @[Lookup.scala 11:37:@6678.4]
  assign _T_666 = _T_154 ? 1'h0 : _T_665; // @[Lookup.scala 11:37:@6679.4]
  assign _T_667 = _T_150 ? 1'h0 : _T_666; // @[Lookup.scala 11:37:@6680.4]
  assign _T_668 = _T_146 ? 1'h0 : _T_667; // @[Lookup.scala 11:37:@6681.4]
  assign _T_669 = _T_142 ? 1'h0 : _T_668; // @[Lookup.scala 11:37:@6682.4]
  assign _T_670 = _T_138 ? 1'h0 : _T_669; // @[Lookup.scala 11:37:@6683.4]
  assign _T_671 = _T_134 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:@6684.4]
  assign _T_672 = _T_130 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:@6685.4]
  assign _T_673 = _T_126 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:@6686.4]
  assign _T_674 = _T_122 ? 1'h0 : _T_673; // @[Lookup.scala 11:37:@6687.4]
  assign _T_675 = _T_118 ? 1'h0 : _T_674; // @[Lookup.scala 11:37:@6688.4]
  assign _T_676 = _T_114 ? 1'h0 : _T_675; // @[Lookup.scala 11:37:@6689.4]
  assign _T_677 = _T_110 ? 1'h0 : _T_676; // @[Lookup.scala 11:37:@6690.4]
  assign _T_678 = _T_106 ? 1'h0 : _T_677; // @[Lookup.scala 11:37:@6691.4]
  assign _T_679 = _T_102 ? 1'h0 : _T_678; // @[Lookup.scala 11:37:@6692.4]
  assign _T_680 = _T_98 ? 1'h0 : _T_679; // @[Lookup.scala 11:37:@6693.4]
  assign _T_681 = _T_94 ? 1'h0 : _T_680; // @[Lookup.scala 11:37:@6694.4]
  assign _T_682 = _T_90 ? 1'h0 : _T_681; // @[Lookup.scala 11:37:@6695.4]
  assign _T_683 = _T_86 ? 1'h0 : _T_682; // @[Lookup.scala 11:37:@6696.4]
  assign _T_684 = _T_82 ? 1'h0 : _T_683; // @[Lookup.scala 11:37:@6697.4]
  assign _T_685 = _T_78 ? 1'h0 : _T_684; // @[Lookup.scala 11:37:@6698.4]
  assign _T_686 = _T_74 ? 1'h0 : _T_685; // @[Lookup.scala 11:37:@6699.4]
  assign _T_687 = _T_70 ? 1'h0 : _T_686; // @[Lookup.scala 11:37:@6700.4]
  assign _T_688 = _T_66 ? 1'h0 : _T_687; // @[Lookup.scala 11:37:@6701.4]
  assign _T_689 = _T_62 ? 1'h0 : _T_688; // @[Lookup.scala 11:37:@6702.4]
  assign _T_690 = _T_58 ? 1'h0 : _T_689; // @[Lookup.scala 11:37:@6703.4]
  assign _T_691 = _T_54 ? 1'h0 : _T_690; // @[Lookup.scala 11:37:@6704.4]
  assign _T_692 = _T_50 ? 1'h0 : _T_691; // @[Lookup.scala 11:37:@6705.4]
  assign _T_693 = _T_46 ? 1'h0 : _T_692; // @[Lookup.scala 11:37:@6706.4]
  assign _T_694 = _T_42 ? 1'h1 : _T_693; // @[Lookup.scala 11:37:@6707.4]
  assign _T_695 = _T_38 ? 1'h1 : _T_694; // @[Lookup.scala 11:37:@6708.4]
  assign _T_696 = _T_34 ? 1'h1 : _T_695; // @[Lookup.scala 11:37:@6709.4]
  assign _T_697 = _T_30 ? 1'h1 : _T_696; // @[Lookup.scala 11:37:@6710.4]
  assign _T_698 = _T_26 ? 1'h1 : _T_697; // @[Lookup.scala 11:37:@6711.4]
  assign _T_699 = _T_22 ? 1'h1 : _T_698; // @[Lookup.scala 11:37:@6712.4]
  assign _T_700 = _T_18 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:@6713.4]
  assign _T_744 = _T_38 ? 1'h1 : _T_42; // @[Lookup.scala 11:37:@6758.4]
  assign _T_745 = _T_34 ? 1'h1 : _T_744; // @[Lookup.scala 11:37:@6759.4]
  assign _T_746 = _T_30 ? 1'h0 : _T_745; // @[Lookup.scala 11:37:@6760.4]
  assign _T_747 = _T_26 ? 1'h0 : _T_746; // @[Lookup.scala 11:37:@6761.4]
  assign _T_748 = _T_22 ? 1'h0 : _T_747; // @[Lookup.scala 11:37:@6762.4]
  assign _T_749 = _T_18 ? 1'h0 : _T_748; // @[Lookup.scala 11:37:@6763.4]
  assign _T_792 = _T_42 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@6807.4]
  assign _T_793 = _T_38 ? 3'h1 : _T_792; // @[Lookup.scala 11:37:@6808.4]
  assign _T_794 = _T_34 ? 3'h3 : _T_793; // @[Lookup.scala 11:37:@6809.4]
  assign _T_795 = _T_30 ? 3'h6 : _T_794; // @[Lookup.scala 11:37:@6810.4]
  assign _T_796 = _T_26 ? 3'h2 : _T_795; // @[Lookup.scala 11:37:@6811.4]
  assign _T_797 = _T_22 ? 3'h5 : _T_796; // @[Lookup.scala 11:37:@6812.4]
  assign _T_798 = _T_18 ? 3'h1 : _T_797; // @[Lookup.scala 11:37:@6813.4]
  assign _T_802 = _T_198 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@6818.4]
  assign _T_803 = _T_194 ? 3'h4 : _T_802; // @[Lookup.scala 11:37:@6819.4]
  assign _T_804 = _T_190 ? 3'h4 : _T_803; // @[Lookup.scala 11:37:@6820.4]
  assign _T_805 = _T_186 ? 3'h4 : _T_804; // @[Lookup.scala 11:37:@6821.4]
  assign _T_806 = _T_182 ? 3'h3 : _T_805; // @[Lookup.scala 11:37:@6822.4]
  assign _T_807 = _T_178 ? 3'h3 : _T_806; // @[Lookup.scala 11:37:@6823.4]
  assign _T_808 = _T_174 ? 3'h2 : _T_807; // @[Lookup.scala 11:37:@6824.4]
  assign _T_809 = _T_170 ? 3'h1 : _T_808; // @[Lookup.scala 11:37:@6825.4]
  assign _T_810 = _T_166 ? 3'h2 : _T_809; // @[Lookup.scala 11:37:@6826.4]
  assign _T_811 = _T_162 ? 3'h1 : _T_810; // @[Lookup.scala 11:37:@6827.4]
  assign _T_812 = _T_158 ? 3'h0 : _T_811; // @[Lookup.scala 11:37:@6828.4]
  assign _T_813 = _T_154 ? 3'h0 : _T_812; // @[Lookup.scala 11:37:@6829.4]
  assign _T_814 = _T_150 ? 3'h0 : _T_813; // @[Lookup.scala 11:37:@6830.4]
  assign _T_815 = _T_146 ? 3'h0 : _T_814; // @[Lookup.scala 11:37:@6831.4]
  assign _T_816 = _T_142 ? 3'h0 : _T_815; // @[Lookup.scala 11:37:@6832.4]
  assign _T_817 = _T_138 ? 3'h0 : _T_816; // @[Lookup.scala 11:37:@6833.4]
  assign _T_818 = _T_134 ? 3'h0 : _T_817; // @[Lookup.scala 11:37:@6834.4]
  assign _T_819 = _T_130 ? 3'h0 : _T_818; // @[Lookup.scala 11:37:@6835.4]
  assign _T_820 = _T_126 ? 3'h0 : _T_819; // @[Lookup.scala 11:37:@6836.4]
  assign _T_821 = _T_122 ? 3'h0 : _T_820; // @[Lookup.scala 11:37:@6837.4]
  assign _T_822 = _T_118 ? 3'h0 : _T_821; // @[Lookup.scala 11:37:@6838.4]
  assign _T_823 = _T_114 ? 3'h0 : _T_822; // @[Lookup.scala 11:37:@6839.4]
  assign _T_824 = _T_110 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@6840.4]
  assign _T_825 = _T_106 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@6841.4]
  assign _T_826 = _T_102 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@6842.4]
  assign _T_827 = _T_98 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@6843.4]
  assign _T_828 = _T_94 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@6844.4]
  assign _T_829 = _T_90 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@6845.4]
  assign _T_830 = _T_86 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@6846.4]
  assign _T_831 = _T_82 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@6847.4]
  assign _T_832 = _T_78 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@6848.4]
  assign _T_833 = _T_74 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@6849.4]
  assign _T_834 = _T_70 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@6850.4]
  assign _T_835 = _T_66 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@6851.4]
  assign _T_836 = _T_62 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@6852.4]
  assign _T_837 = _T_58 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@6853.4]
  assign _T_838 = _T_54 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@6854.4]
  assign _T_839 = _T_50 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@6855.4]
  assign _T_840 = _T_46 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@6856.4]
  assign _T_841 = _T_42 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@6857.4]
  assign _T_842 = _T_38 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@6858.4]
  assign _T_843 = _T_34 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@6859.4]
  assign _T_844 = _T_30 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@6860.4]
  assign _T_845 = _T_26 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@6861.4]
  assign _T_846 = _T_22 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@6862.4]
  assign _T_847 = _T_18 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@6863.4]
  assign _T_850 = _T_202 ? 1'h0 : _T_206; // @[Lookup.scala 11:37:@6867.4]
  assign _T_851 = _T_198 ? 1'h0 : _T_850; // @[Lookup.scala 11:37:@6868.4]
  assign _T_852 = _T_194 ? 1'h0 : _T_851; // @[Lookup.scala 11:37:@6869.4]
  assign _T_853 = _T_190 ? 1'h0 : _T_852; // @[Lookup.scala 11:37:@6870.4]
  assign _T_854 = _T_186 ? 1'h0 : _T_853; // @[Lookup.scala 11:37:@6871.4]
  assign _T_855 = _T_182 ? 1'h0 : _T_854; // @[Lookup.scala 11:37:@6872.4]
  assign _T_856 = _T_178 ? 1'h0 : _T_855; // @[Lookup.scala 11:37:@6873.4]
  assign _T_857 = _T_174 ? 1'h0 : _T_856; // @[Lookup.scala 11:37:@6874.4]
  assign _T_858 = _T_170 ? 1'h0 : _T_857; // @[Lookup.scala 11:37:@6875.4]
  assign _T_859 = _T_166 ? 1'h0 : _T_858; // @[Lookup.scala 11:37:@6876.4]
  assign _T_860 = _T_162 ? 1'h0 : _T_859; // @[Lookup.scala 11:37:@6877.4]
  assign _T_861 = _T_158 ? 1'h0 : _T_860; // @[Lookup.scala 11:37:@6878.4]
  assign _T_862 = _T_154 ? 1'h0 : _T_861; // @[Lookup.scala 11:37:@6879.4]
  assign _T_863 = _T_150 ? 1'h0 : _T_862; // @[Lookup.scala 11:37:@6880.4]
  assign _T_864 = _T_146 ? 1'h0 : _T_863; // @[Lookup.scala 11:37:@6881.4]
  assign _T_865 = _T_142 ? 1'h0 : _T_864; // @[Lookup.scala 11:37:@6882.4]
  assign _T_866 = _T_138 ? 1'h0 : _T_865; // @[Lookup.scala 11:37:@6883.4]
  assign _T_867 = _T_134 ? 1'h0 : _T_866; // @[Lookup.scala 11:37:@6884.4]
  assign _T_868 = _T_130 ? 1'h0 : _T_867; // @[Lookup.scala 11:37:@6885.4]
  assign _T_869 = _T_126 ? 1'h0 : _T_868; // @[Lookup.scala 11:37:@6886.4]
  assign _T_870 = _T_122 ? 1'h0 : _T_869; // @[Lookup.scala 11:37:@6887.4]
  assign _T_871 = _T_118 ? 1'h0 : _T_870; // @[Lookup.scala 11:37:@6888.4]
  assign _T_872 = _T_114 ? 1'h0 : _T_871; // @[Lookup.scala 11:37:@6889.4]
  assign _T_873 = _T_110 ? 1'h0 : _T_872; // @[Lookup.scala 11:37:@6890.4]
  assign _T_874 = _T_106 ? 1'h0 : _T_873; // @[Lookup.scala 11:37:@6891.4]
  assign _T_875 = _T_102 ? 1'h0 : _T_874; // @[Lookup.scala 11:37:@6892.4]
  assign _T_876 = _T_98 ? 1'h0 : _T_875; // @[Lookup.scala 11:37:@6893.4]
  assign _T_877 = _T_94 ? 1'h0 : _T_876; // @[Lookup.scala 11:37:@6894.4]
  assign _T_878 = _T_90 ? 1'h0 : _T_877; // @[Lookup.scala 11:37:@6895.4]
  assign _T_879 = _T_86 ? 1'h0 : _T_878; // @[Lookup.scala 11:37:@6896.4]
  assign _T_880 = _T_82 ? 1'h0 : _T_879; // @[Lookup.scala 11:37:@6897.4]
  assign _T_881 = _T_78 ? 1'h0 : _T_880; // @[Lookup.scala 11:37:@6898.4]
  assign _T_882 = _T_74 ? 1'h0 : _T_881; // @[Lookup.scala 11:37:@6899.4]
  assign _T_883 = _T_70 ? 1'h0 : _T_882; // @[Lookup.scala 11:37:@6900.4]
  assign _T_884 = _T_66 ? 1'h0 : _T_883; // @[Lookup.scala 11:37:@6901.4]
  assign _T_885 = _T_62 ? 1'h0 : _T_884; // @[Lookup.scala 11:37:@6902.4]
  assign _T_886 = _T_58 ? 1'h0 : _T_885; // @[Lookup.scala 11:37:@6903.4]
  assign _T_887 = _T_54 ? 1'h0 : _T_886; // @[Lookup.scala 11:37:@6904.4]
  assign _T_888 = _T_50 ? 1'h0 : _T_887; // @[Lookup.scala 11:37:@6905.4]
  assign _T_889 = _T_46 ? 1'h0 : _T_888; // @[Lookup.scala 11:37:@6906.4]
  assign _T_890 = _T_42 ? 1'h0 : _T_889; // @[Lookup.scala 11:37:@6907.4]
  assign _T_891 = _T_38 ? 1'h0 : _T_890; // @[Lookup.scala 11:37:@6908.4]
  assign _T_892 = _T_34 ? 1'h0 : _T_891; // @[Lookup.scala 11:37:@6909.4]
  assign _T_893 = _T_30 ? 1'h0 : _T_892; // @[Lookup.scala 11:37:@6910.4]
  assign _T_894 = _T_26 ? 1'h0 : _T_893; // @[Lookup.scala 11:37:@6911.4]
  assign _T_895 = _T_22 ? 1'h0 : _T_894; // @[Lookup.scala 11:37:@6912.4]
  assign _T_896 = _T_18 ? 1'h0 : _T_895; // @[Lookup.scala 11:37:@6913.4]
  assign _T_899 = io_inst[19:15]; // @[InstDecoder.scala 131:31:@6930.4]
  assign _T_901 = io_inst[11:7]; // @[InstDecoder.scala 133:31:@6934.4]
  assign func = io_inst[6:2]; // @[InstDecoder.scala 135:21:@6936.4]
  assign _T_903 = func == 5'h18; // @[InstDecoder.scala 139:37:@6937.4]
  assign _T_905 = func == 5'h1b; // @[InstDecoder.scala 137:38:@6938.4]
  assign _T_906 = _T_903 | _T_905; // @[InstDecoder.scala 140:33:@6939.4]
  assign _T_915 = func == 5'h19; // @[InstDecoder.scala 138:39:@6946.4]
  assign _T_916 = _T_905 | _T_915; // @[InstDecoder.scala 142:34:@6947.4]
  assign _T_918 = io_cinfo_wbaddr == 5'h1; // @[InstDecoder.scala 136:37:@6948.4]
  assign _T_920 = io_cinfo_wbaddr == 5'h5; // @[InstDecoder.scala 136:53:@6949.4]
  assign _T_921 = _T_918 | _T_920; // @[InstDecoder.scala 136:45:@6950.4]
  assign _GEN_0 = {{4'd0}, _T_915}; // @[InstDecoder.scala 143:27:@6954.4]
  assign _T_925 = func == _GEN_0; // @[InstDecoder.scala 143:27:@6954.4]
  assign _T_927 = io_cinfo_rs1_addr == 5'h1; // @[InstDecoder.scala 136:37:@6955.4]
  assign _T_929 = io_cinfo_rs1_addr == 5'h5; // @[InstDecoder.scala 136:53:@6956.4]
  assign _T_930 = _T_927 | _T_929; // @[InstDecoder.scala 136:45:@6957.4]
  assign _T_931 = _T_925 & _T_930; // @[InstDecoder.scala 143:44:@6958.4]
  assign _T_938 = _T_921 == 1'h0; // @[InstDecoder.scala 144:6:@6962.4]
  assign _T_939 = io_cinfo_rs1_addr != io_cinfo_wbaddr; // @[InstDecoder.scala 144:50:@6963.4]
  assign _T_940 = _T_938 | _T_939; // @[InstDecoder.scala 144:29:@6964.4]
  assign imm_itype = io_inst[31:20]; // @[InstDecoder.scala 147:27:@6967.4]
  assign _T_942 = io_inst[31:25]; // @[InstDecoder.scala 148:31:@6968.4]
  assign imm_stype = {_T_942,_T_901}; // @[Cat.scala 30:58:@6970.4]
  assign _T_944 = io_inst[31]; // @[InstDecoder.scala 149:31:@6971.4]
  assign _T_945 = io_inst[7]; // @[InstDecoder.scala 149:44:@6972.4]
  assign _T_946 = io_inst[30:25]; // @[InstDecoder.scala 149:56:@6973.4]
  assign _T_947 = io_inst[11:8]; // @[InstDecoder.scala 149:73:@6974.4]
  assign imm_sbtype = {_T_944,_T_945,_T_946,_T_947}; // @[Cat.scala 30:58:@6977.4]
  assign imm_utype = io_inst[31:12]; // @[InstDecoder.scala 150:27:@6978.4]
  assign _T_951 = io_inst[19:12]; // @[InstDecoder.scala 151:44:@6980.4]
  assign _T_952 = io_inst[20]; // @[InstDecoder.scala 151:60:@6981.4]
  assign _T_953 = io_inst[30:21]; // @[InstDecoder.scala 151:73:@6982.4]
  assign imm_ujtype = {_T_944,_T_951,_T_952,_T_953}; // @[Cat.scala 30:58:@6985.4]
  assign _T_956 = imm_itype[11]; // @[InstDecoder.scala 154:43:@6986.4]
  assign _T_960 = _T_956 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@6988.4]
  assign _T_962 = imm_stype[11]; // @[InstDecoder.scala 155:43:@6991.4]
  assign _T_966 = _T_962 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@6993.4]
  assign _T_968 = imm_sbtype[11]; // @[InstDecoder.scala 156:44:@6996.4]
  assign _T_972 = _T_968 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@6998.4]
  assign _T_974 = {_T_972,_T_944,_T_945,_T_946,_T_947}; // @[Cat.scala 30:58:@6999.4]
  assign _T_982 = imm_ujtype[19]; // @[InstDecoder.scala 158:44:@7005.4]
  assign _T_986 = _T_982 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@7007.4]
  assign _T_988 = {_T_986,_T_944,_T_951,_T_952,_T_953}; // @[Cat.scala 30:58:@7008.4]
  assign io_cinfo_br_type = _T_14 ? 4'h0 : _T_308; // @[InstDecoder.scala 116:20:@6915.4]
  assign io_cinfo_op1_sel = _T_14 ? 2'h0 : _T_357; // @[InstDecoder.scala 117:20:@6916.4]
  assign io_cinfo_op2_sel = _T_14 ? 3'h1 : _T_406; // @[InstDecoder.scala 118:20:@6917.4]
  assign io_cinfo_rs1_oen = _T_14 ? 1'h1 : _T_455; // @[InstDecoder.scala 119:20:@6918.4]
  assign io_cinfo_rs2_oen = _T_14 ? 1'h0 : _T_504; // @[InstDecoder.scala 120:20:@6919.4]
  assign io_cinfo_alu_fun = _T_14 ? 4'h0 : _T_553; // @[InstDecoder.scala 121:20:@6920.4]
  assign io_cinfo_wb_sel = _T_14 ? 2'h1 : _T_602; // @[InstDecoder.scala 122:20:@6921.4]
  assign io_cinfo_rf_wen = _T_14 ? 1'h1 : _T_651; // @[InstDecoder.scala 123:20:@6922.4]
  assign io_cinfo_mem_en = _T_14 ? 1'h1 : _T_700; // @[InstDecoder.scala 124:20:@6923.4]
  assign io_cinfo_mem_fcn = _T_14 ? 1'h0 : _T_749; // @[InstDecoder.scala 125:20:@6924.4]
  assign io_cinfo_mem_typ = _T_14 ? 3'h3 : _T_798; // @[InstDecoder.scala 126:20:@6925.4]
  assign io_cinfo_csr_cmd = _T_14 ? 3'h0 : _T_847; // @[InstDecoder.scala 127:20:@6926.4]
  assign io_cinfo_illegal = signals_0 == 1'h0; // @[InstDecoder.scala 128:20:@6928.4]
  assign io_cinfo_fencei = _T_14 ? 1'h0 : _T_896; // @[InstDecoder.scala 129:20:@6929.4]
  assign io_cinfo_branch = func == 5'h18; // @[InstDecoder.scala 141:19:@6944.4]
  assign io_cinfo_push = _T_916 & _T_921; // @[InstDecoder.scala 142:19:@6952.4]
  assign io_cinfo_pop = _T_931 & _T_940; // @[InstDecoder.scala 143:19:@6966.4]
  assign io_cinfo_isBJ = _T_906 | _T_905; // @[InstDecoder.scala 140:19:@6942.4]
  assign io_cinfo_rs1_addr = io_inst[19:15]; // @[InstDecoder.scala 131:21:@6931.4]
  assign io_cinfo_rs2_addr = io_inst[24:20]; // @[InstDecoder.scala 132:21:@6933.4]
  assign io_cinfo_wbaddr = io_inst[11:7]; // @[InstDecoder.scala 133:21:@6935.4]
  assign io_dinfo_imm_i = {_T_960,imm_itype}; // @[InstDecoder.scala 154:19:@6990.4]
  assign io_dinfo_imm_s = {_T_966,imm_stype}; // @[InstDecoder.scala 155:19:@6995.4]
  assign io_dinfo_imm_sb = {_T_974,1'h0}; // @[InstDecoder.scala 156:19:@7001.4]
  assign io_dinfo_imm_u = {imm_utype,12'h0}; // @[InstDecoder.scala 157:19:@7004.4]
  assign io_dinfo_imm_uj = {_T_988,1'h0}; // @[InstDecoder.scala 158:19:@7010.4]
  assign io_dinfo_imm_z = {27'h0,_T_899}; // @[InstDecoder.scala 159:19:@7014.4]
endmodule
module BackEnd( // @[:@7922.2]
  input         clock, // @[:@7923.4]
  input         reset, // @[:@7924.4]
  output        io_mem_req_valid, // @[:@7925.4]
  output [31:0] io_mem_req_bits_addr, // @[:@7925.4]
  output [31:0] io_mem_req_bits_data, // @[:@7925.4]
  output        io_mem_req_bits_fcn, // @[:@7925.4]
  output [2:0]  io_mem_req_bits_typ, // @[:@7925.4]
  input         io_mem_resp_valid, // @[:@7925.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@7925.4]
  output [31:0] io_cyc, // @[:@7925.4]
  output        io_front_xcpt_valid, // @[:@7925.4]
  output [31:0] io_front_xcpt_bits, // @[:@7925.4]
  output        io_front_kill, // @[:@7925.4]
  output        io_front_fence, // @[:@7925.4]
  output        io_front_ras_pop, // @[:@7925.4]
  output        io_front_ras_push_valid, // @[:@7925.4]
  output [31:0] io_front_ras_push_bits, // @[:@7925.4]
  output [31:0] io_front_fb_pc, // @[:@7925.4]
  output [1:0]  io_front_fb_type, // @[:@7925.4]
  output        io_front_feedBack_valid, // @[:@7925.4]
  output        io_front_feedBack_bits_redirect, // @[:@7925.4]
  output [31:0] io_front_feedBack_bits_tgt, // @[:@7925.4]
  output        io_front_forward_0, // @[:@7925.4]
  output        io_front_forward_1, // @[:@7925.4]
  input         io_front_inst_0_valid, // @[:@7925.4]
  input  [31:0] io_front_inst_0_bits, // @[:@7925.4]
  input         io_front_inst_1_valid, // @[:@7925.4]
  input  [31:0] io_front_inst_1_bits, // @[:@7925.4]
  input  [31:0] io_front_pc_0, // @[:@7925.4]
  input  [31:0] io_front_pc_1, // @[:@7925.4]
  input  [31:0] io_front_pred_0, // @[:@7925.4]
  input  [31:0] io_front_pred_1 // @[:@7925.4]
);
  wire  csr_clock; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_reset; // @[BackEnd.scala 80:19:@7927.4]
  wire [2:0] csr_io_rw_cmd; // @[BackEnd.scala 80:19:@7927.4]
  wire [11:0] csr_io_rw_addr; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_rw_rdata; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_rw_wdata; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_eret; // @[BackEnd.scala 80:19:@7927.4]
  wire [1:0] csr_io_status_prv; // @[BackEnd.scala 80:19:@7927.4]
  wire [13:0] csr_io_status_unimp5; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_status_mprv; // @[BackEnd.scala 80:19:@7927.4]
  wire [1:0] csr_io_status_unimp4; // @[BackEnd.scala 80:19:@7927.4]
  wire [1:0] csr_io_status_mpp; // @[BackEnd.scala 80:19:@7927.4]
  wire [2:0] csr_io_status_unimp3; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_status_mpie; // @[BackEnd.scala 80:19:@7927.4]
  wire [2:0] csr_io_status_unimp2; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_status_mie; // @[BackEnd.scala 80:19:@7927.4]
  wire [2:0] csr_io_status_unimp1; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_xcpt; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_cause; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_tval; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_evec; // @[BackEnd.scala 80:19:@7927.4]
  wire  csr_io_illegal; // @[BackEnd.scala 80:19:@7927.4]
  wire [1:0] csr_io_retire; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_pc; // @[BackEnd.scala 80:19:@7927.4]
  wire [31:0] csr_io_time; // @[BackEnd.scala 80:19:@7927.4]
  wire  regfile_clock; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_rs1_addr_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_rs1_addr_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_rs1_data_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_rs1_data_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_rs2_addr_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_rs2_addr_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_rs2_data_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_rs2_data_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_waddr_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [4:0] regfile_io_waddr_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_wdata_0; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] regfile_io_wdata_1; // @[BackEnd.scala 81:23:@7930.4]
  wire  regfile_io_wen_0; // @[BackEnd.scala 81:23:@7930.4]
  wire  regfile_io_wen_1; // @[BackEnd.scala 81:23:@7930.4]
  wire [31:0] ALU_io_op1; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_op2; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_pc; // @[BackEnd.scala 82:33:@7933.4]
  wire [3:0] ALU_io_ctrl_fun; // @[BackEnd.scala 82:33:@7933.4]
  wire [3:0] ALU_io_ctrl_br_type; // @[BackEnd.scala 82:33:@7933.4]
  wire [1:0] ALU_io_ctrl_wb_sel; // @[BackEnd.scala 82:33:@7933.4]
  wire [1:0] ALU_io_ctrl_pc_sel; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_rs2_data; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_result; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_target_brjmp; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_target_jpreg; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_io_target_conti; // @[BackEnd.scala 82:33:@7933.4]
  wire [31:0] ALU_1_io_op1; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_op2; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_pc; // @[BackEnd.scala 82:33:@7936.4]
  wire [3:0] ALU_1_io_ctrl_fun; // @[BackEnd.scala 82:33:@7936.4]
  wire [3:0] ALU_1_io_ctrl_br_type; // @[BackEnd.scala 82:33:@7936.4]
  wire [1:0] ALU_1_io_ctrl_wb_sel; // @[BackEnd.scala 82:33:@7936.4]
  wire [1:0] ALU_1_io_ctrl_pc_sel; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_rs2_data; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_result; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_target_brjmp; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_target_jpreg; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] ALU_1_io_target_conti; // @[BackEnd.scala 82:33:@7936.4]
  wire [31:0] InstDecoder_io_inst; // @[BackEnd.scala 83:33:@7939.4]
  wire [3:0] InstDecoder_io_cinfo_br_type; // @[BackEnd.scala 83:33:@7939.4]
  wire [1:0] InstDecoder_io_cinfo_op1_sel; // @[BackEnd.scala 83:33:@7939.4]
  wire [2:0] InstDecoder_io_cinfo_op2_sel; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 83:33:@7939.4]
  wire [3:0] InstDecoder_io_cinfo_alu_fun; // @[BackEnd.scala 83:33:@7939.4]
  wire [1:0] InstDecoder_io_cinfo_wb_sel; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_mem_en; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_mem_fcn; // @[BackEnd.scala 83:33:@7939.4]
  wire [2:0] InstDecoder_io_cinfo_mem_typ; // @[BackEnd.scala 83:33:@7939.4]
  wire [2:0] InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_illegal; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_fencei; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_branch; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_push; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_pop; // @[BackEnd.scala 83:33:@7939.4]
  wire  InstDecoder_io_cinfo_isBJ; // @[BackEnd.scala 83:33:@7939.4]
  wire [4:0] InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 83:33:@7939.4]
  wire [4:0] InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 83:33:@7939.4]
  wire [4:0] InstDecoder_io_cinfo_wbaddr; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_i; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_s; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_sb; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_u; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_uj; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_io_dinfo_imm_z; // @[BackEnd.scala 83:33:@7939.4]
  wire [31:0] InstDecoder_1_io_inst; // @[BackEnd.scala 83:33:@7942.4]
  wire [3:0] InstDecoder_1_io_cinfo_br_type; // @[BackEnd.scala 83:33:@7942.4]
  wire [1:0] InstDecoder_1_io_cinfo_op1_sel; // @[BackEnd.scala 83:33:@7942.4]
  wire [2:0] InstDecoder_1_io_cinfo_op2_sel; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_rs1_oen; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_rs2_oen; // @[BackEnd.scala 83:33:@7942.4]
  wire [3:0] InstDecoder_1_io_cinfo_alu_fun; // @[BackEnd.scala 83:33:@7942.4]
  wire [1:0] InstDecoder_1_io_cinfo_wb_sel; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_rf_wen; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_mem_en; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_mem_fcn; // @[BackEnd.scala 83:33:@7942.4]
  wire [2:0] InstDecoder_1_io_cinfo_mem_typ; // @[BackEnd.scala 83:33:@7942.4]
  wire [2:0] InstDecoder_1_io_cinfo_csr_cmd; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_illegal; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_fencei; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_branch; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_push; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_pop; // @[BackEnd.scala 83:33:@7942.4]
  wire  InstDecoder_1_io_cinfo_isBJ; // @[BackEnd.scala 83:33:@7942.4]
  wire [4:0] InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 83:33:@7942.4]
  wire [4:0] InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 83:33:@7942.4]
  wire [4:0] InstDecoder_1_io_cinfo_wbaddr; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_i; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_s; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_sb; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_u; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_uj; // @[BackEnd.scala 83:33:@7942.4]
  wire [31:0] InstDecoder_1_io_dinfo_imm_z; // @[BackEnd.scala 83:33:@7942.4]
  reg  exe_0_rf_wen; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_0;
  reg [4:0] exe_0_wbaddr; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_1;
  reg  exe_0_mem_en; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_2;
  reg [2:0] exe_0_csr_cmd; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_3;
  reg  exe_0_illegal; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_4;
  reg [31:0] exe_0_pc; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_5;
  reg [31:0] exe_0_inst; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_6;
  reg [31:0] exe_0_rs2_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_7;
  reg [1:0] exe_0_wb_sel; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_8;
  reg  exe_0_mem_fcn; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_9;
  reg [2:0] exe_0_mem_typ; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_10;
  reg  exe_0_fencei; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_11;
  reg [3:0] exe_0_br_type; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_12;
  reg  exe_0_isBJ; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_13;
  reg [31:0] exe_0_op1_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_14;
  reg [31:0] exe_0_op2_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_15;
  reg [3:0] exe_0_alu_fun; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_16;
  reg  exe_1_rf_wen; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_17;
  reg [4:0] exe_1_wbaddr; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_18;
  reg  exe_1_mem_en; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_19;
  reg [2:0] exe_1_csr_cmd; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_20;
  reg  exe_1_illegal; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_21;
  reg [31:0] exe_1_pc; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_22;
  reg [31:0] exe_1_inst; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_23;
  reg [31:0] exe_1_rs2_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_24;
  reg [1:0] exe_1_wb_sel; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_25;
  reg  exe_1_mem_fcn; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_26;
  reg [2:0] exe_1_mem_typ; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_27;
  reg  exe_1_fencei; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_28;
  reg [3:0] exe_1_br_type; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_29;
  reg  exe_1_isBJ; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_30;
  reg [31:0] exe_1_op1_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_31;
  reg [31:0] exe_1_op2_data; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_32;
  reg [3:0] exe_1_alu_fun; // @[BackEnd.scala 90:22:@7950.4]
  reg [31:0] _RAND_33;
  reg  exe_valid_0; // @[BackEnd.scala 91:26:@7954.4]
  reg [31:0] _RAND_34;
  reg  exe_valid_1; // @[BackEnd.scala 91:26:@7954.4]
  reg [31:0] _RAND_35;
  reg  mem_0_rf_wen; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_36;
  reg [4:0] mem_0_wbaddr; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_37;
  reg  mem_0_mem_en; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_38;
  reg [2:0] mem_0_csr_cmd; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_39;
  reg  mem_0_illegal; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_40;
  reg [31:0] mem_0_pc; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_41;
  reg [31:0] mem_0_inst; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_42;
  reg [1:0] mem_0_wb_sel; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_43;
  reg  mem_0_mem_fcn; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_44;
  reg [2:0] mem_0_mem_typ; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_45;
  reg  mem_1_rf_wen; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_46;
  reg [4:0] mem_1_wbaddr; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_47;
  reg  mem_1_mem_en; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_48;
  reg [2:0] mem_1_csr_cmd; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_49;
  reg  mem_1_illegal; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_50;
  reg [31:0] mem_1_pc; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_51;
  reg [31:0] mem_1_inst; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_52;
  reg [1:0] mem_1_wb_sel; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_53;
  reg  mem_1_mem_fcn; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_54;
  reg [2:0] mem_1_mem_typ; // @[BackEnd.scala 93:22:@7956.4]
  reg [31:0] _RAND_55;
  reg  mem_valid_0; // @[BackEnd.scala 94:26:@7960.4]
  reg [31:0] _RAND_56;
  reg  mem_valid_1; // @[BackEnd.scala 94:26:@7960.4]
  reg [31:0] _RAND_57;
  reg  wb_0_rf_wen; // @[BackEnd.scala 96:22:@7962.4]
  reg [31:0] _RAND_58;
  reg [4:0] wb_0_wbaddr; // @[BackEnd.scala 96:22:@7962.4]
  reg [31:0] _RAND_59;
  reg  wb_1_rf_wen; // @[BackEnd.scala 96:22:@7962.4]
  reg [31:0] _RAND_60;
  reg [4:0] wb_1_wbaddr; // @[BackEnd.scala 96:22:@7962.4]
  reg [31:0] _RAND_61;
  reg  wb_valid_0; // @[BackEnd.scala 97:26:@7966.4]
  reg [31:0] _RAND_62;
  reg  wb_valid_1; // @[BackEnd.scala 97:26:@7966.4]
  reg [31:0] _RAND_63;
  wire  dec_wire_0_fencei; // @[BackEnd.scala 120:51:@7992.4]
  wire  dec_wire_1_fencei; // @[BackEnd.scala 120:51:@8093.4]
  wire  _T_473; // @[BackEnd.scala 100:54:@7968.4]
  wire  exe_wire_0_fencei; // @[BackEnd.scala 211:41:@8247.4]
  wire  exe_wire_1_fencei; // @[BackEnd.scala 211:41:@8286.4]
  wire  _T_474; // @[BackEnd.scala 100:93:@7969.4]
  reg [31:0] wb_wbdata_0; // @[BackEnd.scala 104:23:@7974.4]
  reg [31:0] _RAND_64;
  reg [31:0] wb_wbdata_1; // @[BackEnd.scala 104:23:@7974.4]
  reg [31:0] _RAND_65;
  wire  dec_wire_0_rs1_oen; // @[BackEnd.scala 116:51:@7982.4]
  wire  dec_wire_0_rs2_oen; // @[BackEnd.scala 117:51:@7984.4]
  wire  _T_541; // @[BackEnd.scala 118:51:@7986.4]
  wire  _T_543; // @[BackEnd.scala 118:97:@7987.4]
  wire  dec_wire_0_rf_wen; // @[BackEnd.scala 118:74:@7988.4]
  wire  dec_wire_0_isBJ; // @[BackEnd.scala 119:51:@7990.4]
  wire [2:0] dec_wire_0_csr_cmd; // @[BackEnd.scala 121:31:@7994.4]
  wire  _T_548; // @[BackEnd.scala 129:23:@8000.4]
  wire  _T_749; // @[BackEnd.scala 208:41:@8278.4]
  wire  _T_751; // @[BackEnd.scala 208:75:@8279.4]
  wire  exe_wire_1_rf_wen; // @[BackEnd.scala 208:58:@8280.4]
  wire  _T_549; // @[BackEnd.scala 129:50:@8001.4]
  wire  _T_550; // @[BackEnd.scala 130:23:@8002.4]
  wire  _T_737; // @[BackEnd.scala 208:41:@8239.4]
  wire  _T_739; // @[BackEnd.scala 208:75:@8240.4]
  wire  exe_wire_0_rf_wen; // @[BackEnd.scala 208:58:@8241.4]
  wire  _T_551; // @[BackEnd.scala 130:50:@8003.4]
  wire  _T_552; // @[BackEnd.scala 131:23:@8004.4]
  wire  _T_876; // @[BackEnd.scala 300:41:@8457.4]
  wire  _T_878; // @[BackEnd.scala 300:75:@8458.4]
  wire  mem_wire_1_rf_wen; // @[BackEnd.scala 300:58:@8459.4]
  wire  _T_553; // @[BackEnd.scala 131:50:@8005.4]
  wire  _T_554; // @[BackEnd.scala 132:23:@8006.4]
  wire  _T_857; // @[BackEnd.scala 300:41:@8429.4]
  wire  _T_859; // @[BackEnd.scala 300:75:@8430.4]
  wire  mem_wire_0_rf_wen; // @[BackEnd.scala 300:58:@8431.4]
  wire  _T_555; // @[BackEnd.scala 132:50:@8007.4]
  wire  _T_556; // @[BackEnd.scala 133:23:@8008.4]
  wire  _T_941; // @[BackEnd.scala 373:40:@8646.4]
  wire  _T_943; // @[BackEnd.scala 373:72:@8647.4]
  wire  wb_wire_1_rf_wen; // @[BackEnd.scala 373:56:@8648.4]
  wire  _T_557; // @[BackEnd.scala 133:50:@8009.4]
  wire  _T_558; // @[BackEnd.scala 134:23:@8010.4]
  wire  _T_937; // @[BackEnd.scala 373:40:@8639.4]
  wire  _T_939; // @[BackEnd.scala 373:72:@8640.4]
  wire  wb_wire_0_rf_wen; // @[BackEnd.scala 373:56:@8641.4]
  wire  _T_559; // @[BackEnd.scala 134:50:@8011.4]
  wire [31:0] rf_rs1_data_0; // @[BackEnd.scala 112:25:@7979.4 BackEnd.scala 125:20:@7998.4]
  wire [31:0] _T_560; // @[Mux.scala 61:16:@8012.4]
  wire [31:0] _T_561; // @[Mux.scala 61:16:@8013.4]
  wire  _T_872; // @[BackEnd.scala 312:22:@8448.4]
  wire  _T_873; // @[BackEnd.scala 313:22:@8449.4]
  reg [31:0] mem_reg_wbdata_0; // @[BackEnd.scala 206:28:@8238.4]
  reg [31:0] _RAND_66;
  wire [31:0] _T_874; // @[Mux.scala 61:16:@8450.4]
  wire [31:0] mem_wbdata_0; // @[Mux.scala 61:16:@8451.4]
  wire [31:0] _T_562; // @[Mux.scala 61:16:@8014.4]
  wire  _T_891; // @[BackEnd.scala 312:22:@8476.4]
  wire  _T_892; // @[BackEnd.scala 313:22:@8477.4]
  reg [31:0] mem_reg_wbdata_1; // @[BackEnd.scala 206:28:@8238.4]
  reg [31:0] _RAND_67;
  wire [31:0] _T_893; // @[Mux.scala 61:16:@8478.4]
  wire [31:0] mem_wbdata_1; // @[Mux.scala 61:16:@8479.4]
  wire [31:0] _T_563; // @[Mux.scala 61:16:@8015.4]
  wire [31:0] exe_wbdata_0; // @[BackEnd.scala 102:24:@7972.4 BackEnd.scala 224:19:@8262.4]
  wire [31:0] _T_564; // @[Mux.scala 61:16:@8016.4]
  wire [31:0] exe_wbdata_1; // @[BackEnd.scala 102:24:@7972.4 BackEnd.scala 224:19:@8301.4]
  wire [31:0] dec_rs1_data_0; // @[Mux.scala 61:16:@8017.4]
  wire  _T_566; // @[BackEnd.scala 138:23:@8019.4]
  wire  _T_567; // @[BackEnd.scala 138:50:@8020.4]
  wire  _T_568; // @[BackEnd.scala 139:23:@8021.4]
  wire  _T_569; // @[BackEnd.scala 139:50:@8022.4]
  wire  _T_570; // @[BackEnd.scala 140:23:@8023.4]
  wire  _T_571; // @[BackEnd.scala 140:50:@8024.4]
  wire  _T_572; // @[BackEnd.scala 141:23:@8025.4]
  wire  _T_573; // @[BackEnd.scala 141:50:@8026.4]
  wire  _T_574; // @[BackEnd.scala 142:23:@8027.4]
  wire  _T_575; // @[BackEnd.scala 142:50:@8028.4]
  wire  _T_576; // @[BackEnd.scala 143:23:@8029.4]
  wire  _T_577; // @[BackEnd.scala 143:50:@8030.4]
  wire [31:0] rf_rs2_data_0; // @[BackEnd.scala 113:25:@7980.4 BackEnd.scala 126:20:@7999.4]
  wire [31:0] _T_578; // @[Mux.scala 61:16:@8031.4]
  wire [31:0] _T_579; // @[Mux.scala 61:16:@8032.4]
  wire [31:0] _T_580; // @[Mux.scala 61:16:@8033.4]
  wire [31:0] _T_581; // @[Mux.scala 61:16:@8034.4]
  wire [31:0] _T_582; // @[Mux.scala 61:16:@8035.4]
  wire [31:0] dec_rs2_data_0; // @[Mux.scala 61:16:@8036.4]
  wire  _T_584; // @[BackEnd.scala 147:29:@8038.4]
  wire  _T_585; // @[BackEnd.scala 148:29:@8039.4]
  wire [31:0] _T_586; // @[Mux.scala 61:16:@8040.4]
  wire [31:0] dec_op1_data_0; // @[Mux.scala 61:16:@8041.4]
  wire  _T_588; // @[BackEnd.scala 151:29:@8043.4]
  wire  _T_589; // @[BackEnd.scala 152:29:@8044.4]
  wire  _T_590; // @[BackEnd.scala 153:29:@8045.4]
  wire  _T_591; // @[BackEnd.scala 154:29:@8046.4]
  wire  _T_592; // @[BackEnd.scala 155:29:@8047.4]
  wire [31:0] _T_593; // @[Mux.scala 61:16:@8048.4]
  wire [31:0] _T_594; // @[Mux.scala 61:16:@8049.4]
  wire [31:0] _T_595; // @[Mux.scala 61:16:@8050.4]
  wire [31:0] _T_596; // @[Mux.scala 61:16:@8051.4]
  wire [31:0] dec_op2_data_0; // @[Mux.scala 61:16:@8052.4]
  wire  exe_wire_0_mem_en; // @[BackEnd.scala 209:41:@8243.4]
  wire  exe_wire_1_mem_en; // @[BackEnd.scala 209:41:@8282.4]
  wire  stall_1_1; // @[BackEnd.scala 415:80:@8801.4]
  wire  _T_599; // @[BackEnd.scala 157:11:@8054.4]
  wire [2:0] mem_wire_1_csr_cmd; // @[BackEnd.scala 302:31:@8463.4]
  wire  _T_887; // @[BackEnd.scala 306:39:@8471.4]
  wire  mem_wire_1_mem_en; // @[BackEnd.scala 301:41:@8461.4]
  wire  _T_888; // @[BackEnd.scala 306:49:@8472.4]
  wire  mem_wire_1_illegal; // @[BackEnd.scala 303:41:@8465.4]
  wire  _T_889; // @[BackEnd.scala 307:39:@8473.4]
  reg [31:0] mem_reg_jpnpc; // @[BackEnd.scala 270:31:@8376.4]
  reg [31:0] _RAND_68;
  wire [1:0] _T_883; // @[BackEnd.scala 304:54:@8467.4]
  wire  _T_885; // @[BackEnd.scala 304:60:@8468.4]
  wire  mem_wire_jump_1; // @[BackEnd.scala 304:38:@8469.4]
  wire  mem_sel_1; // @[BackEnd.scala 308:39:@8474.4]
  wire [2:0] mem_wire_0_csr_cmd; // @[BackEnd.scala 302:31:@8435.4]
  wire  _T_868; // @[BackEnd.scala 306:39:@8443.4]
  wire  mem_wire_0_mem_en; // @[BackEnd.scala 301:41:@8433.4]
  wire  _T_869; // @[BackEnd.scala 306:49:@8444.4]
  wire  mem_wire_0_illegal; // @[BackEnd.scala 303:41:@8437.4]
  wire  _T_870; // @[BackEnd.scala 307:39:@8445.4]
  wire  mem_wire_jump_0; // @[BackEnd.scala 304:38:@8441.4]
  wire  mem_sel_0; // @[BackEnd.scala 308:39:@8446.4]
  wire [1:0] _T_1120; // @[BackEnd.scala 417:34:@8807.4]
  wire [1:0] _T_1121; // @[BackEnd.scala 417:41:@8808.4]
  wire  _T_1123; // @[BackEnd.scala 417:41:@8809.4]
  wire  _T_1125; // @[BackEnd.scala 417:72:@8810.4]
  wire  _T_1126; // @[BackEnd.scala 417:69:@8811.4]
  wire  _T_1127; // @[BackEnd.scala 417:46:@8812.4]
  wire  stall_0_2; // @[BackEnd.scala 416:45:@8805.4]
  wire  stall_1_2; // @[BackEnd.scala 417:92:@8813.4]
  wire  _T_601; // @[BackEnd.scala 157:35:@8055.4]
  wire  _T_602; // @[BackEnd.scala 157:32:@8056.4]
  wire  _T_603; // @[BackEnd.scala 161:52:@8060.6]
  wire  _T_604; // @[BackEnd.scala 161:86:@8061.6]
  wire  _T_605; // @[BackEnd.scala 161:62:@8062.6]
  wire  _T_607; // @[BackEnd.scala 162:53:@8063.6]
  wire  _T_608; // @[BackEnd.scala 161:97:@8064.6]
  wire [2:0] _T_609; // @[BackEnd.scala 161:29:@8065.6]
  wire  dec_wire_1_rs1_oen; // @[BackEnd.scala 116:51:@8083.4]
  wire  dec_wire_1_rs2_oen; // @[BackEnd.scala 117:51:@8085.4]
  wire  dec_wire_1_isBJ; // @[BackEnd.scala 119:51:@8091.4]
  wire  _T_619; // @[BackEnd.scala 129:23:@8101.4]
  wire  _T_620; // @[BackEnd.scala 129:50:@8102.4]
  wire  _T_621; // @[BackEnd.scala 130:23:@8103.4]
  wire  _T_622; // @[BackEnd.scala 130:50:@8104.4]
  wire  _T_623; // @[BackEnd.scala 131:23:@8105.4]
  wire  _T_624; // @[BackEnd.scala 131:50:@8106.4]
  wire  _T_625; // @[BackEnd.scala 132:23:@8107.4]
  wire  _T_626; // @[BackEnd.scala 132:50:@8108.4]
  wire  _T_627; // @[BackEnd.scala 133:23:@8109.4]
  wire  _T_628; // @[BackEnd.scala 133:50:@8110.4]
  wire  _T_629; // @[BackEnd.scala 134:23:@8111.4]
  wire  _T_630; // @[BackEnd.scala 134:50:@8112.4]
  wire [31:0] rf_rs1_data_1; // @[BackEnd.scala 112:25:@7979.4 BackEnd.scala 125:20:@8099.4]
  wire [31:0] _T_631; // @[Mux.scala 61:16:@8113.4]
  wire [31:0] _T_632; // @[Mux.scala 61:16:@8114.4]
  wire [31:0] _T_633; // @[Mux.scala 61:16:@8115.4]
  wire [31:0] _T_634; // @[Mux.scala 61:16:@8116.4]
  wire [31:0] _T_635; // @[Mux.scala 61:16:@8117.4]
  wire [31:0] dec_rs1_data_1; // @[Mux.scala 61:16:@8118.4]
  wire  _T_637; // @[BackEnd.scala 138:23:@8120.4]
  wire  _T_638; // @[BackEnd.scala 138:50:@8121.4]
  wire  _T_639; // @[BackEnd.scala 139:23:@8122.4]
  wire  _T_640; // @[BackEnd.scala 139:50:@8123.4]
  wire  _T_641; // @[BackEnd.scala 140:23:@8124.4]
  wire  _T_642; // @[BackEnd.scala 140:50:@8125.4]
  wire  _T_643; // @[BackEnd.scala 141:23:@8126.4]
  wire  _T_644; // @[BackEnd.scala 141:50:@8127.4]
  wire  _T_645; // @[BackEnd.scala 142:23:@8128.4]
  wire  _T_646; // @[BackEnd.scala 142:50:@8129.4]
  wire  _T_647; // @[BackEnd.scala 143:23:@8130.4]
  wire  _T_648; // @[BackEnd.scala 143:50:@8131.4]
  wire [31:0] rf_rs2_data_1; // @[BackEnd.scala 113:25:@7980.4 BackEnd.scala 126:20:@8100.4]
  wire [31:0] _T_649; // @[Mux.scala 61:16:@8132.4]
  wire [31:0] _T_650; // @[Mux.scala 61:16:@8133.4]
  wire [31:0] _T_651; // @[Mux.scala 61:16:@8134.4]
  wire [31:0] _T_652; // @[Mux.scala 61:16:@8135.4]
  wire [31:0] _T_653; // @[Mux.scala 61:16:@8136.4]
  wire [31:0] dec_rs2_data_1; // @[Mux.scala 61:16:@8137.4]
  wire  _T_655; // @[BackEnd.scala 147:29:@8139.4]
  wire  _T_656; // @[BackEnd.scala 148:29:@8140.4]
  wire [31:0] _T_657; // @[Mux.scala 61:16:@8141.4]
  wire [31:0] dec_op1_data_1; // @[Mux.scala 61:16:@8142.4]
  wire  _T_659; // @[BackEnd.scala 151:29:@8144.4]
  wire  _T_660; // @[BackEnd.scala 152:29:@8145.4]
  wire  _T_661; // @[BackEnd.scala 153:29:@8146.4]
  wire  _T_662; // @[BackEnd.scala 154:29:@8147.4]
  wire  _T_663; // @[BackEnd.scala 155:29:@8148.4]
  wire [31:0] _T_664; // @[Mux.scala 61:16:@8149.4]
  wire [31:0] _T_665; // @[Mux.scala 61:16:@8150.4]
  wire [31:0] _T_666; // @[Mux.scala 61:16:@8151.4]
  wire [31:0] _T_667; // @[Mux.scala 61:16:@8152.4]
  wire [31:0] dec_op2_data_1; // @[Mux.scala 61:16:@8153.4]
  wire  _T_674; // @[BackEnd.scala 161:52:@8161.6]
  wire  _T_675; // @[BackEnd.scala 161:86:@8162.6]
  wire  _T_676; // @[BackEnd.scala 161:62:@8163.6]
  wire  _T_678; // @[BackEnd.scala 162:53:@8164.6]
  wire  _T_679; // @[BackEnd.scala 161:97:@8165.6]
  wire [2:0] _T_680; // @[BackEnd.scala 161:29:@8166.6]
  reg [31:0] exe_pred_tgt; // @[BackEnd.scala 179:27:@8183.4]
  reg [31:0] _RAND_69;
  reg  exe_reg_branch; // @[BackEnd.scala 180:27:@8184.4]
  reg [31:0] _RAND_70;
  reg  exe_reg_pop; // @[BackEnd.scala 181:27:@8185.4]
  reg [31:0] _RAND_71;
  reg  exe_reg_push; // @[BackEnd.scala 182:27:@8186.4]
  reg [31:0] _RAND_72;
  wire [31:0] _T_690; // @[BackEnd.scala 184:26:@8191.6]
  wire  _T_691; // @[BackEnd.scala 185:26:@8193.6]
  wire  _T_692; // @[BackEnd.scala 186:26:@8195.6]
  wire  _T_693; // @[BackEnd.scala 187:26:@8197.6]
  wire  rs1_addr_N0_0; // @[BackEnd.scala 398:47:@8730.4]
  wire  _T_1054; // @[BackEnd.scala 401:48:@8735.4]
  wire  _T_1055; // @[BackEnd.scala 401:66:@8736.4]
  wire  _T_1047; // @[BackEnd.scala 397:62:@8727.4]
  wire  exe_load_inst_0; // @[BackEnd.scala 397:44:@8728.4]
  wire  _T_1056; // @[BackEnd.scala 401:89:@8737.4]
  wire  rs2_addr_N0_0; // @[BackEnd.scala 399:47:@8732.4]
  wire  _T_1058; // @[BackEnd.scala 402:48:@8739.4]
  wire  _T_1059; // @[BackEnd.scala 402:66:@8740.4]
  wire  _T_1060; // @[BackEnd.scala 402:89:@8741.4]
  wire  _T_1061; // @[BackEnd.scala 401:110:@8742.4]
  wire  _T_1063; // @[BackEnd.scala 403:48:@8744.4]
  wire  _T_1064; // @[BackEnd.scala 403:66:@8745.4]
  wire  _T_1072; // @[BackEnd.scala 397:62:@8754.4]
  wire  exe_load_inst_1; // @[BackEnd.scala 397:44:@8755.4]
  wire  _T_1065; // @[BackEnd.scala 403:89:@8746.4]
  wire  _T_1066; // @[BackEnd.scala 402:110:@8747.4]
  wire  _T_1068; // @[BackEnd.scala 404:48:@8749.4]
  wire  _T_1069; // @[BackEnd.scala 404:66:@8750.4]
  wire  _T_1070; // @[BackEnd.scala 404:89:@8751.4]
  wire  rAW_0; // @[BackEnd.scala 403:110:@8752.4]
  wire [2:0] exe_wire_0_csr_cmd; // @[BackEnd.scala 213:31:@8251.4]
  wire  _T_1097; // @[BackEnd.scala 407:56:@8781.4]
  wire  _T_1098; // @[BackEnd.scala 407:33:@8782.4]
  wire [2:0] exe_wire_1_csr_cmd; // @[BackEnd.scala 213:31:@8290.4]
  wire  _T_1099; // @[BackEnd.scala 407:89:@8783.4]
  wire  stall_0_0; // @[BackEnd.scala 407:66:@8784.4]
  wire  _T_696; // @[BackEnd.scala 192:31:@8202.4]
  wire  _T_702; // @[BackEnd.scala 192:79:@8206.4]
  wire  ma_jump; // @[BackEnd.scala 344:29:@8602.4]
  wire  mem_en; // @[BackEnd.scala 326:25:@8490.4]
  wire  mem_fcn; // @[BackEnd.scala 327:25:@8491.4]
  wire  _T_907; // @[BackEnd.scala 342:44:@8596.4]
  wire  _T_908; // @[BackEnd.scala 342:33:@8597.4]
  wire [2:0] mem_typ; // @[BackEnd.scala 328:25:@8492.4]
  wire [1:0] _T_896; // @[BackEnd.scala 337:43:@8588.4]
  wire  _T_906; // @[Mux.scala 46:19:@8594.4]
  wire [31:0] mem_exe_out; // @[BackEnd.scala 322:25:@8486.4]
  wire  _T_899; // @[BackEnd.scala 338:23:@8589.4]
  wire  _T_904; // @[Mux.scala 46:19:@8592.4]
  wire [1:0] _T_901; // @[BackEnd.scala 339:23:@8590.4]
  wire  _T_903; // @[BackEnd.scala 339:29:@8591.4]
  wire  _T_905; // @[Mux.scala 46:16:@8593.4]
  wire  ls_addr_ma_valid; // @[Mux.scala 46:16:@8595.4]
  wire  ma_load; // @[BackEnd.scala 342:54:@8598.4]
  wire  _T_928; // @[BackEnd.scala 359:25:@8618.4]
  wire  _T_910; // @[BackEnd.scala 343:33:@8600.4]
  wire  ma_store; // @[BackEnd.scala 343:54:@8601.4]
  wire  _T_929; // @[BackEnd.scala 359:36:@8619.4]
  wire  ma_illegal; // @[BackEnd.scala 345:29:@8603.4]
  wire  _T_930; // @[BackEnd.scala 359:48:@8620.4]
  wire  xcpt_valid; // @[BackEnd.scala 359:62:@8621.4]
  wire  _T_703; // @[BackEnd.scala 192:104:@8207.4]
  wire  not_expect; // @[BackEnd.scala 266:53:@8371.4]
  wire  exe_wire_0_isBJ; // @[BackEnd.scala 210:41:@8245.4]
  wire  exe_wire_1_isBJ; // @[BackEnd.scala 210:41:@8284.4]
  wire  exe_wire_isBJ; // @[BackEnd.scala 245:54:@8321.4]
  wire  mispredict; // @[BackEnd.scala 267:28:@8372.4]
  wire  _T_711; // @[BackEnd.scala 195:47:@8216.8]
  wire  _T_712; // @[BackEnd.scala 195:44:@8217.8]
  wire  _GEN_38; // @[BackEnd.scala 194:60:@8215.6]
  wire  _GEN_39; // @[BackEnd.scala 192:119:@8208.4]
  wire  _T_1101; // @[BackEnd.scala 410:26:@8786.4]
  wire  rs1_addr_N0_1; // @[BackEnd.scala 398:47:@8757.4]
  wire  _T_1102; // @[BackEnd.scala 410:52:@8787.4]
  wire  _T_1103; // @[BackEnd.scala 410:70:@8788.4]
  wire  _T_1104; // @[BackEnd.scala 410:93:@8789.4]
  wire  _T_1105; // @[BackEnd.scala 411:26:@8790.4]
  wire  rs2_addr_N0_1; // @[BackEnd.scala 399:47:@8759.4]
  wire  _T_1106; // @[BackEnd.scala 411:52:@8791.4]
  wire  _T_1107; // @[BackEnd.scala 411:70:@8792.4]
  wire  _T_1108; // @[BackEnd.scala 411:93:@8793.4]
  wire  _T_1109; // @[BackEnd.scala 410:116:@8794.4]
  wire  _T_1110; // @[BackEnd.scala 412:25:@8795.4]
  wire  _T_1111; // @[BackEnd.scala 411:116:@8796.4]
  wire  _T_1079; // @[BackEnd.scala 401:48:@8762.4]
  wire  _T_1080; // @[BackEnd.scala 401:66:@8763.4]
  wire  _T_1081; // @[BackEnd.scala 401:89:@8764.4]
  wire  _T_1083; // @[BackEnd.scala 402:48:@8766.4]
  wire  _T_1084; // @[BackEnd.scala 402:66:@8767.4]
  wire  _T_1085; // @[BackEnd.scala 402:89:@8768.4]
  wire  _T_1086; // @[BackEnd.scala 401:110:@8769.4]
  wire  _T_1088; // @[BackEnd.scala 403:48:@8771.4]
  wire  _T_1089; // @[BackEnd.scala 403:66:@8772.4]
  wire  _T_1090; // @[BackEnd.scala 403:89:@8773.4]
  wire  _T_1091; // @[BackEnd.scala 402:110:@8774.4]
  wire  _T_1093; // @[BackEnd.scala 404:48:@8776.4]
  wire  _T_1094; // @[BackEnd.scala 404:66:@8777.4]
  wire  _T_1095; // @[BackEnd.scala 404:89:@8778.4]
  wire  rAW_1; // @[BackEnd.scala 403:110:@8779.4]
  wire  _T_1112; // @[BackEnd.scala 412:35:@8797.4]
  wire  stall_1_0; // @[BackEnd.scala 412:45:@8798.4]
  wire  _T_715; // @[BackEnd.scala 198:30:@8221.4]
  wire  _T_718; // @[BackEnd.scala 198:54:@8223.4]
  wire  _T_719; // @[BackEnd.scala 198:79:@8224.4]
  wire  exe_cancel; // @[BackEnd.scala 268:28:@8374.4]
  wire  _T_720; // @[BackEnd.scala 198:93:@8225.4]
  wire  _T_729; // @[BackEnd.scala 201:44:@8235.8]
  wire  _GEN_40; // @[BackEnd.scala 200:60:@8233.6]
  wire  _GEN_41; // @[BackEnd.scala 198:108:@8226.4]
  wire [31:0] target_brjmp; // @[BackEnd.scala 241:19:@8317.4]
  wire [31:0] target_jpreg; // @[BackEnd.scala 241:19:@8317.4]
  wire [31:0] target_conti; // @[BackEnd.scala 241:19:@8317.4]
  wire [1:0] pc_sel; // @[BackEnd.scala 242:19:@8318.4]
  wire  exe_wire_branch; // @[BackEnd.scala 246:39:@8322.4]
  wire  exe_wire_pop; // @[BackEnd.scala 247:39:@8323.4]
  wire  exe_wire_push; // @[BackEnd.scala 248:39:@8324.4]
  reg  _T_766; // @[BackEnd.scala 66:27:@8326.4]
  reg [31:0] _RAND_73;
  wire  _GEN_66; // @[BackEnd.scala 68:20:@8331.6]
  wire  _GEN_67; // @[BackEnd.scala 67:20:@8327.4]
  reg  _T_774; // @[BackEnd.scala 66:27:@8337.4]
  reg [31:0] _RAND_74;
  wire  _GEN_68; // @[BackEnd.scala 68:20:@8342.6]
  wire  _GEN_69; // @[BackEnd.scala 67:20:@8338.4]
  reg  _T_782; // @[BackEnd.scala 66:27:@8349.4]
  reg [31:0] _RAND_75;
  wire  _GEN_70; // @[BackEnd.scala 68:20:@8354.6]
  wire  _GEN_71; // @[BackEnd.scala 67:20:@8350.4]
  wire  _T_786; // @[BackEnd.scala 255:45:@8359.4]
  wire  _T_787; // @[BackEnd.scala 255:68:@8360.4]
  wire [31:0] _T_791; // @[BackEnd.scala 258:10:@8365.4]
  wire [1:0] _T_796; // @[BackEnd.scala 264:10:@8368.4]
  wire [31:0] _T_808; // @[Bitwise.scala 72:12:@8381.6]
  wire [31:0] _T_809; // @[BackEnd.scala 273:47:@8382.6]
  wire [31:0] _T_814; // @[Bitwise.scala 72:12:@8385.6]
  wire [31:0] _T_815; // @[BackEnd.scala 274:47:@8386.6]
  wire [31:0] _T_816; // @[BackEnd.scala 273:63:@8387.6]
  wire [31:0] _GEN_72; // @[BackEnd.scala 271:31:@8378.4]
  wire  _T_819; // @[BackEnd.scala 277:57:@8391.4]
  wire  _T_820; // @[BackEnd.scala 277:54:@8392.4]
  wire  _T_821; // @[BackEnd.scala 277:78:@8393.4]
  wire  _GEN_73; // @[BackEnd.scala 279:37:@8399.6]
  wire  _GEN_74; // @[BackEnd.scala 277:93:@8394.4]
  wire  _T_827; // @[BackEnd.scala 283:30:@8403.4]
  wire  _T_828; // @[BackEnd.scala 283:55:@8404.4]
  wire  _T_833; // @[BackEnd.scala 286:37:@8411.8]
  wire  _T_834; // @[BackEnd.scala 286:34:@8412.8]
  wire  _GEN_75; // @[BackEnd.scala 285:37:@8410.6]
  wire  _GEN_76; // @[BackEnd.scala 283:70:@8405.4]
  wire  _T_837; // @[BackEnd.scala 289:69:@8416.4]
  wire [31:0] mem_inst; // @[BackEnd.scala 321:25:@8485.4]
  wire  _T_911; // @[BackEnd.scala 346:27:@8604.4]
  wire  _T_912; // @[BackEnd.scala 346:39:@8605.4]
  wire [2:0] _T_919; // @[Mux.scala 61:16:@8608.4]
  wire [2:0] _T_920; // @[Mux.scala 61:16:@8609.4]
  wire [2:0] _T_921; // @[Mux.scala 61:16:@8610.4]
  wire [2:0] _T_922; // @[Mux.scala 61:16:@8611.4]
  wire [31:0] _T_924; // @[Mux.scala 61:16:@8613.4]
  wire [31:0] _T_925; // @[Mux.scala 61:16:@8614.4]
  wire [31:0] _T_926; // @[Mux.scala 61:16:@8615.4]
  wire  _T_932; // @[BackEnd.scala 362:44:@8624.4]
  wire  _T_933; // @[BackEnd.scala 362:29:@8625.4]
  wire  _GEN_77; // @[BackEnd.scala 362:60:@8626.4]
  wire  _T_935; // @[BackEnd.scala 366:29:@8632.4]
  wire  _GEN_78; // @[BackEnd.scala 366:44:@8633.4]
  wire [1:0] _T_952; // @[BackEnd.scala 385:25:@8654.4]
  wire  retire_0; // @[BackEnd.scala 385:32:@8655.4]
  wire [1:0] _T_955; // @[BackEnd.scala 386:32:@8658.4]
  wire  retire_1; // @[BackEnd.scala 386:32:@8659.4]
  reg  _T_1133; // @[BackEnd.scala 66:27:@8816.4]
  reg [31:0] _RAND_76;
  wire  _GEN_79; // @[BackEnd.scala 68:20:@8821.6]
  wire  _GEN_80; // @[BackEnd.scala 67:20:@8817.4]
  wire  _T_1138; // @[BackEnd.scala 421:26:@8828.4]
  wire  _T_1141; // @[BackEnd.scala 421:47:@8830.4]
  wire  _T_1146; // @[BackEnd.scala 422:26:@8834.4]
  wire  _T_1149; // @[BackEnd.scala 422:47:@8836.4]
  wire  _T_1152; // @[BackEnd.scala 422:71:@8838.4]
  wire  _T_1153; // @[BackEnd.scala 423:35:@8839.4]
  wire  _T_1155; // @[BackEnd.scala 423:5:@8840.4]
  wire [7:0] _T_1159; // @[BackEnd.scala 432:12:@8843.4]
  wire [7:0] _T_1167; // @[BackEnd.scala 434:12:@8845.4]
  wire  _T_1170; // @[BackEnd.scala 435:32:@8846.4]
  wire  _T_1173; // @[BackEnd.scala 436:32:@8847.4]
  wire  _T_1176; // @[BackEnd.scala 437:32:@8848.4]
  wire  _T_1179; // @[BackEnd.scala 438:32:@8849.4]
  wire [7:0] _T_1182; // @[BackEnd.scala 438:12:@8850.4]
  wire [7:0] _T_1183; // @[BackEnd.scala 437:12:@8851.4]
  wire [7:0] _T_1184; // @[BackEnd.scala 436:12:@8852.4]
  wire [7:0] _T_1185; // @[BackEnd.scala 435:12:@8853.4]
  wire [7:0] _T_1189; // @[BackEnd.scala 439:12:@8854.4]
  wire  _T_1192; // @[BackEnd.scala 440:13:@8855.4]
  wire  _T_1193; // @[BackEnd.scala 440:27:@8856.4]
  wire  _T_1199; // @[BackEnd.scala 440:72:@8860.4]
  wire [31:0] _T_1205; // @[BackEnd.scala 440:12:@8864.4]
  wire  _T_1208; // @[BackEnd.scala 427:11:@8866.4]
  wire [7:0] _T_1211; // @[BackEnd.scala 432:12:@8870.4]
  wire [7:0] _T_1215; // @[BackEnd.scala 433:12:@8871.4]
  wire [7:0] _T_1219; // @[BackEnd.scala 434:12:@8872.4]
  wire  _T_1222; // @[BackEnd.scala 435:32:@8873.4]
  wire  _T_1225; // @[BackEnd.scala 436:32:@8874.4]
  wire  _T_1228; // @[BackEnd.scala 437:32:@8875.4]
  wire  _T_1231; // @[BackEnd.scala 438:32:@8876.4]
  wire [7:0] _T_1234; // @[BackEnd.scala 438:12:@8877.4]
  wire [7:0] _T_1235; // @[BackEnd.scala 437:12:@8878.4]
  wire [7:0] _T_1236; // @[BackEnd.scala 436:12:@8879.4]
  wire [7:0] _T_1237; // @[BackEnd.scala 435:12:@8880.4]
  wire  _T_1244; // @[BackEnd.scala 440:13:@8882.4]
  wire  _T_1245; // @[BackEnd.scala 440:27:@8883.4]
  wire  _T_1250; // @[BackEnd.scala 440:41:@8886.4]
  wire  _T_1251; // @[BackEnd.scala 440:72:@8887.4]
  wire  _T_1256; // @[BackEnd.scala 441:29:@8890.4]
  wire [31:0] _T_1257; // @[BackEnd.scala 440:12:@8891.4]
  wire  _T_1267; // @[BackEnd.scala 462:22:@8912.6]
  wire [31:0] _T_1268; // @[BackEnd.scala 463:12:@8913.6]
  CSRFile csr ( // @[BackEnd.scala 80:19:@7927.4]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_status_prv(csr_io_status_prv),
    .io_status_unimp5(csr_io_status_unimp5),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_unimp4(csr_io_status_unimp4),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_unimp3(csr_io_status_unimp3),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_unimp2(csr_io_status_unimp2),
    .io_status_mie(csr_io_status_mie),
    .io_status_unimp1(csr_io_status_unimp1),
    .io_xcpt(csr_io_xcpt),
    .io_cause(csr_io_cause),
    .io_tval(csr_io_tval),
    .io_evec(csr_io_evec),
    .io_illegal(csr_io_illegal),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    .io_time(csr_io_time)
  );
  Regfile regfile ( // @[BackEnd.scala 81:23:@7930.4]
    .clock(regfile_clock),
    .io_rs1_addr_0(regfile_io_rs1_addr_0),
    .io_rs1_addr_1(regfile_io_rs1_addr_1),
    .io_rs1_data_0(regfile_io_rs1_data_0),
    .io_rs1_data_1(regfile_io_rs1_data_1),
    .io_rs2_addr_0(regfile_io_rs2_addr_0),
    .io_rs2_addr_1(regfile_io_rs2_addr_1),
    .io_rs2_data_0(regfile_io_rs2_data_0),
    .io_rs2_data_1(regfile_io_rs2_data_1),
    .io_waddr_0(regfile_io_waddr_0),
    .io_waddr_1(regfile_io_waddr_1),
    .io_wdata_0(regfile_io_wdata_0),
    .io_wdata_1(regfile_io_wdata_1),
    .io_wen_0(regfile_io_wen_0),
    .io_wen_1(regfile_io_wen_1)
  );
  ALU ALU ( // @[BackEnd.scala 82:33:@7933.4]
    .io_op1(ALU_io_op1),
    .io_op2(ALU_io_op2),
    .io_pc(ALU_io_pc),
    .io_ctrl_fun(ALU_io_ctrl_fun),
    .io_ctrl_br_type(ALU_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_io_ctrl_pc_sel),
    .io_rs2_data(ALU_io_rs2_data),
    .io_result(ALU_io_result),
    .io_target_brjmp(ALU_io_target_brjmp),
    .io_target_jpreg(ALU_io_target_jpreg),
    .io_target_conti(ALU_io_target_conti)
  );
  ALU ALU_1 ( // @[BackEnd.scala 82:33:@7936.4]
    .io_op1(ALU_1_io_op1),
    .io_op2(ALU_1_io_op2),
    .io_pc(ALU_1_io_pc),
    .io_ctrl_fun(ALU_1_io_ctrl_fun),
    .io_ctrl_br_type(ALU_1_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_1_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_1_io_ctrl_pc_sel),
    .io_rs2_data(ALU_1_io_rs2_data),
    .io_result(ALU_1_io_result),
    .io_target_brjmp(ALU_1_io_target_brjmp),
    .io_target_jpreg(ALU_1_io_target_jpreg),
    .io_target_conti(ALU_1_io_target_conti)
  );
  InstDecoder InstDecoder ( // @[BackEnd.scala 83:33:@7939.4]
    .io_inst(InstDecoder_io_inst),
    .io_cinfo_br_type(InstDecoder_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_io_cinfo_illegal),
    .io_cinfo_fencei(InstDecoder_io_cinfo_fencei),
    .io_cinfo_branch(InstDecoder_io_cinfo_branch),
    .io_cinfo_push(InstDecoder_io_cinfo_push),
    .io_cinfo_pop(InstDecoder_io_cinfo_pop),
    .io_cinfo_isBJ(InstDecoder_io_cinfo_isBJ),
    .io_cinfo_rs1_addr(InstDecoder_io_cinfo_rs1_addr),
    .io_cinfo_rs2_addr(InstDecoder_io_cinfo_rs2_addr),
    .io_cinfo_wbaddr(InstDecoder_io_cinfo_wbaddr),
    .io_dinfo_imm_i(InstDecoder_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_io_dinfo_imm_z)
  );
  InstDecoder InstDecoder_1 ( // @[BackEnd.scala 83:33:@7942.4]
    .io_inst(InstDecoder_1_io_inst),
    .io_cinfo_br_type(InstDecoder_1_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_1_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_1_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_1_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_1_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_1_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_1_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_1_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_1_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_1_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_1_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_1_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_1_io_cinfo_illegal),
    .io_cinfo_fencei(InstDecoder_1_io_cinfo_fencei),
    .io_cinfo_branch(InstDecoder_1_io_cinfo_branch),
    .io_cinfo_push(InstDecoder_1_io_cinfo_push),
    .io_cinfo_pop(InstDecoder_1_io_cinfo_pop),
    .io_cinfo_isBJ(InstDecoder_1_io_cinfo_isBJ),
    .io_cinfo_rs1_addr(InstDecoder_1_io_cinfo_rs1_addr),
    .io_cinfo_rs2_addr(InstDecoder_1_io_cinfo_rs2_addr),
    .io_cinfo_wbaddr(InstDecoder_1_io_cinfo_wbaddr),
    .io_dinfo_imm_i(InstDecoder_1_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_1_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_1_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_1_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_1_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_1_io_dinfo_imm_z)
  );
  assign dec_wire_0_fencei = io_front_inst_0_valid & InstDecoder_io_cinfo_fencei; // @[BackEnd.scala 120:51:@7992.4]
  assign dec_wire_1_fencei = io_front_inst_1_valid & InstDecoder_1_io_cinfo_fencei; // @[BackEnd.scala 120:51:@8093.4]
  assign _T_473 = dec_wire_0_fencei | dec_wire_1_fencei; // @[BackEnd.scala 100:54:@7968.4]
  assign exe_wire_0_fencei = exe_valid_0 & exe_0_fencei; // @[BackEnd.scala 211:41:@8247.4]
  assign exe_wire_1_fencei = exe_valid_1 & exe_1_fencei; // @[BackEnd.scala 211:41:@8286.4]
  assign _T_474 = exe_wire_0_fencei | exe_wire_1_fencei; // @[BackEnd.scala 100:93:@7969.4]
  assign dec_wire_0_rs1_oen = io_front_inst_0_valid & InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 116:51:@7982.4]
  assign dec_wire_0_rs2_oen = io_front_inst_0_valid & InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 117:51:@7984.4]
  assign _T_541 = io_front_inst_0_valid & InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 118:51:@7986.4]
  assign _T_543 = InstDecoder_io_cinfo_wbaddr != 5'h0; // @[BackEnd.scala 118:97:@7987.4]
  assign dec_wire_0_rf_wen = _T_541 & _T_543; // @[BackEnd.scala 118:74:@7988.4]
  assign dec_wire_0_isBJ = io_front_inst_0_valid & InstDecoder_io_cinfo_isBJ; // @[BackEnd.scala 119:51:@7990.4]
  assign dec_wire_0_csr_cmd = io_front_inst_0_valid ? InstDecoder_io_cinfo_csr_cmd : 3'h0; // @[BackEnd.scala 121:31:@7994.4]
  assign _T_548 = exe_1_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 129:23:@8000.4]
  assign _T_749 = exe_valid_1 & exe_1_rf_wen; // @[BackEnd.scala 208:41:@8278.4]
  assign _T_751 = exe_1_wbaddr != 5'h0; // @[BackEnd.scala 208:75:@8279.4]
  assign exe_wire_1_rf_wen = _T_749 & _T_751; // @[BackEnd.scala 208:58:@8280.4]
  assign _T_549 = _T_548 & exe_wire_1_rf_wen; // @[BackEnd.scala 129:50:@8001.4]
  assign _T_550 = exe_0_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 130:23:@8002.4]
  assign _T_737 = exe_valid_0 & exe_0_rf_wen; // @[BackEnd.scala 208:41:@8239.4]
  assign _T_739 = exe_0_wbaddr != 5'h0; // @[BackEnd.scala 208:75:@8240.4]
  assign exe_wire_0_rf_wen = _T_737 & _T_739; // @[BackEnd.scala 208:58:@8241.4]
  assign _T_551 = _T_550 & exe_wire_0_rf_wen; // @[BackEnd.scala 130:50:@8003.4]
  assign _T_552 = mem_1_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 131:23:@8004.4]
  assign _T_876 = mem_valid_1 & mem_1_rf_wen; // @[BackEnd.scala 300:41:@8457.4]
  assign _T_878 = mem_1_wbaddr != 5'h0; // @[BackEnd.scala 300:75:@8458.4]
  assign mem_wire_1_rf_wen = _T_876 & _T_878; // @[BackEnd.scala 300:58:@8459.4]
  assign _T_553 = _T_552 & mem_wire_1_rf_wen; // @[BackEnd.scala 131:50:@8005.4]
  assign _T_554 = mem_0_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 132:23:@8006.4]
  assign _T_857 = mem_valid_0 & mem_0_rf_wen; // @[BackEnd.scala 300:41:@8429.4]
  assign _T_859 = mem_0_wbaddr != 5'h0; // @[BackEnd.scala 300:75:@8430.4]
  assign mem_wire_0_rf_wen = _T_857 & _T_859; // @[BackEnd.scala 300:58:@8431.4]
  assign _T_555 = _T_554 & mem_wire_0_rf_wen; // @[BackEnd.scala 132:50:@8007.4]
  assign _T_556 = wb_1_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 133:23:@8008.4]
  assign _T_941 = wb_valid_1 & wb_1_rf_wen; // @[BackEnd.scala 373:40:@8646.4]
  assign _T_943 = wb_1_wbaddr != 5'h0; // @[BackEnd.scala 373:72:@8647.4]
  assign wb_wire_1_rf_wen = _T_941 & _T_943; // @[BackEnd.scala 373:56:@8648.4]
  assign _T_557 = _T_556 & wb_wire_1_rf_wen; // @[BackEnd.scala 133:50:@8009.4]
  assign _T_558 = wb_0_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 134:23:@8010.4]
  assign _T_937 = wb_valid_0 & wb_0_rf_wen; // @[BackEnd.scala 373:40:@8639.4]
  assign _T_939 = wb_0_wbaddr != 5'h0; // @[BackEnd.scala 373:72:@8640.4]
  assign wb_wire_0_rf_wen = _T_937 & _T_939; // @[BackEnd.scala 373:56:@8641.4]
  assign _T_559 = _T_558 & wb_wire_0_rf_wen; // @[BackEnd.scala 134:50:@8011.4]
  assign rf_rs1_data_0 = regfile_io_rs1_data_0; // @[BackEnd.scala 112:25:@7979.4 BackEnd.scala 125:20:@7998.4]
  assign _T_560 = _T_559 ? wb_wbdata_0 : rf_rs1_data_0; // @[Mux.scala 61:16:@8012.4]
  assign _T_561 = _T_557 ? wb_wbdata_1 : _T_560; // @[Mux.scala 61:16:@8013.4]
  assign _T_872 = mem_0_wb_sel == 2'h1; // @[BackEnd.scala 312:22:@8448.4]
  assign _T_873 = mem_0_wb_sel == 2'h3; // @[BackEnd.scala 313:22:@8449.4]
  assign _T_874 = _T_873 ? csr_io_rw_rdata : mem_reg_wbdata_0; // @[Mux.scala 61:16:@8450.4]
  assign mem_wbdata_0 = _T_872 ? io_mem_resp_bits_data : _T_874; // @[Mux.scala 61:16:@8451.4]
  assign _T_562 = _T_555 ? mem_wbdata_0 : _T_561; // @[Mux.scala 61:16:@8014.4]
  assign _T_891 = mem_1_wb_sel == 2'h1; // @[BackEnd.scala 312:22:@8476.4]
  assign _T_892 = mem_1_wb_sel == 2'h3; // @[BackEnd.scala 313:22:@8477.4]
  assign _T_893 = _T_892 ? csr_io_rw_rdata : mem_reg_wbdata_1; // @[Mux.scala 61:16:@8478.4]
  assign mem_wbdata_1 = _T_891 ? io_mem_resp_bits_data : _T_893; // @[Mux.scala 61:16:@8479.4]
  assign _T_563 = _T_553 ? mem_wbdata_1 : _T_562; // @[Mux.scala 61:16:@8015.4]
  assign exe_wbdata_0 = ALU_io_result; // @[BackEnd.scala 102:24:@7972.4 BackEnd.scala 224:19:@8262.4]
  assign _T_564 = _T_551 ? exe_wbdata_0 : _T_563; // @[Mux.scala 61:16:@8016.4]
  assign exe_wbdata_1 = ALU_1_io_result; // @[BackEnd.scala 102:24:@7972.4 BackEnd.scala 224:19:@8301.4]
  assign dec_rs1_data_0 = _T_549 ? exe_wbdata_1 : _T_564; // @[Mux.scala 61:16:@8017.4]
  assign _T_566 = exe_1_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 138:23:@8019.4]
  assign _T_567 = _T_566 & exe_wire_1_rf_wen; // @[BackEnd.scala 138:50:@8020.4]
  assign _T_568 = exe_0_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 139:23:@8021.4]
  assign _T_569 = _T_568 & exe_wire_0_rf_wen; // @[BackEnd.scala 139:50:@8022.4]
  assign _T_570 = mem_1_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 140:23:@8023.4]
  assign _T_571 = _T_570 & mem_wire_1_rf_wen; // @[BackEnd.scala 140:50:@8024.4]
  assign _T_572 = mem_0_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 141:23:@8025.4]
  assign _T_573 = _T_572 & mem_wire_0_rf_wen; // @[BackEnd.scala 141:50:@8026.4]
  assign _T_574 = wb_1_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 142:23:@8027.4]
  assign _T_575 = _T_574 & wb_wire_1_rf_wen; // @[BackEnd.scala 142:50:@8028.4]
  assign _T_576 = wb_0_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 143:23:@8029.4]
  assign _T_577 = _T_576 & wb_wire_0_rf_wen; // @[BackEnd.scala 143:50:@8030.4]
  assign rf_rs2_data_0 = regfile_io_rs2_data_0; // @[BackEnd.scala 113:25:@7980.4 BackEnd.scala 126:20:@7999.4]
  assign _T_578 = _T_577 ? wb_wbdata_0 : rf_rs2_data_0; // @[Mux.scala 61:16:@8031.4]
  assign _T_579 = _T_575 ? wb_wbdata_1 : _T_578; // @[Mux.scala 61:16:@8032.4]
  assign _T_580 = _T_573 ? mem_wbdata_0 : _T_579; // @[Mux.scala 61:16:@8033.4]
  assign _T_581 = _T_571 ? mem_wbdata_1 : _T_580; // @[Mux.scala 61:16:@8034.4]
  assign _T_582 = _T_569 ? exe_wbdata_0 : _T_581; // @[Mux.scala 61:16:@8035.4]
  assign dec_rs2_data_0 = _T_567 ? exe_wbdata_1 : _T_582; // @[Mux.scala 61:16:@8036.4]
  assign _T_584 = InstDecoder_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 147:29:@8038.4]
  assign _T_585 = InstDecoder_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 148:29:@8039.4]
  assign _T_586 = _T_585 ? io_front_pc_0 : dec_rs1_data_0; // @[Mux.scala 61:16:@8040.4]
  assign dec_op1_data_0 = _T_584 ? InstDecoder_io_dinfo_imm_z : _T_586; // @[Mux.scala 61:16:@8041.4]
  assign _T_588 = InstDecoder_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 151:29:@8043.4]
  assign _T_589 = InstDecoder_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 152:29:@8044.4]
  assign _T_590 = InstDecoder_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 153:29:@8045.4]
  assign _T_591 = InstDecoder_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 154:29:@8046.4]
  assign _T_592 = InstDecoder_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 155:29:@8047.4]
  assign _T_593 = _T_592 ? InstDecoder_io_dinfo_imm_uj : dec_rs2_data_0; // @[Mux.scala 61:16:@8048.4]
  assign _T_594 = _T_591 ? InstDecoder_io_dinfo_imm_u : _T_593; // @[Mux.scala 61:16:@8049.4]
  assign _T_595 = _T_590 ? InstDecoder_io_dinfo_imm_sb : _T_594; // @[Mux.scala 61:16:@8050.4]
  assign _T_596 = _T_589 ? InstDecoder_io_dinfo_imm_s : _T_595; // @[Mux.scala 61:16:@8051.4]
  assign dec_op2_data_0 = _T_588 ? InstDecoder_io_dinfo_imm_i : _T_596; // @[Mux.scala 61:16:@8052.4]
  assign exe_wire_0_mem_en = exe_valid_0 & exe_0_mem_en; // @[BackEnd.scala 209:41:@8243.4]
  assign exe_wire_1_mem_en = exe_valid_1 & exe_1_mem_en; // @[BackEnd.scala 209:41:@8282.4]
  assign stall_1_1 = exe_wire_0_mem_en & exe_wire_1_mem_en; // @[BackEnd.scala 415:80:@8801.4]
  assign _T_599 = stall_1_1 == 1'h0; // @[BackEnd.scala 157:11:@8054.4]
  assign mem_wire_1_csr_cmd = mem_valid_1 ? mem_1_csr_cmd : 3'h0; // @[BackEnd.scala 302:31:@8463.4]
  assign _T_887 = mem_wire_1_csr_cmd != 3'h0; // @[BackEnd.scala 306:39:@8471.4]
  assign mem_wire_1_mem_en = mem_valid_1 & mem_1_mem_en; // @[BackEnd.scala 301:41:@8461.4]
  assign _T_888 = _T_887 | mem_wire_1_mem_en; // @[BackEnd.scala 306:49:@8472.4]
  assign mem_wire_1_illegal = mem_valid_1 & mem_1_illegal; // @[BackEnd.scala 303:41:@8465.4]
  assign _T_889 = _T_888 | mem_wire_1_illegal; // @[BackEnd.scala 307:39:@8473.4]
  assign _T_883 = mem_reg_jpnpc[1:0]; // @[BackEnd.scala 304:54:@8467.4]
  assign _T_885 = _T_883 != 2'h0; // @[BackEnd.scala 304:60:@8468.4]
  assign mem_wire_jump_1 = mem_valid_1 & _T_885; // @[BackEnd.scala 304:38:@8469.4]
  assign mem_sel_1 = _T_889 | mem_wire_jump_1; // @[BackEnd.scala 308:39:@8474.4]
  assign mem_wire_0_csr_cmd = mem_valid_0 ? mem_0_csr_cmd : 3'h0; // @[BackEnd.scala 302:31:@8435.4]
  assign _T_868 = mem_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 306:39:@8443.4]
  assign mem_wire_0_mem_en = mem_valid_0 & mem_0_mem_en; // @[BackEnd.scala 301:41:@8433.4]
  assign _T_869 = _T_868 | mem_wire_0_mem_en; // @[BackEnd.scala 306:49:@8444.4]
  assign mem_wire_0_illegal = mem_valid_0 & mem_0_illegal; // @[BackEnd.scala 303:41:@8437.4]
  assign _T_870 = _T_869 | mem_wire_0_illegal; // @[BackEnd.scala 307:39:@8445.4]
  assign mem_wire_jump_0 = mem_valid_0 & _T_885; // @[BackEnd.scala 304:38:@8441.4]
  assign mem_sel_0 = _T_870 | mem_wire_jump_0; // @[BackEnd.scala 308:39:@8446.4]
  assign _T_1120 = {mem_sel_1,mem_sel_0}; // @[BackEnd.scala 417:34:@8807.4]
  assign _T_1121 = ~ _T_1120; // @[BackEnd.scala 417:41:@8808.4]
  assign _T_1123 = _T_1121 == 2'h0; // @[BackEnd.scala 417:41:@8809.4]
  assign _T_1125 = io_mem_resp_valid == 1'h0; // @[BackEnd.scala 417:72:@8810.4]
  assign _T_1126 = mem_wire_1_mem_en & _T_1125; // @[BackEnd.scala 417:69:@8811.4]
  assign _T_1127 = _T_1123 | _T_1126; // @[BackEnd.scala 417:46:@8812.4]
  assign stall_0_2 = mem_wire_0_mem_en & _T_1125; // @[BackEnd.scala 416:45:@8805.4]
  assign stall_1_2 = _T_1127 | stall_0_2; // @[BackEnd.scala 417:92:@8813.4]
  assign _T_601 = stall_1_2 == 1'h0; // @[BackEnd.scala 157:35:@8055.4]
  assign _T_602 = _T_599 & _T_601; // @[BackEnd.scala 157:32:@8056.4]
  assign _T_603 = InstDecoder_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 161:52:@8060.6]
  assign _T_604 = InstDecoder_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 161:86:@8061.6]
  assign _T_605 = _T_603 | _T_604; // @[BackEnd.scala 161:62:@8062.6]
  assign _T_607 = InstDecoder_io_cinfo_rs1_addr == 5'h0; // @[BackEnd.scala 162:53:@8063.6]
  assign _T_608 = _T_605 & _T_607; // @[BackEnd.scala 161:97:@8064.6]
  assign _T_609 = _T_608 ? 3'h5 : InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 161:29:@8065.6]
  assign dec_wire_1_rs1_oen = io_front_inst_1_valid & InstDecoder_1_io_cinfo_rs1_oen; // @[BackEnd.scala 116:51:@8083.4]
  assign dec_wire_1_rs2_oen = io_front_inst_1_valid & InstDecoder_1_io_cinfo_rs2_oen; // @[BackEnd.scala 117:51:@8085.4]
  assign dec_wire_1_isBJ = io_front_inst_1_valid & InstDecoder_1_io_cinfo_isBJ; // @[BackEnd.scala 119:51:@8091.4]
  assign _T_619 = exe_1_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 129:23:@8101.4]
  assign _T_620 = _T_619 & exe_wire_1_rf_wen; // @[BackEnd.scala 129:50:@8102.4]
  assign _T_621 = exe_0_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 130:23:@8103.4]
  assign _T_622 = _T_621 & exe_wire_0_rf_wen; // @[BackEnd.scala 130:50:@8104.4]
  assign _T_623 = mem_1_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 131:23:@8105.4]
  assign _T_624 = _T_623 & mem_wire_1_rf_wen; // @[BackEnd.scala 131:50:@8106.4]
  assign _T_625 = mem_0_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 132:23:@8107.4]
  assign _T_626 = _T_625 & mem_wire_0_rf_wen; // @[BackEnd.scala 132:50:@8108.4]
  assign _T_627 = wb_1_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 133:23:@8109.4]
  assign _T_628 = _T_627 & wb_wire_1_rf_wen; // @[BackEnd.scala 133:50:@8110.4]
  assign _T_629 = wb_0_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 134:23:@8111.4]
  assign _T_630 = _T_629 & wb_wire_0_rf_wen; // @[BackEnd.scala 134:50:@8112.4]
  assign rf_rs1_data_1 = regfile_io_rs1_data_1; // @[BackEnd.scala 112:25:@7979.4 BackEnd.scala 125:20:@8099.4]
  assign _T_631 = _T_630 ? wb_wbdata_0 : rf_rs1_data_1; // @[Mux.scala 61:16:@8113.4]
  assign _T_632 = _T_628 ? wb_wbdata_1 : _T_631; // @[Mux.scala 61:16:@8114.4]
  assign _T_633 = _T_626 ? mem_wbdata_0 : _T_632; // @[Mux.scala 61:16:@8115.4]
  assign _T_634 = _T_624 ? mem_wbdata_1 : _T_633; // @[Mux.scala 61:16:@8116.4]
  assign _T_635 = _T_622 ? exe_wbdata_0 : _T_634; // @[Mux.scala 61:16:@8117.4]
  assign dec_rs1_data_1 = _T_620 ? exe_wbdata_1 : _T_635; // @[Mux.scala 61:16:@8118.4]
  assign _T_637 = exe_1_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 138:23:@8120.4]
  assign _T_638 = _T_637 & exe_wire_1_rf_wen; // @[BackEnd.scala 138:50:@8121.4]
  assign _T_639 = exe_0_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 139:23:@8122.4]
  assign _T_640 = _T_639 & exe_wire_0_rf_wen; // @[BackEnd.scala 139:50:@8123.4]
  assign _T_641 = mem_1_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 140:23:@8124.4]
  assign _T_642 = _T_641 & mem_wire_1_rf_wen; // @[BackEnd.scala 140:50:@8125.4]
  assign _T_643 = mem_0_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 141:23:@8126.4]
  assign _T_644 = _T_643 & mem_wire_0_rf_wen; // @[BackEnd.scala 141:50:@8127.4]
  assign _T_645 = wb_1_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 142:23:@8128.4]
  assign _T_646 = _T_645 & wb_wire_1_rf_wen; // @[BackEnd.scala 142:50:@8129.4]
  assign _T_647 = wb_0_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 143:23:@8130.4]
  assign _T_648 = _T_647 & wb_wire_0_rf_wen; // @[BackEnd.scala 143:50:@8131.4]
  assign rf_rs2_data_1 = regfile_io_rs2_data_1; // @[BackEnd.scala 113:25:@7980.4 BackEnd.scala 126:20:@8100.4]
  assign _T_649 = _T_648 ? wb_wbdata_0 : rf_rs2_data_1; // @[Mux.scala 61:16:@8132.4]
  assign _T_650 = _T_646 ? wb_wbdata_1 : _T_649; // @[Mux.scala 61:16:@8133.4]
  assign _T_651 = _T_644 ? mem_wbdata_0 : _T_650; // @[Mux.scala 61:16:@8134.4]
  assign _T_652 = _T_642 ? mem_wbdata_1 : _T_651; // @[Mux.scala 61:16:@8135.4]
  assign _T_653 = _T_640 ? exe_wbdata_0 : _T_652; // @[Mux.scala 61:16:@8136.4]
  assign dec_rs2_data_1 = _T_638 ? exe_wbdata_1 : _T_653; // @[Mux.scala 61:16:@8137.4]
  assign _T_655 = InstDecoder_1_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 147:29:@8139.4]
  assign _T_656 = InstDecoder_1_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 148:29:@8140.4]
  assign _T_657 = _T_656 ? io_front_pc_1 : dec_rs1_data_1; // @[Mux.scala 61:16:@8141.4]
  assign dec_op1_data_1 = _T_655 ? InstDecoder_1_io_dinfo_imm_z : _T_657; // @[Mux.scala 61:16:@8142.4]
  assign _T_659 = InstDecoder_1_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 151:29:@8144.4]
  assign _T_660 = InstDecoder_1_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 152:29:@8145.4]
  assign _T_661 = InstDecoder_1_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 153:29:@8146.4]
  assign _T_662 = InstDecoder_1_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 154:29:@8147.4]
  assign _T_663 = InstDecoder_1_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 155:29:@8148.4]
  assign _T_664 = _T_663 ? InstDecoder_1_io_dinfo_imm_uj : dec_rs2_data_1; // @[Mux.scala 61:16:@8149.4]
  assign _T_665 = _T_662 ? InstDecoder_1_io_dinfo_imm_u : _T_664; // @[Mux.scala 61:16:@8150.4]
  assign _T_666 = _T_661 ? InstDecoder_1_io_dinfo_imm_sb : _T_665; // @[Mux.scala 61:16:@8151.4]
  assign _T_667 = _T_660 ? InstDecoder_1_io_dinfo_imm_s : _T_666; // @[Mux.scala 61:16:@8152.4]
  assign dec_op2_data_1 = _T_659 ? InstDecoder_1_io_dinfo_imm_i : _T_667; // @[Mux.scala 61:16:@8153.4]
  assign _T_674 = InstDecoder_1_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 161:52:@8161.6]
  assign _T_675 = InstDecoder_1_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 161:86:@8162.6]
  assign _T_676 = _T_674 | _T_675; // @[BackEnd.scala 161:62:@8163.6]
  assign _T_678 = InstDecoder_1_io_cinfo_rs1_addr == 5'h0; // @[BackEnd.scala 162:53:@8164.6]
  assign _T_679 = _T_676 & _T_678; // @[BackEnd.scala 161:97:@8165.6]
  assign _T_680 = _T_679 ? 3'h5 : InstDecoder_1_io_cinfo_csr_cmd; // @[BackEnd.scala 161:29:@8166.6]
  assign _T_690 = dec_wire_0_isBJ ? io_front_pred_0 : io_front_pred_1; // @[BackEnd.scala 184:26:@8191.6]
  assign _T_691 = dec_wire_0_isBJ ? InstDecoder_io_cinfo_branch : InstDecoder_1_io_cinfo_branch; // @[BackEnd.scala 185:26:@8193.6]
  assign _T_692 = dec_wire_0_isBJ ? InstDecoder_io_cinfo_pop : InstDecoder_1_io_cinfo_pop; // @[BackEnd.scala 186:26:@8195.6]
  assign _T_693 = dec_wire_0_isBJ ? InstDecoder_io_cinfo_push : InstDecoder_1_io_cinfo_push; // @[BackEnd.scala 187:26:@8197.6]
  assign rs1_addr_N0_0 = InstDecoder_io_cinfo_rs1_addr != 5'h0; // @[BackEnd.scala 398:47:@8730.4]
  assign _T_1054 = _T_550 & rs1_addr_N0_0; // @[BackEnd.scala 401:48:@8735.4]
  assign _T_1055 = _T_1054 & dec_wire_0_rs1_oen; // @[BackEnd.scala 401:66:@8736.4]
  assign _T_1047 = exe_0_mem_fcn == 1'h0; // @[BackEnd.scala 397:62:@8727.4]
  assign exe_load_inst_0 = exe_wire_0_mem_en & _T_1047; // @[BackEnd.scala 397:44:@8728.4]
  assign _T_1056 = _T_1055 & exe_load_inst_0; // @[BackEnd.scala 401:89:@8737.4]
  assign rs2_addr_N0_0 = InstDecoder_io_cinfo_rs2_addr != 5'h0; // @[BackEnd.scala 399:47:@8732.4]
  assign _T_1058 = _T_568 & rs2_addr_N0_0; // @[BackEnd.scala 402:48:@8739.4]
  assign _T_1059 = _T_1058 & dec_wire_0_rs2_oen; // @[BackEnd.scala 402:66:@8740.4]
  assign _T_1060 = _T_1059 & exe_load_inst_0; // @[BackEnd.scala 402:89:@8741.4]
  assign _T_1061 = _T_1056 | _T_1060; // @[BackEnd.scala 401:110:@8742.4]
  assign _T_1063 = _T_548 & rs1_addr_N0_0; // @[BackEnd.scala 403:48:@8744.4]
  assign _T_1064 = _T_1063 & dec_wire_0_rs1_oen; // @[BackEnd.scala 403:66:@8745.4]
  assign _T_1072 = exe_1_mem_fcn == 1'h0; // @[BackEnd.scala 397:62:@8754.4]
  assign exe_load_inst_1 = exe_wire_1_mem_en & _T_1072; // @[BackEnd.scala 397:44:@8755.4]
  assign _T_1065 = _T_1064 & exe_load_inst_1; // @[BackEnd.scala 403:89:@8746.4]
  assign _T_1066 = _T_1061 | _T_1065; // @[BackEnd.scala 402:110:@8747.4]
  assign _T_1068 = _T_566 & rs2_addr_N0_0; // @[BackEnd.scala 404:48:@8749.4]
  assign _T_1069 = _T_1068 & dec_wire_0_rs2_oen; // @[BackEnd.scala 404:66:@8750.4]
  assign _T_1070 = _T_1069 & exe_load_inst_1; // @[BackEnd.scala 404:89:@8751.4]
  assign rAW_0 = _T_1066 | _T_1070; // @[BackEnd.scala 403:110:@8752.4]
  assign exe_wire_0_csr_cmd = exe_valid_0 ? exe_0_csr_cmd : 3'h0; // @[BackEnd.scala 213:31:@8251.4]
  assign _T_1097 = exe_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 407:56:@8781.4]
  assign _T_1098 = rAW_0 | _T_1097; // @[BackEnd.scala 407:33:@8782.4]
  assign exe_wire_1_csr_cmd = exe_valid_1 ? exe_1_csr_cmd : 3'h0; // @[BackEnd.scala 213:31:@8290.4]
  assign _T_1099 = exe_wire_1_csr_cmd != 3'h0; // @[BackEnd.scala 407:89:@8783.4]
  assign stall_0_0 = _T_1098 | _T_1099; // @[BackEnd.scala 407:66:@8784.4]
  assign _T_696 = stall_0_0 | stall_1_1; // @[BackEnd.scala 192:31:@8202.4]
  assign _T_702 = _T_696 & _T_601; // @[BackEnd.scala 192:79:@8206.4]
  assign ma_jump = mem_sel_0 ? mem_wire_jump_0 : mem_wire_jump_1; // @[BackEnd.scala 344:29:@8602.4]
  assign mem_en = mem_sel_0 ? mem_wire_0_mem_en : mem_wire_1_mem_en; // @[BackEnd.scala 326:25:@8490.4]
  assign mem_fcn = mem_sel_0 ? mem_0_mem_fcn : mem_1_mem_fcn; // @[BackEnd.scala 327:25:@8491.4]
  assign _T_907 = mem_fcn == 1'h0; // @[BackEnd.scala 342:44:@8596.4]
  assign _T_908 = mem_en & _T_907; // @[BackEnd.scala 342:33:@8597.4]
  assign mem_typ = mem_sel_0 ? mem_0_mem_typ : mem_1_mem_typ; // @[BackEnd.scala 328:25:@8492.4]
  assign _T_896 = mem_typ[1:0]; // @[BackEnd.scala 337:43:@8588.4]
  assign _T_906 = 2'h2 == _T_896; // @[Mux.scala 46:19:@8594.4]
  assign mem_exe_out = mem_sel_0 ? mem_reg_wbdata_0 : mem_reg_wbdata_1; // @[BackEnd.scala 322:25:@8486.4]
  assign _T_899 = mem_exe_out[0]; // @[BackEnd.scala 338:23:@8589.4]
  assign _T_904 = 2'h3 == _T_896; // @[Mux.scala 46:19:@8592.4]
  assign _T_901 = mem_exe_out[1:0]; // @[BackEnd.scala 339:23:@8590.4]
  assign _T_903 = _T_901 != 2'h0; // @[BackEnd.scala 339:29:@8591.4]
  assign _T_905 = _T_904 ? _T_903 : 1'h0; // @[Mux.scala 46:16:@8593.4]
  assign ls_addr_ma_valid = _T_906 ? _T_899 : _T_905; // @[Mux.scala 46:16:@8595.4]
  assign ma_load = _T_908 & ls_addr_ma_valid; // @[BackEnd.scala 342:54:@8598.4]
  assign _T_928 = ma_jump | ma_load; // @[BackEnd.scala 359:25:@8618.4]
  assign _T_910 = mem_en & mem_fcn; // @[BackEnd.scala 343:33:@8600.4]
  assign ma_store = _T_910 & ls_addr_ma_valid; // @[BackEnd.scala 343:54:@8601.4]
  assign _T_929 = _T_928 | ma_store; // @[BackEnd.scala 359:36:@8619.4]
  assign ma_illegal = mem_sel_0 ? mem_wire_0_illegal : mem_wire_1_illegal; // @[BackEnd.scala 345:29:@8603.4]
  assign _T_930 = _T_929 | ma_illegal; // @[BackEnd.scala 359:48:@8620.4]
  assign xcpt_valid = _T_930 | csr_io_eret; // @[BackEnd.scala 359:62:@8621.4]
  assign _T_703 = _T_702 | xcpt_valid; // @[BackEnd.scala 192:104:@8207.4]
  assign not_expect = io_front_feedBack_bits_tgt != exe_pred_tgt; // @[BackEnd.scala 266:53:@8371.4]
  assign exe_wire_0_isBJ = exe_valid_0 & exe_0_isBJ; // @[BackEnd.scala 210:41:@8245.4]
  assign exe_wire_1_isBJ = exe_valid_1 & exe_1_isBJ; // @[BackEnd.scala 210:41:@8284.4]
  assign exe_wire_isBJ = exe_wire_0_isBJ | exe_wire_1_isBJ; // @[BackEnd.scala 245:54:@8321.4]
  assign mispredict = not_expect & exe_wire_isBJ; // @[BackEnd.scala 267:28:@8372.4]
  assign _T_711 = mispredict == 1'h0; // @[BackEnd.scala 195:47:@8216.8]
  assign _T_712 = io_front_inst_0_valid & _T_711; // @[BackEnd.scala 195:44:@8217.8]
  assign _GEN_38 = _T_602 ? _T_712 : exe_valid_0; // @[BackEnd.scala 194:60:@8215.6]
  assign _GEN_39 = _T_703 ? 1'h0 : _GEN_38; // @[BackEnd.scala 192:119:@8208.4]
  assign _T_1101 = InstDecoder_io_cinfo_wbaddr == InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 410:26:@8786.4]
  assign rs1_addr_N0_1 = InstDecoder_1_io_cinfo_rs1_addr != 5'h0; // @[BackEnd.scala 398:47:@8757.4]
  assign _T_1102 = _T_1101 & rs1_addr_N0_1; // @[BackEnd.scala 410:52:@8787.4]
  assign _T_1103 = _T_1102 & dec_wire_1_rs1_oen; // @[BackEnd.scala 410:70:@8788.4]
  assign _T_1104 = _T_1103 & dec_wire_0_rf_wen; // @[BackEnd.scala 410:93:@8789.4]
  assign _T_1105 = InstDecoder_io_cinfo_wbaddr == InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 411:26:@8790.4]
  assign rs2_addr_N0_1 = InstDecoder_1_io_cinfo_rs2_addr != 5'h0; // @[BackEnd.scala 399:47:@8759.4]
  assign _T_1106 = _T_1105 & rs2_addr_N0_1; // @[BackEnd.scala 411:52:@8791.4]
  assign _T_1107 = _T_1106 & dec_wire_1_rs2_oen; // @[BackEnd.scala 411:70:@8792.4]
  assign _T_1108 = _T_1107 & dec_wire_0_rf_wen; // @[BackEnd.scala 411:93:@8793.4]
  assign _T_1109 = _T_1104 | _T_1108; // @[BackEnd.scala 410:116:@8794.4]
  assign _T_1110 = dec_wire_0_csr_cmd != 3'h0; // @[BackEnd.scala 412:25:@8795.4]
  assign _T_1111 = _T_1109 | _T_1110; // @[BackEnd.scala 411:116:@8796.4]
  assign _T_1079 = _T_621 & rs1_addr_N0_1; // @[BackEnd.scala 401:48:@8762.4]
  assign _T_1080 = _T_1079 & dec_wire_1_rs1_oen; // @[BackEnd.scala 401:66:@8763.4]
  assign _T_1081 = _T_1080 & exe_load_inst_0; // @[BackEnd.scala 401:89:@8764.4]
  assign _T_1083 = _T_639 & rs2_addr_N0_1; // @[BackEnd.scala 402:48:@8766.4]
  assign _T_1084 = _T_1083 & dec_wire_1_rs2_oen; // @[BackEnd.scala 402:66:@8767.4]
  assign _T_1085 = _T_1084 & exe_load_inst_0; // @[BackEnd.scala 402:89:@8768.4]
  assign _T_1086 = _T_1081 | _T_1085; // @[BackEnd.scala 401:110:@8769.4]
  assign _T_1088 = _T_619 & rs1_addr_N0_1; // @[BackEnd.scala 403:48:@8771.4]
  assign _T_1089 = _T_1088 & dec_wire_1_rs1_oen; // @[BackEnd.scala 403:66:@8772.4]
  assign _T_1090 = _T_1089 & exe_load_inst_1; // @[BackEnd.scala 403:89:@8773.4]
  assign _T_1091 = _T_1086 | _T_1090; // @[BackEnd.scala 402:110:@8774.4]
  assign _T_1093 = _T_637 & rs2_addr_N0_1; // @[BackEnd.scala 404:48:@8776.4]
  assign _T_1094 = _T_1093 & dec_wire_1_rs2_oen; // @[BackEnd.scala 404:66:@8777.4]
  assign _T_1095 = _T_1094 & exe_load_inst_1; // @[BackEnd.scala 404:89:@8778.4]
  assign rAW_1 = _T_1091 | _T_1095; // @[BackEnd.scala 403:110:@8779.4]
  assign _T_1112 = _T_1111 | rAW_1; // @[BackEnd.scala 412:35:@8797.4]
  assign stall_1_0 = _T_1112 | stall_0_0; // @[BackEnd.scala 412:45:@8798.4]
  assign _T_715 = stall_1_0 & _T_599; // @[BackEnd.scala 198:30:@8221.4]
  assign _T_718 = _T_715 & _T_601; // @[BackEnd.scala 198:54:@8223.4]
  assign _T_719 = _T_718 | xcpt_valid; // @[BackEnd.scala 198:79:@8224.4]
  assign exe_cancel = not_expect & exe_wire_0_isBJ; // @[BackEnd.scala 268:28:@8374.4]
  assign _T_720 = _T_719 | exe_cancel; // @[BackEnd.scala 198:93:@8225.4]
  assign _T_729 = io_front_inst_1_valid & _T_711; // @[BackEnd.scala 201:44:@8235.8]
  assign _GEN_40 = _T_602 ? _T_729 : exe_valid_1; // @[BackEnd.scala 200:60:@8233.6]
  assign _GEN_41 = _T_720 ? 1'h0 : _GEN_40; // @[BackEnd.scala 198:108:@8226.4]
  assign target_brjmp = exe_wire_0_isBJ ? ALU_io_target_brjmp : ALU_1_io_target_brjmp; // @[BackEnd.scala 241:19:@8317.4]
  assign target_jpreg = exe_wire_0_isBJ ? ALU_io_target_jpreg : ALU_1_io_target_jpreg; // @[BackEnd.scala 241:19:@8317.4]
  assign target_conti = exe_wire_0_isBJ ? ALU_io_target_conti : ALU_1_io_target_conti; // @[BackEnd.scala 241:19:@8317.4]
  assign pc_sel = exe_wire_0_isBJ ? ALU_io_ctrl_pc_sel : ALU_1_io_ctrl_pc_sel; // @[BackEnd.scala 242:19:@8318.4]
  assign exe_wire_branch = exe_wire_isBJ & exe_reg_branch; // @[BackEnd.scala 246:39:@8322.4]
  assign exe_wire_pop = exe_wire_isBJ & exe_reg_pop; // @[BackEnd.scala 247:39:@8323.4]
  assign exe_wire_push = exe_wire_isBJ & exe_reg_push; // @[BackEnd.scala 248:39:@8324.4]
  assign _GEN_66 = exe_wire_pop ? 1'h0 : _T_766; // @[BackEnd.scala 68:20:@8331.6]
  assign _GEN_67 = _T_601 ? 1'h1 : _GEN_66; // @[BackEnd.scala 67:20:@8327.4]
  assign _GEN_68 = exe_wire_push ? 1'h0 : _T_774; // @[BackEnd.scala 68:20:@8342.6]
  assign _GEN_69 = _T_601 ? 1'h1 : _GEN_68; // @[BackEnd.scala 67:20:@8338.4]
  assign _GEN_70 = exe_wire_isBJ ? 1'h0 : _T_782; // @[BackEnd.scala 68:20:@8354.6]
  assign _GEN_71 = _T_601 ? 1'h1 : _GEN_70; // @[BackEnd.scala 67:20:@8350.4]
  assign _T_786 = pc_sel == 2'h1; // @[BackEnd.scala 255:45:@8359.4]
  assign _T_787 = pc_sel == 2'h2; // @[BackEnd.scala 255:68:@8360.4]
  assign _T_791 = _T_787 ? target_jpreg : target_conti; // @[BackEnd.scala 258:10:@8365.4]
  assign _T_796 = exe_wire_pop ? 2'h1 : 2'h3; // @[BackEnd.scala 264:10:@8368.4]
  assign _T_808 = _T_786 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@8381.6]
  assign _T_809 = _T_808 & target_brjmp; // @[BackEnd.scala 273:47:@8382.6]
  assign _T_814 = _T_787 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@8385.6]
  assign _T_815 = _T_814 & target_jpreg; // @[BackEnd.scala 274:47:@8386.6]
  assign _T_816 = _T_809 | _T_815; // @[BackEnd.scala 273:63:@8387.6]
  assign _GEN_72 = _T_601 ? _T_816 : mem_reg_jpnpc; // @[BackEnd.scala 271:31:@8378.4]
  assign _T_819 = stall_0_2 == 1'h0; // @[BackEnd.scala 277:57:@8391.4]
  assign _T_820 = stall_1_2 & _T_819; // @[BackEnd.scala 277:54:@8392.4]
  assign _T_821 = _T_820 | xcpt_valid; // @[BackEnd.scala 277:78:@8393.4]
  assign _GEN_73 = _T_601 ? exe_valid_0 : mem_valid_0; // @[BackEnd.scala 279:37:@8399.6]
  assign _GEN_74 = _T_821 ? 1'h0 : _GEN_73; // @[BackEnd.scala 277:93:@8394.4]
  assign _T_827 = stall_1_1 & _T_601; // @[BackEnd.scala 283:30:@8403.4]
  assign _T_828 = _T_827 | xcpt_valid; // @[BackEnd.scala 283:55:@8404.4]
  assign _T_833 = exe_cancel == 1'h0; // @[BackEnd.scala 286:37:@8411.8]
  assign _T_834 = exe_valid_1 & _T_833; // @[BackEnd.scala 286:34:@8412.8]
  assign _GEN_75 = _T_601 ? _T_834 : mem_valid_1; // @[BackEnd.scala 285:37:@8410.6]
  assign _GEN_76 = _T_828 ? 1'h0 : _GEN_75; // @[BackEnd.scala 283:70:@8405.4]
  assign _T_837 = exe_wire_1_mem_en & _T_833; // @[BackEnd.scala 289:69:@8416.4]
  assign mem_inst = mem_sel_0 ? mem_0_inst : mem_1_inst; // @[BackEnd.scala 321:25:@8485.4]
  assign _T_911 = ma_load | ma_store; // @[BackEnd.scala 346:27:@8604.4]
  assign _T_912 = _T_911 | ma_jump; // @[BackEnd.scala 346:39:@8605.4]
  assign _T_919 = ma_store ? 3'h6 : 3'h0; // @[Mux.scala 61:16:@8608.4]
  assign _T_920 = ma_load ? 3'h4 : _T_919; // @[Mux.scala 61:16:@8609.4]
  assign _T_921 = ma_illegal ? 3'h2 : _T_920; // @[Mux.scala 61:16:@8610.4]
  assign _T_922 = ma_jump ? 3'h0 : _T_921; // @[Mux.scala 61:16:@8611.4]
  assign _T_924 = ma_store ? mem_exe_out : 32'h0; // @[Mux.scala 61:16:@8613.4]
  assign _T_925 = ma_load ? mem_exe_out : _T_924; // @[Mux.scala 61:16:@8614.4]
  assign _T_926 = ma_illegal ? mem_inst : _T_925; // @[Mux.scala 61:16:@8615.4]
  assign _T_932 = xcpt_valid & mem_sel_0; // @[BackEnd.scala 362:44:@8624.4]
  assign _T_933 = stall_0_2 | _T_932; // @[BackEnd.scala 362:29:@8625.4]
  assign _GEN_77 = _T_933 ? 1'h0 : mem_valid_0; // @[BackEnd.scala 362:60:@8626.4]
  assign _T_935 = stall_1_2 | xcpt_valid; // @[BackEnd.scala 366:29:@8632.4]
  assign _GEN_78 = _T_935 ? 1'h0 : mem_valid_1; // @[BackEnd.scala 366:44:@8633.4]
  assign _T_952 = {wb_valid_1,wb_valid_0}; // @[BackEnd.scala 385:25:@8654.4]
  assign retire_0 = ^_T_952; // @[BackEnd.scala 385:32:@8655.4]
  assign _T_955 = ~ _T_952; // @[BackEnd.scala 386:32:@8658.4]
  assign retire_1 = _T_955 == 2'h0; // @[BackEnd.scala 386:32:@8659.4]
  assign _GEN_79 = mispredict ? 1'h0 : _T_1133; // @[BackEnd.scala 68:20:@8821.6]
  assign _GEN_80 = _T_601 ? 1'h1 : _GEN_79; // @[BackEnd.scala 67:20:@8817.4]
  assign _T_1138 = stall_0_0 == 1'h0; // @[BackEnd.scala 421:26:@8828.4]
  assign _T_1141 = _T_1138 & _T_599; // @[BackEnd.scala 421:47:@8830.4]
  assign _T_1146 = stall_1_0 == 1'h0; // @[BackEnd.scala 422:26:@8834.4]
  assign _T_1149 = _T_1146 & _T_599; // @[BackEnd.scala 422:47:@8836.4]
  assign _T_1152 = _T_1149 & _T_601; // @[BackEnd.scala 422:71:@8838.4]
  assign _T_1153 = dec_wire_0_isBJ & dec_wire_1_isBJ; // @[BackEnd.scala 423:35:@8839.4]
  assign _T_1155 = _T_1153 == 1'h0; // @[BackEnd.scala 423:5:@8840.4]
  assign _T_1159 = stall_0_2 ? 8'h4d : 8'h20; // @[BackEnd.scala 432:12:@8843.4]
  assign _T_1167 = stall_0_0 ? 8'h44 : 8'h20; // @[BackEnd.scala 434:12:@8845.4]
  assign _T_1170 = ALU_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 435:32:@8846.4]
  assign _T_1173 = ALU_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 436:32:@8847.4]
  assign _T_1176 = ALU_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 437:32:@8848.4]
  assign _T_1179 = ALU_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 438:32:@8849.4]
  assign _T_1182 = _T_1179 ? 8'h20 : 8'h3f; // @[BackEnd.scala 438:12:@8850.4]
  assign _T_1183 = _T_1176 ? 8'h45 : _T_1182; // @[BackEnd.scala 437:12:@8851.4]
  assign _T_1184 = _T_1173 ? 8'h4a : _T_1183; // @[BackEnd.scala 436:12:@8852.4]
  assign _T_1185 = _T_1170 ? 8'h42 : _T_1184; // @[BackEnd.scala 435:12:@8853.4]
  assign _T_1189 = csr_io_illegal ? 8'h58 : 8'h20; // @[BackEnd.scala 439:12:@8854.4]
  assign _T_1192 = exe_valid_0 == 1'h0; // @[BackEnd.scala 440:13:@8855.4]
  assign _T_1193 = _T_1192 | xcpt_valid; // @[BackEnd.scala 440:27:@8856.4]
  assign _T_1199 = _T_1193 | stall_1_2; // @[BackEnd.scala 440:72:@8860.4]
  assign _T_1205 = _T_1199 ? 32'h4033 : exe_0_inst; // @[BackEnd.scala 440:12:@8864.4]
  assign _T_1208 = reset == 1'h0; // @[BackEnd.scala 427:11:@8866.4]
  assign _T_1211 = stall_1_2 ? 8'h4d : 8'h20; // @[BackEnd.scala 432:12:@8870.4]
  assign _T_1215 = stall_1_1 ? 8'h45 : 8'h20; // @[BackEnd.scala 433:12:@8871.4]
  assign _T_1219 = stall_1_0 ? 8'h44 : 8'h20; // @[BackEnd.scala 434:12:@8872.4]
  assign _T_1222 = ALU_1_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 435:32:@8873.4]
  assign _T_1225 = ALU_1_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 436:32:@8874.4]
  assign _T_1228 = ALU_1_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 437:32:@8875.4]
  assign _T_1231 = ALU_1_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 438:32:@8876.4]
  assign _T_1234 = _T_1231 ? 8'h20 : 8'h3f; // @[BackEnd.scala 438:12:@8877.4]
  assign _T_1235 = _T_1228 ? 8'h45 : _T_1234; // @[BackEnd.scala 437:12:@8878.4]
  assign _T_1236 = _T_1225 ? 8'h4a : _T_1235; // @[BackEnd.scala 436:12:@8879.4]
  assign _T_1237 = _T_1222 ? 8'h42 : _T_1236; // @[BackEnd.scala 435:12:@8880.4]
  assign _T_1244 = exe_valid_1 == 1'h0; // @[BackEnd.scala 440:13:@8882.4]
  assign _T_1245 = _T_1244 | xcpt_valid; // @[BackEnd.scala 440:27:@8883.4]
  assign _T_1250 = _T_1245 | exe_cancel; // @[BackEnd.scala 440:41:@8886.4]
  assign _T_1251 = _T_1250 | stall_1_2; // @[BackEnd.scala 440:72:@8887.4]
  assign _T_1256 = _T_1251 | stall_1_1; // @[BackEnd.scala 441:29:@8890.4]
  assign _T_1257 = _T_1256 ? 32'h4033 : exe_1_inst; // @[BackEnd.scala 440:12:@8891.4]
  assign _T_1267 = exe_pred_tgt != target_conti; // @[BackEnd.scala 462:22:@8912.6]
  assign _T_1268 = exe_wire_0_isBJ ? exe_0_inst : exe_1_inst; // @[BackEnd.scala 463:12:@8913.6]
  assign io_mem_req_valid = exe_wire_0_mem_en | _T_837; // @[BackEnd.scala 289:24:@8418.4]
  assign io_mem_req_bits_addr = exe_wire_0_mem_en ? exe_wbdata_0 : exe_wbdata_1; // @[BackEnd.scala 290:24:@8420.4]
  assign io_mem_req_bits_data = exe_wire_0_mem_en ? exe_0_rs2_data : exe_1_rs2_data; // @[BackEnd.scala 293:24:@8426.4]
  assign io_mem_req_bits_fcn = exe_wire_0_mem_en ? exe_0_mem_fcn : exe_1_mem_fcn; // @[BackEnd.scala 291:24:@8422.4]
  assign io_mem_req_bits_typ = exe_wire_0_mem_en ? exe_0_mem_typ : exe_1_mem_typ; // @[BackEnd.scala 292:24:@8424.4]
  assign io_cyc = csr_io_time; // @[BackEnd.scala 84:10:@7946.4]
  assign io_front_xcpt_valid = _T_930 | csr_io_eret; // @[BackEnd.scala 420:17:@8827.4]
  assign io_front_xcpt_bits = csr_io_evec; // @[BackEnd.scala 420:17:@8826.4]
  assign io_front_kill = mispredict & _T_1133; // @[BackEnd.scala 419:17:@8825.4]
  assign io_front_fence = _T_473 | _T_474; // @[BackEnd.scala 100:20:@7971.4]
  assign io_front_ras_pop = exe_wire_pop & _T_766; // @[BackEnd.scala 250:27:@8335.4]
  assign io_front_ras_push_valid = exe_wire_push & _T_774; // @[BackEnd.scala 251:27:@8346.4]
  assign io_front_ras_push_bits = exe_wire_0_isBJ ? ALU_io_target_conti : ALU_1_io_target_conti; // @[BackEnd.scala 252:27:@8347.4]
  assign io_front_fb_pc = exe_wire_0_isBJ ? exe_0_pc : exe_1_pc; // @[BackEnd.scala 243:18:@8320.4]
  assign io_front_fb_type = exe_wire_branch ? 2'h2 : _T_796; // @[BackEnd.scala 262:20:@8370.4]
  assign io_front_feedBack_valid = exe_wire_isBJ & _T_782; // @[BackEnd.scala 254:27:@8358.4]
  assign io_front_feedBack_bits_redirect = _T_786 | _T_787; // @[BackEnd.scala 255:35:@8362.4]
  assign io_front_feedBack_bits_tgt = _T_786 ? target_brjmp : _T_791; // @[BackEnd.scala 256:30:@8367.4]
  assign io_front_forward_0 = _T_1141 & _T_601; // @[BackEnd.scala 421:23:@8833.4]
  assign io_front_forward_1 = _T_1152 & _T_1155; // @[BackEnd.scala 422:23:@8842.4]
  assign csr_clock = clock; // @[:@7928.4]
  assign csr_reset = reset; // @[:@7929.4]
  assign csr_io_rw_cmd = mem_sel_0 ? mem_wire_0_csr_cmd : mem_wire_1_csr_cmd; // @[BackEnd.scala 334:19:@8586.4]
  assign csr_io_rw_addr = mem_inst[31:20]; // @[BackEnd.scala 332:19:@8584.4]
  assign csr_io_rw_wdata = mem_sel_0 ? mem_reg_wbdata_0 : mem_reg_wbdata_1; // @[BackEnd.scala 333:19:@8585.4]
  assign csr_io_xcpt = _T_912 | ma_illegal; // @[BackEnd.scala 346:16:@8607.4]
  assign csr_io_cause = {{29'd0}, _T_922}; // @[BackEnd.scala 347:16:@8612.4]
  assign csr_io_tval = ma_jump ? mem_reg_jpnpc : _T_926; // @[BackEnd.scala 353:16:@8617.4]
  assign csr_io_illegal = 1'h0;
  assign csr_io_retire = {retire_1,retire_0}; // @[BackEnd.scala 387:17:@8662.4]
  assign csr_io_pc = mem_sel_0 ? mem_0_pc : mem_1_pc; // @[BackEnd.scala 335:19:@8587.4]
  assign regfile_clock = clock; // @[:@7931.4]
  assign regfile_io_rs1_addr_0 = InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 123:28:@7996.4]
  assign regfile_io_rs1_addr_1 = InstDecoder_1_io_cinfo_rs1_addr; // @[BackEnd.scala 123:28:@8097.4]
  assign regfile_io_rs2_addr_0 = InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 124:28:@7997.4]
  assign regfile_io_rs2_addr_1 = InstDecoder_1_io_cinfo_rs2_addr; // @[BackEnd.scala 124:28:@8098.4]
  assign regfile_io_waddr_0 = wb_0_wbaddr; // @[BackEnd.scala 374:25:@8643.4]
  assign regfile_io_waddr_1 = wb_1_wbaddr; // @[BackEnd.scala 374:25:@8650.4]
  assign regfile_io_wdata_0 = wb_wbdata_0; // @[BackEnd.scala 375:25:@8644.4]
  assign regfile_io_wdata_1 = wb_wbdata_1; // @[BackEnd.scala 375:25:@8651.4]
  assign regfile_io_wen_0 = _T_937 & _T_939; // @[BackEnd.scala 376:25:@8645.4]
  assign regfile_io_wen_1 = _T_941 & _T_943; // @[BackEnd.scala 376:25:@8652.4]
  assign ALU_io_op1 = exe_0_op1_data; // @[BackEnd.scala 216:25:@8255.4]
  assign ALU_io_op2 = exe_0_op2_data; // @[BackEnd.scala 217:25:@8256.4]
  assign ALU_io_pc = exe_0_pc; // @[BackEnd.scala 218:25:@8257.4]
  assign ALU_io_ctrl_fun = exe_0_alu_fun; // @[BackEnd.scala 220:25:@8259.4]
  assign ALU_io_ctrl_br_type = exe_valid_0 ? exe_0_br_type : 4'h0; // @[BackEnd.scala 221:25:@8260.4]
  assign ALU_io_ctrl_wb_sel = exe_0_wb_sel; // @[BackEnd.scala 222:25:@8261.4]
  assign ALU_io_rs2_data = exe_0_rs2_data; // @[BackEnd.scala 219:25:@8258.4]
  assign ALU_1_io_op1 = exe_1_op1_data; // @[BackEnd.scala 216:25:@8294.4]
  assign ALU_1_io_op2 = exe_1_op2_data; // @[BackEnd.scala 217:25:@8295.4]
  assign ALU_1_io_pc = exe_1_pc; // @[BackEnd.scala 218:25:@8296.4]
  assign ALU_1_io_ctrl_fun = exe_1_alu_fun; // @[BackEnd.scala 220:25:@8298.4]
  assign ALU_1_io_ctrl_br_type = exe_valid_1 ? exe_1_br_type : 4'h0; // @[BackEnd.scala 221:25:@8299.4]
  assign ALU_1_io_ctrl_wb_sel = exe_1_wb_sel; // @[BackEnd.scala 222:25:@8300.4]
  assign ALU_1_io_rs2_data = exe_1_rs2_data; // @[BackEnd.scala 219:25:@8297.4]
  assign InstDecoder_io_inst = io_front_inst_0_bits; // @[BackEnd.scala 115:18:@7981.4]
  assign InstDecoder_1_io_inst = io_front_inst_1_bits; // @[BackEnd.scala 115:18:@8082.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exe_0_rf_wen = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  exe_0_wbaddr = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  exe_0_mem_en = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  exe_0_csr_cmd = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  exe_0_illegal = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  exe_0_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  exe_0_inst = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  exe_0_rs2_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  exe_0_wb_sel = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  exe_0_mem_fcn = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  exe_0_mem_typ = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  exe_0_fencei = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  exe_0_br_type = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  exe_0_isBJ = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  exe_0_op1_data = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  exe_0_op2_data = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  exe_0_alu_fun = _RAND_16[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  exe_1_rf_wen = _RAND_17[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  exe_1_wbaddr = _RAND_18[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  exe_1_mem_en = _RAND_19[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  exe_1_csr_cmd = _RAND_20[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  exe_1_illegal = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  exe_1_pc = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  exe_1_inst = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  exe_1_rs2_data = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  exe_1_wb_sel = _RAND_25[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  exe_1_mem_fcn = _RAND_26[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  exe_1_mem_typ = _RAND_27[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  exe_1_fencei = _RAND_28[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  exe_1_br_type = _RAND_29[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  exe_1_isBJ = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  exe_1_op1_data = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  exe_1_op2_data = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  exe_1_alu_fun = _RAND_33[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  exe_valid_0 = _RAND_34[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  exe_valid_1 = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_0_rf_wen = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  mem_0_wbaddr = _RAND_37[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  mem_0_mem_en = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  mem_0_csr_cmd = _RAND_39[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  mem_0_illegal = _RAND_40[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  mem_0_pc = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  mem_0_inst = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  mem_0_wb_sel = _RAND_43[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  mem_0_mem_fcn = _RAND_44[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  mem_0_mem_typ = _RAND_45[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  mem_1_rf_wen = _RAND_46[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  mem_1_wbaddr = _RAND_47[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  mem_1_mem_en = _RAND_48[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  mem_1_csr_cmd = _RAND_49[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  mem_1_illegal = _RAND_50[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  mem_1_pc = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  mem_1_inst = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  mem_1_wb_sel = _RAND_53[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  mem_1_mem_fcn = _RAND_54[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  mem_1_mem_typ = _RAND_55[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  mem_valid_0 = _RAND_56[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  mem_valid_1 = _RAND_57[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  wb_0_rf_wen = _RAND_58[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  wb_0_wbaddr = _RAND_59[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  wb_1_rf_wen = _RAND_60[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  wb_1_wbaddr = _RAND_61[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  wb_valid_0 = _RAND_62[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  wb_valid_1 = _RAND_63[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  wb_wbdata_0 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  wb_wbdata_1 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  mem_reg_wbdata_0 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  mem_reg_wbdata_1 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  mem_reg_jpnpc = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  exe_pred_tgt = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  exe_reg_branch = _RAND_70[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  exe_reg_pop = _RAND_71[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  exe_reg_push = _RAND_72[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  _T_766 = _RAND_73[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  _T_774 = _RAND_74[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  _T_782 = _RAND_75[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  _T_1133 = _RAND_76[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (_T_602) begin
      exe_0_rf_wen <= InstDecoder_io_cinfo_rf_wen;
    end
    if (_T_602) begin
      exe_0_wbaddr <= InstDecoder_io_cinfo_wbaddr;
    end
    if (_T_602) begin
      exe_0_mem_en <= InstDecoder_io_cinfo_mem_en;
    end
    if (_T_602) begin
      if (_T_608) begin
        exe_0_csr_cmd <= 3'h5;
      end else begin
        exe_0_csr_cmd <= InstDecoder_io_cinfo_csr_cmd;
      end
    end
    if (_T_602) begin
      exe_0_illegal <= InstDecoder_io_cinfo_illegal;
    end
    if (_T_602) begin
      exe_0_pc <= io_front_pc_0;
    end
    if (_T_602) begin
      exe_0_inst <= InstDecoder_io_inst;
    end
    if (_T_602) begin
      if (_T_567) begin
        exe_0_rs2_data <= exe_wbdata_1;
      end else begin
        if (_T_569) begin
          exe_0_rs2_data <= exe_wbdata_0;
        end else begin
          if (_T_571) begin
            if (_T_891) begin
              exe_0_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_892) begin
                exe_0_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_0_rs2_data <= mem_reg_wbdata_1;
              end
            end
          end else begin
            if (_T_573) begin
              if (_T_872) begin
                exe_0_rs2_data <= io_mem_resp_bits_data;
              end else begin
                if (_T_873) begin
                  exe_0_rs2_data <= csr_io_rw_rdata;
                end else begin
                  exe_0_rs2_data <= mem_reg_wbdata_0;
                end
              end
            end else begin
              if (_T_575) begin
                exe_0_rs2_data <= wb_wbdata_1;
              end else begin
                if (_T_577) begin
                  exe_0_rs2_data <= wb_wbdata_0;
                end else begin
                  exe_0_rs2_data <= rf_rs2_data_0;
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      exe_0_wb_sel <= InstDecoder_io_cinfo_wb_sel;
    end
    if (_T_602) begin
      exe_0_mem_fcn <= InstDecoder_io_cinfo_mem_fcn;
    end
    if (_T_602) begin
      exe_0_mem_typ <= InstDecoder_io_cinfo_mem_typ;
    end
    if (_T_602) begin
      exe_0_fencei <= InstDecoder_io_cinfo_fencei;
    end
    if (_T_602) begin
      exe_0_br_type <= InstDecoder_io_cinfo_br_type;
    end
    if (_T_602) begin
      exe_0_isBJ <= InstDecoder_io_cinfo_isBJ;
    end
    if (_T_602) begin
      if (_T_584) begin
        exe_0_op1_data <= InstDecoder_io_dinfo_imm_z;
      end else begin
        if (_T_585) begin
          exe_0_op1_data <= io_front_pc_0;
        end else begin
          if (_T_549) begin
            exe_0_op1_data <= exe_wbdata_1;
          end else begin
            if (_T_551) begin
              exe_0_op1_data <= exe_wbdata_0;
            end else begin
              if (_T_553) begin
                if (_T_891) begin
                  exe_0_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_892) begin
                    exe_0_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_0_op1_data <= mem_reg_wbdata_1;
                  end
                end
              end else begin
                if (_T_555) begin
                  if (_T_872) begin
                    exe_0_op1_data <= io_mem_resp_bits_data;
                  end else begin
                    if (_T_873) begin
                      exe_0_op1_data <= csr_io_rw_rdata;
                    end else begin
                      exe_0_op1_data <= mem_reg_wbdata_0;
                    end
                  end
                end else begin
                  if (_T_557) begin
                    exe_0_op1_data <= wb_wbdata_1;
                  end else begin
                    if (_T_559) begin
                      exe_0_op1_data <= wb_wbdata_0;
                    end else begin
                      exe_0_op1_data <= rf_rs1_data_0;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      if (_T_588) begin
        exe_0_op2_data <= InstDecoder_io_dinfo_imm_i;
      end else begin
        if (_T_589) begin
          exe_0_op2_data <= InstDecoder_io_dinfo_imm_s;
        end else begin
          if (_T_590) begin
            exe_0_op2_data <= InstDecoder_io_dinfo_imm_sb;
          end else begin
            if (_T_591) begin
              exe_0_op2_data <= InstDecoder_io_dinfo_imm_u;
            end else begin
              if (_T_592) begin
                exe_0_op2_data <= InstDecoder_io_dinfo_imm_uj;
              end else begin
                if (_T_567) begin
                  exe_0_op2_data <= exe_wbdata_1;
                end else begin
                  if (_T_569) begin
                    exe_0_op2_data <= exe_wbdata_0;
                  end else begin
                    if (_T_571) begin
                      if (_T_891) begin
                        exe_0_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_892) begin
                          exe_0_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_0_op2_data <= mem_reg_wbdata_1;
                        end
                      end
                    end else begin
                      if (_T_573) begin
                        if (_T_872) begin
                          exe_0_op2_data <= io_mem_resp_bits_data;
                        end else begin
                          if (_T_873) begin
                            exe_0_op2_data <= csr_io_rw_rdata;
                          end else begin
                            exe_0_op2_data <= mem_reg_wbdata_0;
                          end
                        end
                      end else begin
                        if (_T_575) begin
                          exe_0_op2_data <= wb_wbdata_1;
                        end else begin
                          if (_T_577) begin
                            exe_0_op2_data <= wb_wbdata_0;
                          end else begin
                            exe_0_op2_data <= rf_rs2_data_0;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      exe_0_alu_fun <= InstDecoder_io_cinfo_alu_fun;
    end
    if (_T_602) begin
      exe_1_rf_wen <= InstDecoder_1_io_cinfo_rf_wen;
    end
    if (_T_602) begin
      exe_1_wbaddr <= InstDecoder_1_io_cinfo_wbaddr;
    end
    if (_T_602) begin
      exe_1_mem_en <= InstDecoder_1_io_cinfo_mem_en;
    end
    if (_T_602) begin
      if (_T_679) begin
        exe_1_csr_cmd <= 3'h5;
      end else begin
        exe_1_csr_cmd <= InstDecoder_1_io_cinfo_csr_cmd;
      end
    end
    if (_T_602) begin
      exe_1_illegal <= InstDecoder_1_io_cinfo_illegal;
    end
    if (_T_602) begin
      exe_1_pc <= io_front_pc_1;
    end
    if (_T_602) begin
      exe_1_inst <= InstDecoder_1_io_inst;
    end
    if (_T_602) begin
      if (_T_638) begin
        exe_1_rs2_data <= exe_wbdata_1;
      end else begin
        if (_T_640) begin
          exe_1_rs2_data <= exe_wbdata_0;
        end else begin
          if (_T_642) begin
            if (_T_891) begin
              exe_1_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_892) begin
                exe_1_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_1_rs2_data <= mem_reg_wbdata_1;
              end
            end
          end else begin
            if (_T_644) begin
              if (_T_872) begin
                exe_1_rs2_data <= io_mem_resp_bits_data;
              end else begin
                if (_T_873) begin
                  exe_1_rs2_data <= csr_io_rw_rdata;
                end else begin
                  exe_1_rs2_data <= mem_reg_wbdata_0;
                end
              end
            end else begin
              if (_T_646) begin
                exe_1_rs2_data <= wb_wbdata_1;
              end else begin
                if (_T_648) begin
                  exe_1_rs2_data <= wb_wbdata_0;
                end else begin
                  exe_1_rs2_data <= rf_rs2_data_1;
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      exe_1_wb_sel <= InstDecoder_1_io_cinfo_wb_sel;
    end
    if (_T_602) begin
      exe_1_mem_fcn <= InstDecoder_1_io_cinfo_mem_fcn;
    end
    if (_T_602) begin
      exe_1_mem_typ <= InstDecoder_1_io_cinfo_mem_typ;
    end
    if (_T_602) begin
      exe_1_fencei <= InstDecoder_1_io_cinfo_fencei;
    end
    if (_T_602) begin
      exe_1_br_type <= InstDecoder_1_io_cinfo_br_type;
    end
    if (_T_602) begin
      exe_1_isBJ <= InstDecoder_1_io_cinfo_isBJ;
    end
    if (_T_602) begin
      if (_T_655) begin
        exe_1_op1_data <= InstDecoder_1_io_dinfo_imm_z;
      end else begin
        if (_T_656) begin
          exe_1_op1_data <= io_front_pc_1;
        end else begin
          if (_T_620) begin
            exe_1_op1_data <= exe_wbdata_1;
          end else begin
            if (_T_622) begin
              exe_1_op1_data <= exe_wbdata_0;
            end else begin
              if (_T_624) begin
                if (_T_891) begin
                  exe_1_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_892) begin
                    exe_1_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_1_op1_data <= mem_reg_wbdata_1;
                  end
                end
              end else begin
                if (_T_626) begin
                  if (_T_872) begin
                    exe_1_op1_data <= io_mem_resp_bits_data;
                  end else begin
                    if (_T_873) begin
                      exe_1_op1_data <= csr_io_rw_rdata;
                    end else begin
                      exe_1_op1_data <= mem_reg_wbdata_0;
                    end
                  end
                end else begin
                  if (_T_628) begin
                    exe_1_op1_data <= wb_wbdata_1;
                  end else begin
                    if (_T_630) begin
                      exe_1_op1_data <= wb_wbdata_0;
                    end else begin
                      exe_1_op1_data <= rf_rs1_data_1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      if (_T_659) begin
        exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_i;
      end else begin
        if (_T_660) begin
          exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_s;
        end else begin
          if (_T_661) begin
            exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_sb;
          end else begin
            if (_T_662) begin
              exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_u;
            end else begin
              if (_T_663) begin
                exe_1_op2_data <= InstDecoder_1_io_dinfo_imm_uj;
              end else begin
                if (_T_638) begin
                  exe_1_op2_data <= exe_wbdata_1;
                end else begin
                  if (_T_640) begin
                    exe_1_op2_data <= exe_wbdata_0;
                  end else begin
                    if (_T_642) begin
                      if (_T_891) begin
                        exe_1_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_892) begin
                          exe_1_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_1_op2_data <= mem_reg_wbdata_1;
                        end
                      end
                    end else begin
                      if (_T_644) begin
                        if (_T_872) begin
                          exe_1_op2_data <= io_mem_resp_bits_data;
                        end else begin
                          if (_T_873) begin
                            exe_1_op2_data <= csr_io_rw_rdata;
                          end else begin
                            exe_1_op2_data <= mem_reg_wbdata_0;
                          end
                        end
                      end else begin
                        if (_T_646) begin
                          exe_1_op2_data <= wb_wbdata_1;
                        end else begin
                          if (_T_648) begin
                            exe_1_op2_data <= wb_wbdata_0;
                          end else begin
                            exe_1_op2_data <= rf_rs2_data_1;
                          end
                        end
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (_T_602) begin
      exe_1_alu_fun <= InstDecoder_1_io_cinfo_alu_fun;
    end
    if (reset) begin
      exe_valid_0 <= 1'h0;
    end else begin
      if (_T_703) begin
        exe_valid_0 <= 1'h0;
      end else begin
        if (_T_602) begin
          exe_valid_0 <= _T_712;
        end
      end
    end
    if (reset) begin
      exe_valid_1 <= 1'h0;
    end else begin
      if (_T_720) begin
        exe_valid_1 <= 1'h0;
      end else begin
        if (_T_602) begin
          exe_valid_1 <= _T_729;
        end
      end
    end
    if (_T_601) begin
      mem_0_rf_wen <= exe_0_rf_wen;
    end
    if (_T_601) begin
      mem_0_wbaddr <= exe_0_wbaddr;
    end
    if (_T_601) begin
      mem_0_mem_en <= exe_0_mem_en;
    end
    if (_T_601) begin
      mem_0_csr_cmd <= exe_0_csr_cmd;
    end
    if (_T_601) begin
      mem_0_illegal <= exe_0_illegal;
    end
    if (_T_601) begin
      mem_0_pc <= exe_0_pc;
    end
    if (_T_601) begin
      mem_0_inst <= exe_0_inst;
    end
    if (_T_601) begin
      mem_0_wb_sel <= exe_0_wb_sel;
    end
    if (_T_601) begin
      mem_0_mem_fcn <= exe_0_mem_fcn;
    end
    if (_T_601) begin
      mem_0_mem_typ <= exe_0_mem_typ;
    end
    if (_T_601) begin
      mem_1_rf_wen <= exe_1_rf_wen;
    end
    if (_T_601) begin
      mem_1_wbaddr <= exe_1_wbaddr;
    end
    if (_T_601) begin
      mem_1_mem_en <= exe_1_mem_en;
    end
    if (_T_601) begin
      mem_1_csr_cmd <= exe_1_csr_cmd;
    end
    if (_T_601) begin
      mem_1_illegal <= exe_1_illegal;
    end
    if (_T_601) begin
      mem_1_pc <= exe_1_pc;
    end
    if (_T_601) begin
      mem_1_inst <= exe_1_inst;
    end
    if (_T_601) begin
      mem_1_wb_sel <= exe_1_wb_sel;
    end
    if (_T_601) begin
      mem_1_mem_fcn <= exe_1_mem_fcn;
    end
    if (_T_601) begin
      mem_1_mem_typ <= exe_1_mem_typ;
    end
    if (reset) begin
      mem_valid_0 <= 1'h0;
    end else begin
      if (_T_821) begin
        mem_valid_0 <= 1'h0;
      end else begin
        if (_T_601) begin
          mem_valid_0 <= exe_valid_0;
        end
      end
    end
    if (reset) begin
      mem_valid_1 <= 1'h0;
    end else begin
      if (_T_828) begin
        mem_valid_1 <= 1'h0;
      end else begin
        if (_T_601) begin
          mem_valid_1 <= _T_834;
        end
      end
    end
    wb_0_rf_wen <= mem_0_rf_wen;
    wb_0_wbaddr <= mem_0_wbaddr;
    wb_1_rf_wen <= mem_1_rf_wen;
    wb_1_wbaddr <= mem_1_wbaddr;
    if (reset) begin
      wb_valid_0 <= 1'h0;
    end else begin
      if (_T_933) begin
        wb_valid_0 <= 1'h0;
      end else begin
        wb_valid_0 <= mem_valid_0;
      end
    end
    if (reset) begin
      wb_valid_1 <= 1'h0;
    end else begin
      if (_T_935) begin
        wb_valid_1 <= 1'h0;
      end else begin
        wb_valid_1 <= mem_valid_1;
      end
    end
    if (_T_872) begin
      wb_wbdata_0 <= io_mem_resp_bits_data;
    end else begin
      if (_T_873) begin
        wb_wbdata_0 <= csr_io_rw_rdata;
      end else begin
        wb_wbdata_0 <= mem_reg_wbdata_0;
      end
    end
    if (_T_891) begin
      wb_wbdata_1 <= io_mem_resp_bits_data;
    end else begin
      if (_T_892) begin
        wb_wbdata_1 <= csr_io_rw_rdata;
      end else begin
        wb_wbdata_1 <= mem_reg_wbdata_1;
      end
    end
    if (_T_601) begin
      mem_reg_wbdata_0 <= exe_wbdata_0;
    end
    if (_T_601) begin
      mem_reg_wbdata_1 <= exe_wbdata_1;
    end
    if (reset) begin
      mem_reg_jpnpc <= 32'h0;
    end else begin
      if (_T_601) begin
        mem_reg_jpnpc <= _T_816;
      end
    end
    if (_T_602) begin
      if (dec_wire_0_isBJ) begin
        exe_pred_tgt <= io_front_pred_0;
      end else begin
        exe_pred_tgt <= io_front_pred_1;
      end
    end
    if (_T_602) begin
      if (dec_wire_0_isBJ) begin
        exe_reg_branch <= InstDecoder_io_cinfo_branch;
      end else begin
        exe_reg_branch <= InstDecoder_1_io_cinfo_branch;
      end
    end
    if (_T_602) begin
      if (dec_wire_0_isBJ) begin
        exe_reg_pop <= InstDecoder_io_cinfo_pop;
      end else begin
        exe_reg_pop <= InstDecoder_1_io_cinfo_pop;
      end
    end
    if (_T_602) begin
      if (dec_wire_0_isBJ) begin
        exe_reg_push <= InstDecoder_io_cinfo_push;
      end else begin
        exe_reg_push <= InstDecoder_1_io_cinfo_push;
      end
    end
    if (reset) begin
      _T_766 <= 1'h1;
    end else begin
      if (_T_601) begin
        _T_766 <= 1'h1;
      end else begin
        if (exe_wire_pop) begin
          _T_766 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_774 <= 1'h1;
    end else begin
      if (_T_601) begin
        _T_774 <= 1'h1;
      end else begin
        if (exe_wire_push) begin
          _T_774 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_782 <= 1'h1;
    end else begin
      if (_T_601) begin
        _T_782 <= 1'h1;
      end else begin
        if (exe_wire_isBJ) begin
          _T_782 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_1133 <= 1'h1;
    end else begin
      if (_T_601) begin
        _T_1133 <= 1'h1;
      end else begin
        if (mispredict) begin
          _T_1133 <= 1'h0;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1208) begin
          $fwrite(32'h80000002,"Core: Cyc= %d PC(%x, %x, %x) [%c%c %c%c %c%c] %c%c %c%c Exe: DASM(%x)\n",io_cyc,io_front_pc_0,exe_0_pc,mem_0_pc,_T_1159,8'h30,8'h20,8'h30,_T_1167,8'h30,_T_1185,8'h30,_T_1189,8'h30,_T_1205); // @[BackEnd.scala 427:11:@8868.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_1208) begin
          $fwrite(32'h80000002,"Core: Cyc= %d PC(%x, %x, %x) [%c%c %c%c %c%c] %c%c %c%c Exe: DASM(%x)\n",io_cyc,io_front_pc_1,exe_1_pc,mem_1_pc,_T_1211,8'h31,_T_1215,8'h31,_T_1219,8'h31,_T_1237,8'h31,_T_1189,8'h31,_T_1257); // @[BackEnd.scala 427:11:@8895.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid_0 & _T_1208) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_0_rf_wen,wb_0_wbaddr,regfile_io_wdata_0); // @[BackEnd.scala 446:13:@8901.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid_1 & _T_1208) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_1_rf_wen,wb_1_wbaddr,regfile_io_wdata_1); // @[BackEnd.scala 446:13:@8908.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_front_feedBack_valid & _T_1208) begin
          $fwrite(32'h80000002,"BranchJump: Cyc= %d kill %x pc %x tgt %x actual %x expect %x inst DASM(%x)\n",io_cyc,mispredict,io_front_fb_pc,io_front_feedBack_bits_tgt,io_front_feedBack_bits_redirect,_T_1267,_T_1268); // @[BackEnd.scala 456:11:@8917.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module rv32_ttoy( // @[:@8921.2]
  input         clock, // @[:@8922.4]
  input         reset, // @[:@8923.4]
  input         io_imem_addr_ready, // @[:@8924.4]
  output        io_imem_addr_valid, // @[:@8924.4]
  output [31:0] io_imem_addr_bits, // @[:@8924.4]
  input         io_imem_inst_0_valid, // @[:@8924.4]
  input  [31:0] io_imem_inst_0_bits, // @[:@8924.4]
  input         io_imem_inst_1_valid, // @[:@8924.4]
  input  [31:0] io_imem_inst_1_bits, // @[:@8924.4]
  output        io_dmem_req_valid, // @[:@8924.4]
  output [31:0] io_dmem_req_bits_addr, // @[:@8924.4]
  output [31:0] io_dmem_req_bits_data, // @[:@8924.4]
  output        io_dmem_req_bits_fcn, // @[:@8924.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:@8924.4]
  input         io_dmem_resp_valid, // @[:@8924.4]
  input  [31:0] io_dmem_resp_bits_data // @[:@8924.4]
);
  wire  frontEnd_clock; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_reset; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_cyc; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_mem_addr_ready; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_mem_addr_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_mem_addr_bits; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_mem_inst_0_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_mem_inst_0_bits; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_mem_inst_1_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_mem_inst_1_bits; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_xcpt_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_xcpt_bits; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_kill; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_fence; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_ras_pop; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_ras_push_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_ras_push_bits; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_fb_pc; // @[Core.scala 35:24:@8926.4]
  wire [1:0] frontEnd_io_back_fb_type; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_feedBack_valid; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_feedBack_bits_redirect; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_feedBack_bits_tgt; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_forward_0; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_forward_1; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_inst_0_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_inst_0_bits; // @[Core.scala 35:24:@8926.4]
  wire  frontEnd_io_back_inst_1_valid; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_inst_1_bits; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_pc_0; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_pc_1; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_pred_0; // @[Core.scala 35:24:@8926.4]
  wire [31:0] frontEnd_io_back_pred_1; // @[Core.scala 35:24:@8926.4]
  wire  backEnd_clock; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_reset; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_mem_req_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_mem_req_bits_addr; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_mem_req_bits_data; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_mem_req_bits_fcn; // @[Core.scala 36:24:@8929.4]
  wire [2:0] backEnd_io_mem_req_bits_typ; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_mem_resp_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_mem_resp_bits_data; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_cyc; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_xcpt_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_xcpt_bits; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_kill; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_fence; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_ras_pop; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_ras_push_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_ras_push_bits; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_fb_pc; // @[Core.scala 36:24:@8929.4]
  wire [1:0] backEnd_io_front_fb_type; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_feedBack_valid; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_feedBack_bits_redirect; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_feedBack_bits_tgt; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_forward_0; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_forward_1; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_inst_0_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_inst_0_bits; // @[Core.scala 36:24:@8929.4]
  wire  backEnd_io_front_inst_1_valid; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_inst_1_bits; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_pc_0; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_pc_1; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_pred_0; // @[Core.scala 36:24:@8929.4]
  wire [31:0] backEnd_io_front_pred_1; // @[Core.scala 36:24:@8929.4]
  FrontEnd frontEnd ( // @[Core.scala 35:24:@8926.4]
    .clock(frontEnd_clock),
    .reset(frontEnd_reset),
    .io_cyc(frontEnd_io_cyc),
    .io_mem_addr_ready(frontEnd_io_mem_addr_ready),
    .io_mem_addr_valid(frontEnd_io_mem_addr_valid),
    .io_mem_addr_bits(frontEnd_io_mem_addr_bits),
    .io_mem_inst_0_valid(frontEnd_io_mem_inst_0_valid),
    .io_mem_inst_0_bits(frontEnd_io_mem_inst_0_bits),
    .io_mem_inst_1_valid(frontEnd_io_mem_inst_1_valid),
    .io_mem_inst_1_bits(frontEnd_io_mem_inst_1_bits),
    .io_back_xcpt_valid(frontEnd_io_back_xcpt_valid),
    .io_back_xcpt_bits(frontEnd_io_back_xcpt_bits),
    .io_back_kill(frontEnd_io_back_kill),
    .io_back_fence(frontEnd_io_back_fence),
    .io_back_ras_pop(frontEnd_io_back_ras_pop),
    .io_back_ras_push_valid(frontEnd_io_back_ras_push_valid),
    .io_back_ras_push_bits(frontEnd_io_back_ras_push_bits),
    .io_back_fb_pc(frontEnd_io_back_fb_pc),
    .io_back_fb_type(frontEnd_io_back_fb_type),
    .io_back_feedBack_valid(frontEnd_io_back_feedBack_valid),
    .io_back_feedBack_bits_redirect(frontEnd_io_back_feedBack_bits_redirect),
    .io_back_feedBack_bits_tgt(frontEnd_io_back_feedBack_bits_tgt),
    .io_back_forward_0(frontEnd_io_back_forward_0),
    .io_back_forward_1(frontEnd_io_back_forward_1),
    .io_back_inst_0_valid(frontEnd_io_back_inst_0_valid),
    .io_back_inst_0_bits(frontEnd_io_back_inst_0_bits),
    .io_back_inst_1_valid(frontEnd_io_back_inst_1_valid),
    .io_back_inst_1_bits(frontEnd_io_back_inst_1_bits),
    .io_back_pc_0(frontEnd_io_back_pc_0),
    .io_back_pc_1(frontEnd_io_back_pc_1),
    .io_back_pred_0(frontEnd_io_back_pred_0),
    .io_back_pred_1(frontEnd_io_back_pred_1)
  );
  BackEnd backEnd ( // @[Core.scala 36:24:@8929.4]
    .clock(backEnd_clock),
    .reset(backEnd_reset),
    .io_mem_req_valid(backEnd_io_mem_req_valid),
    .io_mem_req_bits_addr(backEnd_io_mem_req_bits_addr),
    .io_mem_req_bits_data(backEnd_io_mem_req_bits_data),
    .io_mem_req_bits_fcn(backEnd_io_mem_req_bits_fcn),
    .io_mem_req_bits_typ(backEnd_io_mem_req_bits_typ),
    .io_mem_resp_valid(backEnd_io_mem_resp_valid),
    .io_mem_resp_bits_data(backEnd_io_mem_resp_bits_data),
    .io_cyc(backEnd_io_cyc),
    .io_front_xcpt_valid(backEnd_io_front_xcpt_valid),
    .io_front_xcpt_bits(backEnd_io_front_xcpt_bits),
    .io_front_kill(backEnd_io_front_kill),
    .io_front_fence(backEnd_io_front_fence),
    .io_front_ras_pop(backEnd_io_front_ras_pop),
    .io_front_ras_push_valid(backEnd_io_front_ras_push_valid),
    .io_front_ras_push_bits(backEnd_io_front_ras_push_bits),
    .io_front_fb_pc(backEnd_io_front_fb_pc),
    .io_front_fb_type(backEnd_io_front_fb_type),
    .io_front_feedBack_valid(backEnd_io_front_feedBack_valid),
    .io_front_feedBack_bits_redirect(backEnd_io_front_feedBack_bits_redirect),
    .io_front_feedBack_bits_tgt(backEnd_io_front_feedBack_bits_tgt),
    .io_front_forward_0(backEnd_io_front_forward_0),
    .io_front_forward_1(backEnd_io_front_forward_1),
    .io_front_inst_0_valid(backEnd_io_front_inst_0_valid),
    .io_front_inst_0_bits(backEnd_io_front_inst_0_bits),
    .io_front_inst_1_valid(backEnd_io_front_inst_1_valid),
    .io_front_inst_1_bits(backEnd_io_front_inst_1_bits),
    .io_front_pc_0(backEnd_io_front_pc_0),
    .io_front_pc_1(backEnd_io_front_pc_1),
    .io_front_pred_0(backEnd_io_front_pred_0),
    .io_front_pred_1(backEnd_io_front_pred_1)
  );
  assign io_imem_addr_valid = frontEnd_io_mem_addr_valid; // @[Core.scala 37:19:@8937.4]
  assign io_imem_addr_bits = frontEnd_io_mem_addr_bits; // @[Core.scala 37:19:@8936.4]
  assign io_dmem_req_valid = backEnd_io_mem_req_valid; // @[Core.scala 38:20:@8945.4]
  assign io_dmem_req_bits_addr = backEnd_io_mem_req_bits_addr; // @[Core.scala 38:20:@8944.4]
  assign io_dmem_req_bits_data = backEnd_io_mem_req_bits_data; // @[Core.scala 38:20:@8943.4]
  assign io_dmem_req_bits_fcn = backEnd_io_mem_req_bits_fcn; // @[Core.scala 38:20:@8942.4]
  assign io_dmem_req_bits_typ = backEnd_io_mem_req_bits_typ; // @[Core.scala 38:20:@8941.4]
  assign frontEnd_clock = clock; // @[:@8927.4]
  assign frontEnd_reset = reset; // @[:@8928.4]
  assign frontEnd_io_cyc = backEnd_io_cyc; // @[Core.scala 41:20:@8969.4]
  assign frontEnd_io_mem_addr_ready = io_imem_addr_ready; // @[Core.scala 37:19:@8938.4]
  assign frontEnd_io_mem_inst_0_valid = io_imem_inst_0_valid; // @[Core.scala 37:19:@8933.4]
  assign frontEnd_io_mem_inst_0_bits = io_imem_inst_0_bits; // @[Core.scala 37:19:@8932.4]
  assign frontEnd_io_mem_inst_1_valid = io_imem_inst_1_valid; // @[Core.scala 37:19:@8935.4]
  assign frontEnd_io_mem_inst_1_bits = io_imem_inst_1_bits; // @[Core.scala 37:19:@8934.4]
  assign frontEnd_io_back_xcpt_valid = backEnd_io_front_xcpt_valid; // @[Core.scala 40:20:@8968.4]
  assign frontEnd_io_back_xcpt_bits = backEnd_io_front_xcpt_bits; // @[Core.scala 40:20:@8967.4]
  assign frontEnd_io_back_kill = backEnd_io_front_kill; // @[Core.scala 40:20:@8966.4]
  assign frontEnd_io_back_fence = backEnd_io_front_fence; // @[Core.scala 40:20:@8965.4]
  assign frontEnd_io_back_ras_pop = backEnd_io_front_ras_pop; // @[Core.scala 40:20:@8964.4]
  assign frontEnd_io_back_ras_push_valid = backEnd_io_front_ras_push_valid; // @[Core.scala 40:20:@8963.4]
  assign frontEnd_io_back_ras_push_bits = backEnd_io_front_ras_push_bits; // @[Core.scala 40:20:@8962.4]
  assign frontEnd_io_back_fb_pc = backEnd_io_front_fb_pc; // @[Core.scala 40:20:@8961.4]
  assign frontEnd_io_back_fb_type = backEnd_io_front_fb_type; // @[Core.scala 40:20:@8960.4]
  assign frontEnd_io_back_feedBack_valid = backEnd_io_front_feedBack_valid; // @[Core.scala 40:20:@8959.4]
  assign frontEnd_io_back_feedBack_bits_redirect = backEnd_io_front_feedBack_bits_redirect; // @[Core.scala 40:20:@8958.4]
  assign frontEnd_io_back_feedBack_bits_tgt = backEnd_io_front_feedBack_bits_tgt; // @[Core.scala 40:20:@8957.4]
  assign frontEnd_io_back_forward_0 = backEnd_io_front_forward_0; // @[Core.scala 40:20:@8955.4]
  assign frontEnd_io_back_forward_1 = backEnd_io_front_forward_1; // @[Core.scala 40:20:@8956.4]
  assign backEnd_clock = clock; // @[:@8930.4]
  assign backEnd_reset = reset; // @[:@8931.4]
  assign backEnd_io_mem_resp_valid = io_dmem_resp_valid; // @[Core.scala 38:20:@8940.4]
  assign backEnd_io_mem_resp_bits_data = io_dmem_resp_bits_data; // @[Core.scala 38:20:@8939.4]
  assign backEnd_io_front_inst_0_valid = frontEnd_io_back_inst_0_valid; // @[Core.scala 40:20:@8952.4]
  assign backEnd_io_front_inst_0_bits = frontEnd_io_back_inst_0_bits; // @[Core.scala 40:20:@8951.4]
  assign backEnd_io_front_inst_1_valid = frontEnd_io_back_inst_1_valid; // @[Core.scala 40:20:@8954.4]
  assign backEnd_io_front_inst_1_bits = frontEnd_io_back_inst_1_bits; // @[Core.scala 40:20:@8953.4]
  assign backEnd_io_front_pc_0 = frontEnd_io_back_pc_0; // @[Core.scala 40:20:@8949.4]
  assign backEnd_io_front_pc_1 = frontEnd_io_back_pc_1; // @[Core.scala 40:20:@8950.4]
  assign backEnd_io_front_pred_0 = frontEnd_io_back_pred_0; // @[Core.scala 40:20:@8947.4]
  assign backEnd_io_front_pred_1 = frontEnd_io_back_pred_1; // @[Core.scala 40:20:@8948.4]
endmodule