module FetchInst( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  output        io_mem_req_valid, // @[:@6.4]
  output [31:0] io_mem_req_bits_addr, // @[:@6.4]
  input         io_mem_resp_valid, // @[:@6.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@6.4]
  input         io_if_kill, // @[:@6.4]
  input         io_if_fence, // @[:@6.4]
  input         io_dec_forward, // @[:@6.4]
  input         io_dec_kill, // @[:@6.4]
  input  [31:0] io_if_target, // @[:@6.4]
  input  [31:0] io_btb_target, // @[:@6.4]
  output        io_if_forward, // @[:@6.4]
  output [31:0] io_if_pc, // @[:@6.4]
  output        io_dec_inst_valid, // @[:@6.4]
  output [31:0] io_dec_inst_bits // @[:@6.4]
);
  reg [31:0] if_reg_pc; // @[FetchInst.scala 24:27:@8.4]
  reg [31:0] _RAND_0;
  wire [31:0] if_pc_next; // @[FetchInst.scala 29:22:@11.4]
  wire  _T_144; // @[FetchInst.scala 35:20:@14.4]
  wire [31:0] _GEN_0; // @[FetchInst.scala 35:58:@15.4]
  reg  pc_state; // @[FetchInst.scala 40:25:@18.4]
  reg [31:0] _RAND_1;
  wire  _T_148; // @[FetchInst.scala 41:56:@20.4]
  wire  _T_149; // @[FetchInst.scala 41:53:@21.4]
  wire  _T_151; // @[FetchInst.scala 41:71:@22.4]
  wire  pc_ready; // @[FetchInst.scala 41:68:@23.4]
  wire  inst_yback; // @[FetchInst.scala 42:43:@25.4]
  wire  _T_155; // @[FetchInst.scala 43:46:@27.4]
  wire  inst_nback; // @[FetchInst.scala 43:43:@28.4]
  wire  _T_156; // @[Conditional.scala 37:30:@29.4]
  wire  _GEN_1; // @[FetchInst.scala 45:38:@31.6]
  wire  _GEN_2; // @[FetchInst.scala 48:46:@38.8]
  wire  _GEN_3; // @[Conditional.scala 39:67:@37.6]
  wire  _GEN_4; // @[Conditional.scala 40:58:@30.4]
  wire  _T_161; // @[FetchInst.scala 55:42:@45.4]
  reg [1:0] inst_state; // @[FetchInst.scala 64:27:@53.4]
  reg [31:0] _RAND_2;
  wire  _T_166; // @[Conditional.scala 37:30:@54.4]
  wire  _T_167; // @[FetchInst.scala 67:25:@56.6]
  wire  _T_169; // @[FetchInst.scala 69:18:@61.8]
  wire  _T_170; // @[FetchInst.scala 69:31:@62.8]
  wire  _T_172; // @[FetchInst.scala 69:48:@63.8]
  wire  _T_173; // @[FetchInst.scala 69:45:@64.8]
  wire [1:0] _GEN_5; // @[FetchInst.scala 69:65:@65.8]
  wire [1:0] _GEN_6; // @[FetchInst.scala 67:40:@57.6]
  wire  _T_174; // @[Conditional.scala 37:30:@70.6]
  wire  _T_175; // @[FetchInst.scala 74:28:@72.8]
  wire [1:0] _GEN_7; // @[FetchInst.scala 74:44:@73.8]
  wire  _T_176; // @[Conditional.scala 37:30:@78.8]
  wire [1:0] _GEN_8; // @[FetchInst.scala 79:32:@80.10]
  wire [1:0] _GEN_9; // @[Conditional.scala 39:67:@79.8]
  wire [1:0] _GEN_10; // @[Conditional.scala 39:67:@71.6]
  wire [1:0] _GEN_11; // @[Conditional.scala 40:58:@55.4]
  reg [31:0] reg_inst; // @[FetchInst.scala 84:21:@84.4]
  reg [31:0] _RAND_3;
  wire  _T_178; // @[FetchInst.scala 88:39:@88.4]
  wire  _T_180; // @[FetchInst.scala 89:35:@91.4]
  wire  _T_181; // @[FetchInst.scala 89:45:@92.4]
  assign if_pc_next = io_if_kill ? io_if_target : io_btb_target; // @[FetchInst.scala 29:22:@11.4]
  assign _T_144 = io_if_kill | io_if_forward; // @[FetchInst.scala 35:20:@14.4]
  assign _GEN_0 = _T_144 ? if_pc_next : if_reg_pc; // @[FetchInst.scala 35:58:@15.4]
  assign _T_148 = io_if_kill == 1'h0; // @[FetchInst.scala 41:56:@20.4]
  assign _T_149 = io_dec_forward & _T_148; // @[FetchInst.scala 41:53:@21.4]
  assign _T_151 = io_if_fence == 1'h0; // @[FetchInst.scala 41:71:@22.4]
  assign pc_ready = _T_149 & _T_151; // @[FetchInst.scala 41:68:@23.4]
  assign inst_yback = pc_state & io_mem_resp_valid; // @[FetchInst.scala 42:43:@25.4]
  assign _T_155 = io_mem_resp_valid == 1'h0; // @[FetchInst.scala 43:46:@27.4]
  assign inst_nback = pc_state & _T_155; // @[FetchInst.scala 43:43:@28.4]
  assign _T_156 = 1'h0 == pc_state; // @[Conditional.scala 37:30:@29.4]
  assign _GEN_1 = pc_ready ? 1'h1 : pc_state; // @[FetchInst.scala 45:38:@31.6]
  assign _GEN_2 = io_mem_resp_valid ? pc_ready : pc_state; // @[FetchInst.scala 48:46:@38.8]
  assign _GEN_3 = pc_state ? _GEN_2 : pc_state; // @[Conditional.scala 39:67:@37.6]
  assign _GEN_4 = _T_156 ? _GEN_1 : _GEN_3; // @[Conditional.scala 40:58:@30.4]
  assign _T_161 = io_dec_forward & io_mem_req_valid; // @[FetchInst.scala 55:42:@45.4]
  assign _T_166 = 2'h0 == inst_state; // @[Conditional.scala 37:30:@54.4]
  assign _T_167 = io_dec_kill & inst_nback; // @[FetchInst.scala 67:25:@56.6]
  assign _T_169 = io_dec_kill == 1'h0; // @[FetchInst.scala 69:18:@61.8]
  assign _T_170 = _T_169 & inst_yback; // @[FetchInst.scala 69:31:@62.8]
  assign _T_172 = io_dec_forward == 1'h0; // @[FetchInst.scala 69:48:@63.8]
  assign _T_173 = _T_170 & _T_172; // @[FetchInst.scala 69:45:@64.8]
  assign _GEN_5 = _T_173 ? 2'h1 : inst_state; // @[FetchInst.scala 69:65:@65.8]
  assign _GEN_6 = _T_167 ? 2'h2 : _GEN_5; // @[FetchInst.scala 67:40:@57.6]
  assign _T_174 = 2'h1 == inst_state; // @[Conditional.scala 37:30:@70.6]
  assign _T_175 = io_dec_forward | io_dec_kill; // @[FetchInst.scala 74:28:@72.8]
  assign _GEN_7 = _T_175 ? 2'h0 : inst_state; // @[FetchInst.scala 74:44:@73.8]
  assign _T_176 = 2'h2 == inst_state; // @[Conditional.scala 37:30:@78.8]
  assign _GEN_8 = io_mem_resp_valid ? 2'h0 : inst_state; // @[FetchInst.scala 79:32:@80.10]
  assign _GEN_9 = _T_176 ? _GEN_8 : inst_state; // @[Conditional.scala 39:67:@79.8]
  assign _GEN_10 = _T_174 ? _GEN_7 : _GEN_9; // @[Conditional.scala 39:67:@71.6]
  assign _GEN_11 = _T_166 ? _GEN_6 : _GEN_10; // @[Conditional.scala 40:58:@55.4]
  assign _T_178 = inst_state == 2'h1; // @[FetchInst.scala 88:39:@88.4]
  assign _T_180 = inst_state == 2'h0; // @[FetchInst.scala 89:35:@91.4]
  assign _T_181 = _T_180 & inst_yback; // @[FetchInst.scala 89:45:@92.4]
  assign io_mem_req_valid = inst_nback == 1'h0; // @[FetchInst.scala 53:24:@44.4]
  assign io_mem_req_bits_addr = if_reg_pc; // @[FetchInst.scala 56:24:@49.4]
  assign io_if_forward = _T_161 & _T_151; // @[FetchInst.scala 55:24:@48.4]
  assign io_if_pc = if_reg_pc; // @[FetchInst.scala 25:13:@9.4]
  assign io_dec_inst_valid = _T_181 | _T_178; // @[FetchInst.scala 89:21:@95.4]
  assign io_dec_inst_bits = _T_178 ? reg_inst : io_mem_resp_bits_data; // @[FetchInst.scala 88:21:@90.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  if_reg_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pc_state = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  inst_state = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_inst = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      if_reg_pc <= 32'h80000000;
    end else begin
      if (_T_144) begin
        if (io_if_kill) begin
          if_reg_pc <= io_if_target;
        end else begin
          if_reg_pc <= io_btb_target;
        end
      end
    end
    if (reset) begin
      pc_state <= 1'h0;
    end else begin
      if (_T_156) begin
        if (pc_ready) begin
          pc_state <= 1'h1;
        end
      end else begin
        if (pc_state) begin
          if (io_mem_resp_valid) begin
            pc_state <= pc_ready;
          end
        end
      end
    end
    if (reset) begin
      inst_state <= 2'h0;
    end else begin
      if (_T_166) begin
        if (_T_167) begin
          inst_state <= 2'h2;
        end else begin
          if (_T_173) begin
            inst_state <= 2'h1;
          end
        end
      end else begin
        if (_T_174) begin
          if (_T_175) begin
            inst_state <= 2'h0;
          end
        end else begin
          if (_T_176) begin
            if (io_mem_resp_valid) begin
              inst_state <= 2'h0;
            end
          end
        end
      end
    end
    if (inst_yback) begin
      reg_inst <= io_mem_resp_bits_data;
    end
  end
endmodule
module BTB( // @[:@97.2]
  input         clock, // @[:@98.4]
  input         reset, // @[:@99.4]
  input  [31:0] io_if_pc, // @[:@100.4]
  input  [31:0] io_ras_peek, // @[:@100.4]
  output [31:0] io_pred_pc, // @[:@100.4]
  input  [31:0] io_fb_pc, // @[:@100.4]
  input  [1:0]  io_fb_type, // @[:@100.4]
  input         io_feedBack_valid, // @[:@100.4]
  input         io_feedBack_bits_redirect, // @[:@100.4]
  input  [31:0] io_feedBack_bits_tgt // @[:@100.4]
);
  reg [31:0] btb_pc_0; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_0;
  reg [31:0] btb_pc_1; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_1;
  reg [31:0] btb_pc_2; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_2;
  reg [31:0] btb_pc_3; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_3;
  reg [31:0] btb_pc_4; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_4;
  reg [31:0] btb_pc_5; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_5;
  reg [31:0] btb_pc_6; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_6;
  reg [31:0] btb_pc_7; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_7;
  reg [31:0] btb_pc_8; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_8;
  reg [31:0] btb_pc_9; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_9;
  reg [31:0] btb_pc_10; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_10;
  reg [31:0] btb_pc_11; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_11;
  reg [31:0] btb_pc_12; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_12;
  reg [31:0] btb_pc_13; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_13;
  reg [31:0] btb_pc_14; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_14;
  reg [31:0] btb_pc_15; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_15;
  reg [31:0] btb_pc_16; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_16;
  reg [31:0] btb_pc_17; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_17;
  reg [31:0] btb_pc_18; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_18;
  reg [31:0] btb_pc_19; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_19;
  reg [31:0] btb_pc_20; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_20;
  reg [31:0] btb_pc_21; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_21;
  reg [31:0] btb_pc_22; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_22;
  reg [31:0] btb_pc_23; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_23;
  reg [31:0] btb_pc_24; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_24;
  reg [31:0] btb_pc_25; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_25;
  reg [31:0] btb_pc_26; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_26;
  reg [31:0] btb_pc_27; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_27;
  reg [31:0] btb_pc_28; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_28;
  reg [31:0] btb_pc_29; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_29;
  reg [31:0] btb_pc_30; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_30;
  reg [31:0] btb_pc_31; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_31;
  reg [31:0] btb_pc_32; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_32;
  reg [31:0] btb_pc_33; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_33;
  reg [31:0] btb_pc_34; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_34;
  reg [31:0] btb_pc_35; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_35;
  reg [31:0] btb_pc_36; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_36;
  reg [31:0] btb_pc_37; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_37;
  reg [31:0] btb_pc_38; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_38;
  reg [31:0] btb_pc_39; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_39;
  reg [31:0] btb_pc_40; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_40;
  reg [31:0] btb_pc_41; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_41;
  reg [31:0] btb_pc_42; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_42;
  reg [31:0] btb_pc_43; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_43;
  reg [31:0] btb_pc_44; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_44;
  reg [31:0] btb_pc_45; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_45;
  reg [31:0] btb_pc_46; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_46;
  reg [31:0] btb_pc_47; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_47;
  reg [31:0] btb_pc_48; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_48;
  reg [31:0] btb_pc_49; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_49;
  reg [31:0] btb_pc_50; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_50;
  reg [31:0] btb_pc_51; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_51;
  reg [31:0] btb_pc_52; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_52;
  reg [31:0] btb_pc_53; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_53;
  reg [31:0] btb_pc_54; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_54;
  reg [31:0] btb_pc_55; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_55;
  reg [31:0] btb_pc_56; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_56;
  reg [31:0] btb_pc_57; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_57;
  reg [31:0] btb_pc_58; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_58;
  reg [31:0] btb_pc_59; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_59;
  reg [31:0] btb_pc_60; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_60;
  reg [31:0] btb_pc_61; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_61;
  reg [31:0] btb_pc_62; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_62;
  reg [31:0] btb_pc_63; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_63;
  reg [31:0] btb_target_0; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_64;
  reg [31:0] btb_target_1; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_65;
  reg [31:0] btb_target_2; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_66;
  reg [31:0] btb_target_3; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_67;
  reg [31:0] btb_target_4; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_68;
  reg [31:0] btb_target_5; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_69;
  reg [31:0] btb_target_6; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_70;
  reg [31:0] btb_target_7; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_71;
  reg [31:0] btb_target_8; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_72;
  reg [31:0] btb_target_9; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_73;
  reg [31:0] btb_target_10; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_74;
  reg [31:0] btb_target_11; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_75;
  reg [31:0] btb_target_12; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_76;
  reg [31:0] btb_target_13; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_77;
  reg [31:0] btb_target_14; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_78;
  reg [31:0] btb_target_15; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_79;
  reg [31:0] btb_target_16; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_80;
  reg [31:0] btb_target_17; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_81;
  reg [31:0] btb_target_18; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_82;
  reg [31:0] btb_target_19; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_83;
  reg [31:0] btb_target_20; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_84;
  reg [31:0] btb_target_21; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_85;
  reg [31:0] btb_target_22; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_86;
  reg [31:0] btb_target_23; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_87;
  reg [31:0] btb_target_24; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_88;
  reg [31:0] btb_target_25; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_89;
  reg [31:0] btb_target_26; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_90;
  reg [31:0] btb_target_27; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_91;
  reg [31:0] btb_target_28; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_92;
  reg [31:0] btb_target_29; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_93;
  reg [31:0] btb_target_30; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_94;
  reg [31:0] btb_target_31; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_95;
  reg [31:0] btb_target_32; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_96;
  reg [31:0] btb_target_33; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_97;
  reg [31:0] btb_target_34; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_98;
  reg [31:0] btb_target_35; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_99;
  reg [31:0] btb_target_36; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_100;
  reg [31:0] btb_target_37; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_101;
  reg [31:0] btb_target_38; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_102;
  reg [31:0] btb_target_39; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_103;
  reg [31:0] btb_target_40; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_104;
  reg [31:0] btb_target_41; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_105;
  reg [31:0] btb_target_42; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_106;
  reg [31:0] btb_target_43; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_107;
  reg [31:0] btb_target_44; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_108;
  reg [31:0] btb_target_45; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_109;
  reg [31:0] btb_target_46; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_110;
  reg [31:0] btb_target_47; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_111;
  reg [31:0] btb_target_48; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_112;
  reg [31:0] btb_target_49; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_113;
  reg [31:0] btb_target_50; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_114;
  reg [31:0] btb_target_51; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_115;
  reg [31:0] btb_target_52; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_116;
  reg [31:0] btb_target_53; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_117;
  reg [31:0] btb_target_54; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_118;
  reg [31:0] btb_target_55; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_119;
  reg [31:0] btb_target_56; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_120;
  reg [31:0] btb_target_57; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_121;
  reg [31:0] btb_target_58; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_122;
  reg [31:0] btb_target_59; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_123;
  reg [31:0] btb_target_60; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_124;
  reg [31:0] btb_target_61; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_125;
  reg [31:0] btb_target_62; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_126;
  reg [31:0] btb_target_63; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_127;
  reg [1:0] btb_hcount_0; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_128;
  reg [1:0] btb_hcount_1; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_129;
  reg [1:0] btb_hcount_2; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_130;
  reg [1:0] btb_hcount_3; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_131;
  reg [1:0] btb_hcount_4; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_132;
  reg [1:0] btb_hcount_5; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_133;
  reg [1:0] btb_hcount_6; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_134;
  reg [1:0] btb_hcount_7; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_135;
  reg [1:0] btb_hcount_8; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_136;
  reg [1:0] btb_hcount_9; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_137;
  reg [1:0] btb_hcount_10; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_138;
  reg [1:0] btb_hcount_11; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_139;
  reg [1:0] btb_hcount_12; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_140;
  reg [1:0] btb_hcount_13; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_141;
  reg [1:0] btb_hcount_14; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_142;
  reg [1:0] btb_hcount_15; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_143;
  reg [1:0] btb_hcount_16; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_144;
  reg [1:0] btb_hcount_17; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_145;
  reg [1:0] btb_hcount_18; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_146;
  reg [1:0] btb_hcount_19; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_147;
  reg [1:0] btb_hcount_20; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_148;
  reg [1:0] btb_hcount_21; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_149;
  reg [1:0] btb_hcount_22; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_150;
  reg [1:0] btb_hcount_23; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_151;
  reg [1:0] btb_hcount_24; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_152;
  reg [1:0] btb_hcount_25; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_153;
  reg [1:0] btb_hcount_26; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_154;
  reg [1:0] btb_hcount_27; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_155;
  reg [1:0] btb_hcount_28; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_156;
  reg [1:0] btb_hcount_29; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_157;
  reg [1:0] btb_hcount_30; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_158;
  reg [1:0] btb_hcount_31; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_159;
  reg [1:0] btb_hcount_32; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_160;
  reg [1:0] btb_hcount_33; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_161;
  reg [1:0] btb_hcount_34; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_162;
  reg [1:0] btb_hcount_35; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_163;
  reg [1:0] btb_hcount_36; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_164;
  reg [1:0] btb_hcount_37; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_165;
  reg [1:0] btb_hcount_38; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_166;
  reg [1:0] btb_hcount_39; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_167;
  reg [1:0] btb_hcount_40; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_168;
  reg [1:0] btb_hcount_41; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_169;
  reg [1:0] btb_hcount_42; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_170;
  reg [1:0] btb_hcount_43; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_171;
  reg [1:0] btb_hcount_44; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_172;
  reg [1:0] btb_hcount_45; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_173;
  reg [1:0] btb_hcount_46; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_174;
  reg [1:0] btb_hcount_47; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_175;
  reg [1:0] btb_hcount_48; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_176;
  reg [1:0] btb_hcount_49; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_177;
  reg [1:0] btb_hcount_50; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_178;
  reg [1:0] btb_hcount_51; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_179;
  reg [1:0] btb_hcount_52; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_180;
  reg [1:0] btb_hcount_53; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_181;
  reg [1:0] btb_hcount_54; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_182;
  reg [1:0] btb_hcount_55; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_183;
  reg [1:0] btb_hcount_56; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_184;
  reg [1:0] btb_hcount_57; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_185;
  reg [1:0] btb_hcount_58; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_186;
  reg [1:0] btb_hcount_59; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_187;
  reg [1:0] btb_hcount_60; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_188;
  reg [1:0] btb_hcount_61; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_189;
  reg [1:0] btb_hcount_62; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_190;
  reg [1:0] btb_hcount_63; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_191;
  reg [1:0] btb_btype_0; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_192;
  reg [1:0] btb_btype_1; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_193;
  reg [1:0] btb_btype_2; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_194;
  reg [1:0] btb_btype_3; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_195;
  reg [1:0] btb_btype_4; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_196;
  reg [1:0] btb_btype_5; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_197;
  reg [1:0] btb_btype_6; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_198;
  reg [1:0] btb_btype_7; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_199;
  reg [1:0] btb_btype_8; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_200;
  reg [1:0] btb_btype_9; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_201;
  reg [1:0] btb_btype_10; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_202;
  reg [1:0] btb_btype_11; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_203;
  reg [1:0] btb_btype_12; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_204;
  reg [1:0] btb_btype_13; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_205;
  reg [1:0] btb_btype_14; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_206;
  reg [1:0] btb_btype_15; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_207;
  reg [1:0] btb_btype_16; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_208;
  reg [1:0] btb_btype_17; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_209;
  reg [1:0] btb_btype_18; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_210;
  reg [1:0] btb_btype_19; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_211;
  reg [1:0] btb_btype_20; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_212;
  reg [1:0] btb_btype_21; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_213;
  reg [1:0] btb_btype_22; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_214;
  reg [1:0] btb_btype_23; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_215;
  reg [1:0] btb_btype_24; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_216;
  reg [1:0] btb_btype_25; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_217;
  reg [1:0] btb_btype_26; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_218;
  reg [1:0] btb_btype_27; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_219;
  reg [1:0] btb_btype_28; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_220;
  reg [1:0] btb_btype_29; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_221;
  reg [1:0] btb_btype_30; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_222;
  reg [1:0] btb_btype_31; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_223;
  reg [1:0] btb_btype_32; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_224;
  reg [1:0] btb_btype_33; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_225;
  reg [1:0] btb_btype_34; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_226;
  reg [1:0] btb_btype_35; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_227;
  reg [1:0] btb_btype_36; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_228;
  reg [1:0] btb_btype_37; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_229;
  reg [1:0] btb_btype_38; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_230;
  reg [1:0] btb_btype_39; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_231;
  reg [1:0] btb_btype_40; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_232;
  reg [1:0] btb_btype_41; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_233;
  reg [1:0] btb_btype_42; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_234;
  reg [1:0] btb_btype_43; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_235;
  reg [1:0] btb_btype_44; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_236;
  reg [1:0] btb_btype_45; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_237;
  reg [1:0] btb_btype_46; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_238;
  reg [1:0] btb_btype_47; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_239;
  reg [1:0] btb_btype_48; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_240;
  reg [1:0] btb_btype_49; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_241;
  reg [1:0] btb_btype_50; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_242;
  reg [1:0] btb_btype_51; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_243;
  reg [1:0] btb_btype_52; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_244;
  reg [1:0] btb_btype_53; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_245;
  reg [1:0] btb_btype_54; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_246;
  reg [1:0] btb_btype_55; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_247;
  reg [1:0] btb_btype_56; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_248;
  reg [1:0] btb_btype_57; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_249;
  reg [1:0] btb_btype_58; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_250;
  reg [1:0] btb_btype_59; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_251;
  reg [1:0] btb_btype_60; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_252;
  reg [1:0] btb_btype_61; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_253;
  reg [1:0] btb_btype_62; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_254;
  reg [1:0] btb_btype_63; // @[BTB.scala 44:20:@359.4]
  reg [31:0] _RAND_255;
  wire  _T_125; // @[BTB.scala 70:42:@361.4]
  wire  _T_126; // @[BTB.scala 70:42:@362.4]
  wire  _T_127; // @[BTB.scala 70:42:@363.4]
  wire  _T_128; // @[BTB.scala 70:42:@364.4]
  wire  _T_129; // @[BTB.scala 70:42:@365.4]
  wire  _T_130; // @[BTB.scala 70:42:@366.4]
  wire  _T_131; // @[BTB.scala 70:42:@367.4]
  wire  _T_132; // @[BTB.scala 70:42:@368.4]
  wire  _T_133; // @[BTB.scala 70:42:@369.4]
  wire  _T_134; // @[BTB.scala 70:42:@370.4]
  wire  _T_135; // @[BTB.scala 70:42:@371.4]
  wire  _T_136; // @[BTB.scala 70:42:@372.4]
  wire  _T_137; // @[BTB.scala 70:42:@373.4]
  wire  _T_138; // @[BTB.scala 70:42:@374.4]
  wire  _T_139; // @[BTB.scala 70:42:@375.4]
  wire  _T_140; // @[BTB.scala 70:42:@376.4]
  wire  _T_141; // @[BTB.scala 70:42:@377.4]
  wire  _T_142; // @[BTB.scala 70:42:@378.4]
  wire  _T_143; // @[BTB.scala 70:42:@379.4]
  wire  _T_144; // @[BTB.scala 70:42:@380.4]
  wire  _T_145; // @[BTB.scala 70:42:@381.4]
  wire  _T_146; // @[BTB.scala 70:42:@382.4]
  wire  _T_147; // @[BTB.scala 70:42:@383.4]
  wire  _T_148; // @[BTB.scala 70:42:@384.4]
  wire  _T_149; // @[BTB.scala 70:42:@385.4]
  wire  _T_150; // @[BTB.scala 70:42:@386.4]
  wire  _T_151; // @[BTB.scala 70:42:@387.4]
  wire  _T_152; // @[BTB.scala 70:42:@388.4]
  wire  _T_153; // @[BTB.scala 70:42:@389.4]
  wire  _T_154; // @[BTB.scala 70:42:@390.4]
  wire  _T_155; // @[BTB.scala 70:42:@391.4]
  wire  _T_156; // @[BTB.scala 70:42:@392.4]
  wire  _T_157; // @[BTB.scala 70:42:@393.4]
  wire  _T_158; // @[BTB.scala 70:42:@394.4]
  wire  _T_159; // @[BTB.scala 70:42:@395.4]
  wire  _T_160; // @[BTB.scala 70:42:@396.4]
  wire  _T_161; // @[BTB.scala 70:42:@397.4]
  wire  _T_162; // @[BTB.scala 70:42:@398.4]
  wire  _T_163; // @[BTB.scala 70:42:@399.4]
  wire  _T_164; // @[BTB.scala 70:42:@400.4]
  wire  _T_165; // @[BTB.scala 70:42:@401.4]
  wire  _T_166; // @[BTB.scala 70:42:@402.4]
  wire  _T_167; // @[BTB.scala 70:42:@403.4]
  wire  _T_168; // @[BTB.scala 70:42:@404.4]
  wire  _T_169; // @[BTB.scala 70:42:@405.4]
  wire  _T_170; // @[BTB.scala 70:42:@406.4]
  wire  _T_171; // @[BTB.scala 70:42:@407.4]
  wire  _T_172; // @[BTB.scala 70:42:@408.4]
  wire  _T_173; // @[BTB.scala 70:42:@409.4]
  wire  _T_174; // @[BTB.scala 70:42:@410.4]
  wire  _T_175; // @[BTB.scala 70:42:@411.4]
  wire  _T_176; // @[BTB.scala 70:42:@412.4]
  wire  _T_177; // @[BTB.scala 70:42:@413.4]
  wire  _T_178; // @[BTB.scala 70:42:@414.4]
  wire  _T_179; // @[BTB.scala 70:42:@415.4]
  wire  _T_180; // @[BTB.scala 70:42:@416.4]
  wire  _T_181; // @[BTB.scala 70:42:@417.4]
  wire  _T_182; // @[BTB.scala 70:42:@418.4]
  wire  _T_183; // @[BTB.scala 70:42:@419.4]
  wire  _T_184; // @[BTB.scala 70:42:@420.4]
  wire  _T_185; // @[BTB.scala 70:42:@421.4]
  wire  _T_186; // @[BTB.scala 70:42:@422.4]
  wire  _T_187; // @[BTB.scala 70:42:@423.4]
  wire  _T_188; // @[BTB.scala 70:42:@424.4]
  wire [7:0] _T_265; // @[BTB.scala 70:57:@496.4]
  wire [15:0] _T_273; // @[BTB.scala 70:57:@504.4]
  wire [7:0] _T_280; // @[BTB.scala 70:57:@511.4]
  wire [31:0] _T_289; // @[BTB.scala 70:57:@520.4]
  wire [7:0] _T_296; // @[BTB.scala 70:57:@527.4]
  wire [15:0] _T_304; // @[BTB.scala 70:57:@535.4]
  wire [7:0] _T_311; // @[BTB.scala 70:57:@542.4]
  wire [31:0] _T_320; // @[BTB.scala 70:57:@551.4]
  wire [63:0] _T_321; // @[BTB.scala 70:57:@552.4]
  wire  _T_323; // @[BTB.scala 50:66:@553.4]
  wire  _T_325; // @[BTB.scala 50:66:@554.4]
  wire  _T_327; // @[BTB.scala 50:66:@555.4]
  wire  _T_329; // @[BTB.scala 50:66:@556.4]
  wire  _T_331; // @[BTB.scala 50:66:@557.4]
  wire  _T_333; // @[BTB.scala 50:66:@558.4]
  wire  _T_335; // @[BTB.scala 50:66:@559.4]
  wire  _T_337; // @[BTB.scala 50:66:@560.4]
  wire  _T_339; // @[BTB.scala 50:66:@561.4]
  wire  _T_341; // @[BTB.scala 50:66:@562.4]
  wire  _T_343; // @[BTB.scala 50:66:@563.4]
  wire  _T_345; // @[BTB.scala 50:66:@564.4]
  wire  _T_347; // @[BTB.scala 50:66:@565.4]
  wire  _T_349; // @[BTB.scala 50:66:@566.4]
  wire  _T_351; // @[BTB.scala 50:66:@567.4]
  wire  _T_353; // @[BTB.scala 50:66:@568.4]
  wire  _T_355; // @[BTB.scala 50:66:@569.4]
  wire  _T_357; // @[BTB.scala 50:66:@570.4]
  wire  _T_359; // @[BTB.scala 50:66:@571.4]
  wire  _T_361; // @[BTB.scala 50:66:@572.4]
  wire  _T_363; // @[BTB.scala 50:66:@573.4]
  wire  _T_365; // @[BTB.scala 50:66:@574.4]
  wire  _T_367; // @[BTB.scala 50:66:@575.4]
  wire  _T_369; // @[BTB.scala 50:66:@576.4]
  wire  _T_371; // @[BTB.scala 50:66:@577.4]
  wire  _T_373; // @[BTB.scala 50:66:@578.4]
  wire  _T_375; // @[BTB.scala 50:66:@579.4]
  wire  _T_377; // @[BTB.scala 50:66:@580.4]
  wire  _T_379; // @[BTB.scala 50:66:@581.4]
  wire  _T_381; // @[BTB.scala 50:66:@582.4]
  wire  _T_383; // @[BTB.scala 50:66:@583.4]
  wire  _T_385; // @[BTB.scala 50:66:@584.4]
  wire  _T_387; // @[BTB.scala 50:66:@585.4]
  wire  _T_389; // @[BTB.scala 50:66:@586.4]
  wire  _T_391; // @[BTB.scala 50:66:@587.4]
  wire  _T_393; // @[BTB.scala 50:66:@588.4]
  wire  _T_395; // @[BTB.scala 50:66:@589.4]
  wire  _T_397; // @[BTB.scala 50:66:@590.4]
  wire  _T_399; // @[BTB.scala 50:66:@591.4]
  wire  _T_401; // @[BTB.scala 50:66:@592.4]
  wire  _T_403; // @[BTB.scala 50:66:@593.4]
  wire  _T_405; // @[BTB.scala 50:66:@594.4]
  wire  _T_407; // @[BTB.scala 50:66:@595.4]
  wire  _T_409; // @[BTB.scala 50:66:@596.4]
  wire  _T_411; // @[BTB.scala 50:66:@597.4]
  wire  _T_413; // @[BTB.scala 50:66:@598.4]
  wire  _T_415; // @[BTB.scala 50:66:@599.4]
  wire  _T_417; // @[BTB.scala 50:66:@600.4]
  wire  _T_419; // @[BTB.scala 50:66:@601.4]
  wire  _T_421; // @[BTB.scala 50:66:@602.4]
  wire  _T_423; // @[BTB.scala 50:66:@603.4]
  wire  _T_425; // @[BTB.scala 50:66:@604.4]
  wire  _T_427; // @[BTB.scala 50:66:@605.4]
  wire  _T_429; // @[BTB.scala 50:66:@606.4]
  wire  _T_431; // @[BTB.scala 50:66:@607.4]
  wire  _T_433; // @[BTB.scala 50:66:@608.4]
  wire  _T_435; // @[BTB.scala 50:66:@609.4]
  wire  _T_437; // @[BTB.scala 50:66:@610.4]
  wire  _T_439; // @[BTB.scala 50:66:@611.4]
  wire  _T_441; // @[BTB.scala 50:66:@612.4]
  wire  _T_443; // @[BTB.scala 50:66:@613.4]
  wire  _T_445; // @[BTB.scala 50:66:@614.4]
  wire  _T_447; // @[BTB.scala 50:66:@615.4]
  wire  _T_449; // @[BTB.scala 50:66:@616.4]
  wire [7:0] _T_526; // @[BTB.scala 50:72:@688.4]
  wire [15:0] _T_534; // @[BTB.scala 50:72:@696.4]
  wire [7:0] _T_541; // @[BTB.scala 50:72:@703.4]
  wire [31:0] _T_550; // @[BTB.scala 50:72:@712.4]
  wire [7:0] _T_557; // @[BTB.scala 50:72:@719.4]
  wire [15:0] _T_565; // @[BTB.scala 50:72:@727.4]
  wire [7:0] _T_572; // @[BTB.scala 50:72:@734.4]
  wire [31:0] _T_581; // @[BTB.scala 50:72:@743.4]
  wire [63:0] _T_582; // @[BTB.scala 50:72:@744.4]
  wire [63:0] predict_lookup; // @[BTB.scala 70:64:@745.4]
  wire [32:0] _T_585; // @[BTB.scala 71:32:@747.4]
  wire [31:0] predict_cont_tgt; // @[BTB.scala 71:32:@748.4]
  wire  _T_587; // @[Mux.scala 21:36:@750.4]
  wire  _T_588; // @[Mux.scala 21:36:@751.4]
  wire  _T_589; // @[Mux.scala 21:36:@752.4]
  wire  _T_590; // @[Mux.scala 21:36:@753.4]
  wire  _T_591; // @[Mux.scala 21:36:@754.4]
  wire  _T_592; // @[Mux.scala 21:36:@755.4]
  wire  _T_593; // @[Mux.scala 21:36:@756.4]
  wire  _T_594; // @[Mux.scala 21:36:@757.4]
  wire  _T_595; // @[Mux.scala 21:36:@758.4]
  wire  _T_596; // @[Mux.scala 21:36:@759.4]
  wire  _T_597; // @[Mux.scala 21:36:@760.4]
  wire  _T_598; // @[Mux.scala 21:36:@761.4]
  wire  _T_599; // @[Mux.scala 21:36:@762.4]
  wire  _T_600; // @[Mux.scala 21:36:@763.4]
  wire  _T_601; // @[Mux.scala 21:36:@764.4]
  wire  _T_602; // @[Mux.scala 21:36:@765.4]
  wire  _T_603; // @[Mux.scala 21:36:@766.4]
  wire  _T_604; // @[Mux.scala 21:36:@767.4]
  wire  _T_605; // @[Mux.scala 21:36:@768.4]
  wire  _T_606; // @[Mux.scala 21:36:@769.4]
  wire  _T_607; // @[Mux.scala 21:36:@770.4]
  wire  _T_608; // @[Mux.scala 21:36:@771.4]
  wire  _T_609; // @[Mux.scala 21:36:@772.4]
  wire  _T_610; // @[Mux.scala 21:36:@773.4]
  wire  _T_611; // @[Mux.scala 21:36:@774.4]
  wire  _T_612; // @[Mux.scala 21:36:@775.4]
  wire  _T_613; // @[Mux.scala 21:36:@776.4]
  wire  _T_614; // @[Mux.scala 21:36:@777.4]
  wire  _T_615; // @[Mux.scala 21:36:@778.4]
  wire  _T_616; // @[Mux.scala 21:36:@779.4]
  wire  _T_617; // @[Mux.scala 21:36:@780.4]
  wire  _T_618; // @[Mux.scala 21:36:@781.4]
  wire  _T_619; // @[Mux.scala 21:36:@782.4]
  wire  _T_620; // @[Mux.scala 21:36:@783.4]
  wire  _T_621; // @[Mux.scala 21:36:@784.4]
  wire  _T_622; // @[Mux.scala 21:36:@785.4]
  wire  _T_623; // @[Mux.scala 21:36:@786.4]
  wire  _T_624; // @[Mux.scala 21:36:@787.4]
  wire  _T_625; // @[Mux.scala 21:36:@788.4]
  wire  _T_626; // @[Mux.scala 21:36:@789.4]
  wire  _T_627; // @[Mux.scala 21:36:@790.4]
  wire  _T_628; // @[Mux.scala 21:36:@791.4]
  wire  _T_629; // @[Mux.scala 21:36:@792.4]
  wire  _T_630; // @[Mux.scala 21:36:@793.4]
  wire  _T_631; // @[Mux.scala 21:36:@794.4]
  wire  _T_632; // @[Mux.scala 21:36:@795.4]
  wire  _T_633; // @[Mux.scala 21:36:@796.4]
  wire  _T_634; // @[Mux.scala 21:36:@797.4]
  wire  _T_635; // @[Mux.scala 21:36:@798.4]
  wire  _T_636; // @[Mux.scala 21:36:@799.4]
  wire  _T_637; // @[Mux.scala 21:36:@800.4]
  wire  _T_638; // @[Mux.scala 21:36:@801.4]
  wire  _T_639; // @[Mux.scala 21:36:@802.4]
  wire  _T_640; // @[Mux.scala 21:36:@803.4]
  wire  _T_641; // @[Mux.scala 21:36:@804.4]
  wire  _T_642; // @[Mux.scala 21:36:@805.4]
  wire  _T_643; // @[Mux.scala 21:36:@806.4]
  wire  _T_644; // @[Mux.scala 21:36:@807.4]
  wire  _T_645; // @[Mux.scala 21:36:@808.4]
  wire  _T_646; // @[Mux.scala 21:36:@809.4]
  wire  _T_647; // @[Mux.scala 21:36:@810.4]
  wire  _T_648; // @[Mux.scala 21:36:@811.4]
  wire  _T_649; // @[Mux.scala 21:36:@812.4]
  wire  _T_650; // @[Mux.scala 21:36:@813.4]
  wire [31:0] _T_653; // @[Mux.scala 19:72:@814.4]
  wire [31:0] _T_655; // @[Mux.scala 19:72:@815.4]
  wire [31:0] _T_657; // @[Mux.scala 19:72:@816.4]
  wire [31:0] _T_659; // @[Mux.scala 19:72:@817.4]
  wire [31:0] _T_661; // @[Mux.scala 19:72:@818.4]
  wire [31:0] _T_663; // @[Mux.scala 19:72:@819.4]
  wire [31:0] _T_665; // @[Mux.scala 19:72:@820.4]
  wire [31:0] _T_667; // @[Mux.scala 19:72:@821.4]
  wire [31:0] _T_669; // @[Mux.scala 19:72:@822.4]
  wire [31:0] _T_671; // @[Mux.scala 19:72:@823.4]
  wire [31:0] _T_673; // @[Mux.scala 19:72:@824.4]
  wire [31:0] _T_675; // @[Mux.scala 19:72:@825.4]
  wire [31:0] _T_677; // @[Mux.scala 19:72:@826.4]
  wire [31:0] _T_679; // @[Mux.scala 19:72:@827.4]
  wire [31:0] _T_681; // @[Mux.scala 19:72:@828.4]
  wire [31:0] _T_683; // @[Mux.scala 19:72:@829.4]
  wire [31:0] _T_685; // @[Mux.scala 19:72:@830.4]
  wire [31:0] _T_687; // @[Mux.scala 19:72:@831.4]
  wire [31:0] _T_689; // @[Mux.scala 19:72:@832.4]
  wire [31:0] _T_691; // @[Mux.scala 19:72:@833.4]
  wire [31:0] _T_693; // @[Mux.scala 19:72:@834.4]
  wire [31:0] _T_695; // @[Mux.scala 19:72:@835.4]
  wire [31:0] _T_697; // @[Mux.scala 19:72:@836.4]
  wire [31:0] _T_699; // @[Mux.scala 19:72:@837.4]
  wire [31:0] _T_701; // @[Mux.scala 19:72:@838.4]
  wire [31:0] _T_703; // @[Mux.scala 19:72:@839.4]
  wire [31:0] _T_705; // @[Mux.scala 19:72:@840.4]
  wire [31:0] _T_707; // @[Mux.scala 19:72:@841.4]
  wire [31:0] _T_709; // @[Mux.scala 19:72:@842.4]
  wire [31:0] _T_711; // @[Mux.scala 19:72:@843.4]
  wire [31:0] _T_713; // @[Mux.scala 19:72:@844.4]
  wire [31:0] _T_715; // @[Mux.scala 19:72:@845.4]
  wire [31:0] _T_717; // @[Mux.scala 19:72:@846.4]
  wire [31:0] _T_719; // @[Mux.scala 19:72:@847.4]
  wire [31:0] _T_721; // @[Mux.scala 19:72:@848.4]
  wire [31:0] _T_723; // @[Mux.scala 19:72:@849.4]
  wire [31:0] _T_725; // @[Mux.scala 19:72:@850.4]
  wire [31:0] _T_727; // @[Mux.scala 19:72:@851.4]
  wire [31:0] _T_729; // @[Mux.scala 19:72:@852.4]
  wire [31:0] _T_731; // @[Mux.scala 19:72:@853.4]
  wire [31:0] _T_733; // @[Mux.scala 19:72:@854.4]
  wire [31:0] _T_735; // @[Mux.scala 19:72:@855.4]
  wire [31:0] _T_737; // @[Mux.scala 19:72:@856.4]
  wire [31:0] _T_739; // @[Mux.scala 19:72:@857.4]
  wire [31:0] _T_741; // @[Mux.scala 19:72:@858.4]
  wire [31:0] _T_743; // @[Mux.scala 19:72:@859.4]
  wire [31:0] _T_745; // @[Mux.scala 19:72:@860.4]
  wire [31:0] _T_747; // @[Mux.scala 19:72:@861.4]
  wire [31:0] _T_749; // @[Mux.scala 19:72:@862.4]
  wire [31:0] _T_751; // @[Mux.scala 19:72:@863.4]
  wire [31:0] _T_753; // @[Mux.scala 19:72:@864.4]
  wire [31:0] _T_755; // @[Mux.scala 19:72:@865.4]
  wire [31:0] _T_757; // @[Mux.scala 19:72:@866.4]
  wire [31:0] _T_759; // @[Mux.scala 19:72:@867.4]
  wire [31:0] _T_761; // @[Mux.scala 19:72:@868.4]
  wire [31:0] _T_763; // @[Mux.scala 19:72:@869.4]
  wire [31:0] _T_765; // @[Mux.scala 19:72:@870.4]
  wire [31:0] _T_767; // @[Mux.scala 19:72:@871.4]
  wire [31:0] _T_769; // @[Mux.scala 19:72:@872.4]
  wire [31:0] _T_771; // @[Mux.scala 19:72:@873.4]
  wire [31:0] _T_773; // @[Mux.scala 19:72:@874.4]
  wire [31:0] _T_775; // @[Mux.scala 19:72:@875.4]
  wire [31:0] _T_777; // @[Mux.scala 19:72:@876.4]
  wire [31:0] _T_779; // @[Mux.scala 19:72:@877.4]
  wire [31:0] _T_780; // @[Mux.scala 19:72:@878.4]
  wire [31:0] _T_781; // @[Mux.scala 19:72:@879.4]
  wire [31:0] _T_782; // @[Mux.scala 19:72:@880.4]
  wire [31:0] _T_783; // @[Mux.scala 19:72:@881.4]
  wire [31:0] _T_784; // @[Mux.scala 19:72:@882.4]
  wire [31:0] _T_785; // @[Mux.scala 19:72:@883.4]
  wire [31:0] _T_786; // @[Mux.scala 19:72:@884.4]
  wire [31:0] _T_787; // @[Mux.scala 19:72:@885.4]
  wire [31:0] _T_788; // @[Mux.scala 19:72:@886.4]
  wire [31:0] _T_789; // @[Mux.scala 19:72:@887.4]
  wire [31:0] _T_790; // @[Mux.scala 19:72:@888.4]
  wire [31:0] _T_791; // @[Mux.scala 19:72:@889.4]
  wire [31:0] _T_792; // @[Mux.scala 19:72:@890.4]
  wire [31:0] _T_793; // @[Mux.scala 19:72:@891.4]
  wire [31:0] _T_794; // @[Mux.scala 19:72:@892.4]
  wire [31:0] _T_795; // @[Mux.scala 19:72:@893.4]
  wire [31:0] _T_796; // @[Mux.scala 19:72:@894.4]
  wire [31:0] _T_797; // @[Mux.scala 19:72:@895.4]
  wire [31:0] _T_798; // @[Mux.scala 19:72:@896.4]
  wire [31:0] _T_799; // @[Mux.scala 19:72:@897.4]
  wire [31:0] _T_800; // @[Mux.scala 19:72:@898.4]
  wire [31:0] _T_801; // @[Mux.scala 19:72:@899.4]
  wire [31:0] _T_802; // @[Mux.scala 19:72:@900.4]
  wire [31:0] _T_803; // @[Mux.scala 19:72:@901.4]
  wire [31:0] _T_804; // @[Mux.scala 19:72:@902.4]
  wire [31:0] _T_805; // @[Mux.scala 19:72:@903.4]
  wire [31:0] _T_806; // @[Mux.scala 19:72:@904.4]
  wire [31:0] _T_807; // @[Mux.scala 19:72:@905.4]
  wire [31:0] _T_808; // @[Mux.scala 19:72:@906.4]
  wire [31:0] _T_809; // @[Mux.scala 19:72:@907.4]
  wire [31:0] _T_810; // @[Mux.scala 19:72:@908.4]
  wire [31:0] _T_811; // @[Mux.scala 19:72:@909.4]
  wire [31:0] _T_812; // @[Mux.scala 19:72:@910.4]
  wire [31:0] _T_813; // @[Mux.scala 19:72:@911.4]
  wire [31:0] _T_814; // @[Mux.scala 19:72:@912.4]
  wire [31:0] _T_815; // @[Mux.scala 19:72:@913.4]
  wire [31:0] _T_816; // @[Mux.scala 19:72:@914.4]
  wire [31:0] _T_817; // @[Mux.scala 19:72:@915.4]
  wire [31:0] _T_818; // @[Mux.scala 19:72:@916.4]
  wire [31:0] _T_819; // @[Mux.scala 19:72:@917.4]
  wire [31:0] _T_820; // @[Mux.scala 19:72:@918.4]
  wire [31:0] _T_821; // @[Mux.scala 19:72:@919.4]
  wire [31:0] _T_822; // @[Mux.scala 19:72:@920.4]
  wire [31:0] _T_823; // @[Mux.scala 19:72:@921.4]
  wire [31:0] _T_824; // @[Mux.scala 19:72:@922.4]
  wire [31:0] _T_825; // @[Mux.scala 19:72:@923.4]
  wire [31:0] _T_826; // @[Mux.scala 19:72:@924.4]
  wire [31:0] _T_827; // @[Mux.scala 19:72:@925.4]
  wire [31:0] _T_828; // @[Mux.scala 19:72:@926.4]
  wire [31:0] _T_829; // @[Mux.scala 19:72:@927.4]
  wire [31:0] _T_830; // @[Mux.scala 19:72:@928.4]
  wire [31:0] _T_831; // @[Mux.scala 19:72:@929.4]
  wire [31:0] _T_832; // @[Mux.scala 19:72:@930.4]
  wire [31:0] _T_833; // @[Mux.scala 19:72:@931.4]
  wire [31:0] _T_834; // @[Mux.scala 19:72:@932.4]
  wire [31:0] _T_835; // @[Mux.scala 19:72:@933.4]
  wire [31:0] _T_836; // @[Mux.scala 19:72:@934.4]
  wire [31:0] _T_837; // @[Mux.scala 19:72:@935.4]
  wire [31:0] _T_838; // @[Mux.scala 19:72:@936.4]
  wire [31:0] _T_839; // @[Mux.scala 19:72:@937.4]
  wire [31:0] _T_840; // @[Mux.scala 19:72:@938.4]
  wire [31:0] _T_841; // @[Mux.scala 19:72:@939.4]
  wire [31:0] predict_jump_tgt; // @[Mux.scala 19:72:@940.4]
  wire [1:0] _T_911; // @[Mux.scala 19:72:@1008.4]
  wire [1:0] _T_913; // @[Mux.scala 19:72:@1009.4]
  wire [1:0] _T_915; // @[Mux.scala 19:72:@1010.4]
  wire [1:0] _T_917; // @[Mux.scala 19:72:@1011.4]
  wire [1:0] _T_919; // @[Mux.scala 19:72:@1012.4]
  wire [1:0] _T_921; // @[Mux.scala 19:72:@1013.4]
  wire [1:0] _T_923; // @[Mux.scala 19:72:@1014.4]
  wire [1:0] _T_925; // @[Mux.scala 19:72:@1015.4]
  wire [1:0] _T_927; // @[Mux.scala 19:72:@1016.4]
  wire [1:0] _T_929; // @[Mux.scala 19:72:@1017.4]
  wire [1:0] _T_931; // @[Mux.scala 19:72:@1018.4]
  wire [1:0] _T_933; // @[Mux.scala 19:72:@1019.4]
  wire [1:0] _T_935; // @[Mux.scala 19:72:@1020.4]
  wire [1:0] _T_937; // @[Mux.scala 19:72:@1021.4]
  wire [1:0] _T_939; // @[Mux.scala 19:72:@1022.4]
  wire [1:0] _T_941; // @[Mux.scala 19:72:@1023.4]
  wire [1:0] _T_943; // @[Mux.scala 19:72:@1024.4]
  wire [1:0] _T_945; // @[Mux.scala 19:72:@1025.4]
  wire [1:0] _T_947; // @[Mux.scala 19:72:@1026.4]
  wire [1:0] _T_949; // @[Mux.scala 19:72:@1027.4]
  wire [1:0] _T_951; // @[Mux.scala 19:72:@1028.4]
  wire [1:0] _T_953; // @[Mux.scala 19:72:@1029.4]
  wire [1:0] _T_955; // @[Mux.scala 19:72:@1030.4]
  wire [1:0] _T_957; // @[Mux.scala 19:72:@1031.4]
  wire [1:0] _T_959; // @[Mux.scala 19:72:@1032.4]
  wire [1:0] _T_961; // @[Mux.scala 19:72:@1033.4]
  wire [1:0] _T_963; // @[Mux.scala 19:72:@1034.4]
  wire [1:0] _T_965; // @[Mux.scala 19:72:@1035.4]
  wire [1:0] _T_967; // @[Mux.scala 19:72:@1036.4]
  wire [1:0] _T_969; // @[Mux.scala 19:72:@1037.4]
  wire [1:0] _T_971; // @[Mux.scala 19:72:@1038.4]
  wire [1:0] _T_973; // @[Mux.scala 19:72:@1039.4]
  wire [1:0] _T_975; // @[Mux.scala 19:72:@1040.4]
  wire [1:0] _T_977; // @[Mux.scala 19:72:@1041.4]
  wire [1:0] _T_979; // @[Mux.scala 19:72:@1042.4]
  wire [1:0] _T_981; // @[Mux.scala 19:72:@1043.4]
  wire [1:0] _T_983; // @[Mux.scala 19:72:@1044.4]
  wire [1:0] _T_985; // @[Mux.scala 19:72:@1045.4]
  wire [1:0] _T_987; // @[Mux.scala 19:72:@1046.4]
  wire [1:0] _T_989; // @[Mux.scala 19:72:@1047.4]
  wire [1:0] _T_991; // @[Mux.scala 19:72:@1048.4]
  wire [1:0] _T_993; // @[Mux.scala 19:72:@1049.4]
  wire [1:0] _T_995; // @[Mux.scala 19:72:@1050.4]
  wire [1:0] _T_997; // @[Mux.scala 19:72:@1051.4]
  wire [1:0] _T_999; // @[Mux.scala 19:72:@1052.4]
  wire [1:0] _T_1001; // @[Mux.scala 19:72:@1053.4]
  wire [1:0] _T_1003; // @[Mux.scala 19:72:@1054.4]
  wire [1:0] _T_1005; // @[Mux.scala 19:72:@1055.4]
  wire [1:0] _T_1007; // @[Mux.scala 19:72:@1056.4]
  wire [1:0] _T_1009; // @[Mux.scala 19:72:@1057.4]
  wire [1:0] _T_1011; // @[Mux.scala 19:72:@1058.4]
  wire [1:0] _T_1013; // @[Mux.scala 19:72:@1059.4]
  wire [1:0] _T_1015; // @[Mux.scala 19:72:@1060.4]
  wire [1:0] _T_1017; // @[Mux.scala 19:72:@1061.4]
  wire [1:0] _T_1019; // @[Mux.scala 19:72:@1062.4]
  wire [1:0] _T_1021; // @[Mux.scala 19:72:@1063.4]
  wire [1:0] _T_1023; // @[Mux.scala 19:72:@1064.4]
  wire [1:0] _T_1025; // @[Mux.scala 19:72:@1065.4]
  wire [1:0] _T_1027; // @[Mux.scala 19:72:@1066.4]
  wire [1:0] _T_1029; // @[Mux.scala 19:72:@1067.4]
  wire [1:0] _T_1031; // @[Mux.scala 19:72:@1068.4]
  wire [1:0] _T_1033; // @[Mux.scala 19:72:@1069.4]
  wire [1:0] _T_1035; // @[Mux.scala 19:72:@1070.4]
  wire [1:0] _T_1037; // @[Mux.scala 19:72:@1071.4]
  wire [1:0] _T_1038; // @[Mux.scala 19:72:@1072.4]
  wire [1:0] _T_1039; // @[Mux.scala 19:72:@1073.4]
  wire [1:0] _T_1040; // @[Mux.scala 19:72:@1074.4]
  wire [1:0] _T_1041; // @[Mux.scala 19:72:@1075.4]
  wire [1:0] _T_1042; // @[Mux.scala 19:72:@1076.4]
  wire [1:0] _T_1043; // @[Mux.scala 19:72:@1077.4]
  wire [1:0] _T_1044; // @[Mux.scala 19:72:@1078.4]
  wire [1:0] _T_1045; // @[Mux.scala 19:72:@1079.4]
  wire [1:0] _T_1046; // @[Mux.scala 19:72:@1080.4]
  wire [1:0] _T_1047; // @[Mux.scala 19:72:@1081.4]
  wire [1:0] _T_1048; // @[Mux.scala 19:72:@1082.4]
  wire [1:0] _T_1049; // @[Mux.scala 19:72:@1083.4]
  wire [1:0] _T_1050; // @[Mux.scala 19:72:@1084.4]
  wire [1:0] _T_1051; // @[Mux.scala 19:72:@1085.4]
  wire [1:0] _T_1052; // @[Mux.scala 19:72:@1086.4]
  wire [1:0] _T_1053; // @[Mux.scala 19:72:@1087.4]
  wire [1:0] _T_1054; // @[Mux.scala 19:72:@1088.4]
  wire [1:0] _T_1055; // @[Mux.scala 19:72:@1089.4]
  wire [1:0] _T_1056; // @[Mux.scala 19:72:@1090.4]
  wire [1:0] _T_1057; // @[Mux.scala 19:72:@1091.4]
  wire [1:0] _T_1058; // @[Mux.scala 19:72:@1092.4]
  wire [1:0] _T_1059; // @[Mux.scala 19:72:@1093.4]
  wire [1:0] _T_1060; // @[Mux.scala 19:72:@1094.4]
  wire [1:0] _T_1061; // @[Mux.scala 19:72:@1095.4]
  wire [1:0] _T_1062; // @[Mux.scala 19:72:@1096.4]
  wire [1:0] _T_1063; // @[Mux.scala 19:72:@1097.4]
  wire [1:0] _T_1064; // @[Mux.scala 19:72:@1098.4]
  wire [1:0] _T_1065; // @[Mux.scala 19:72:@1099.4]
  wire [1:0] _T_1066; // @[Mux.scala 19:72:@1100.4]
  wire [1:0] _T_1067; // @[Mux.scala 19:72:@1101.4]
  wire [1:0] _T_1068; // @[Mux.scala 19:72:@1102.4]
  wire [1:0] _T_1069; // @[Mux.scala 19:72:@1103.4]
  wire [1:0] _T_1070; // @[Mux.scala 19:72:@1104.4]
  wire [1:0] _T_1071; // @[Mux.scala 19:72:@1105.4]
  wire [1:0] _T_1072; // @[Mux.scala 19:72:@1106.4]
  wire [1:0] _T_1073; // @[Mux.scala 19:72:@1107.4]
  wire [1:0] _T_1074; // @[Mux.scala 19:72:@1108.4]
  wire [1:0] _T_1075; // @[Mux.scala 19:72:@1109.4]
  wire [1:0] _T_1076; // @[Mux.scala 19:72:@1110.4]
  wire [1:0] _T_1077; // @[Mux.scala 19:72:@1111.4]
  wire [1:0] _T_1078; // @[Mux.scala 19:72:@1112.4]
  wire [1:0] _T_1079; // @[Mux.scala 19:72:@1113.4]
  wire [1:0] _T_1080; // @[Mux.scala 19:72:@1114.4]
  wire [1:0] _T_1081; // @[Mux.scala 19:72:@1115.4]
  wire [1:0] _T_1082; // @[Mux.scala 19:72:@1116.4]
  wire [1:0] _T_1083; // @[Mux.scala 19:72:@1117.4]
  wire [1:0] _T_1084; // @[Mux.scala 19:72:@1118.4]
  wire [1:0] _T_1085; // @[Mux.scala 19:72:@1119.4]
  wire [1:0] _T_1086; // @[Mux.scala 19:72:@1120.4]
  wire [1:0] _T_1087; // @[Mux.scala 19:72:@1121.4]
  wire [1:0] _T_1088; // @[Mux.scala 19:72:@1122.4]
  wire [1:0] _T_1089; // @[Mux.scala 19:72:@1123.4]
  wire [1:0] _T_1090; // @[Mux.scala 19:72:@1124.4]
  wire [1:0] _T_1091; // @[Mux.scala 19:72:@1125.4]
  wire [1:0] _T_1092; // @[Mux.scala 19:72:@1126.4]
  wire [1:0] _T_1093; // @[Mux.scala 19:72:@1127.4]
  wire [1:0] _T_1094; // @[Mux.scala 19:72:@1128.4]
  wire [1:0] _T_1095; // @[Mux.scala 19:72:@1129.4]
  wire [1:0] _T_1096; // @[Mux.scala 19:72:@1130.4]
  wire [1:0] _T_1097; // @[Mux.scala 19:72:@1131.4]
  wire [1:0] _T_1098; // @[Mux.scala 19:72:@1132.4]
  wire [1:0] _T_1099; // @[Mux.scala 19:72:@1133.4]
  wire [1:0] predict_btype; // @[Mux.scala 19:72:@1134.4]
  wire [1:0] _T_1169; // @[Mux.scala 19:72:@1202.4]
  wire [1:0] _T_1171; // @[Mux.scala 19:72:@1203.4]
  wire [1:0] _T_1173; // @[Mux.scala 19:72:@1204.4]
  wire [1:0] _T_1175; // @[Mux.scala 19:72:@1205.4]
  wire [1:0] _T_1177; // @[Mux.scala 19:72:@1206.4]
  wire [1:0] _T_1179; // @[Mux.scala 19:72:@1207.4]
  wire [1:0] _T_1181; // @[Mux.scala 19:72:@1208.4]
  wire [1:0] _T_1183; // @[Mux.scala 19:72:@1209.4]
  wire [1:0] _T_1185; // @[Mux.scala 19:72:@1210.4]
  wire [1:0] _T_1187; // @[Mux.scala 19:72:@1211.4]
  wire [1:0] _T_1189; // @[Mux.scala 19:72:@1212.4]
  wire [1:0] _T_1191; // @[Mux.scala 19:72:@1213.4]
  wire [1:0] _T_1193; // @[Mux.scala 19:72:@1214.4]
  wire [1:0] _T_1195; // @[Mux.scala 19:72:@1215.4]
  wire [1:0] _T_1197; // @[Mux.scala 19:72:@1216.4]
  wire [1:0] _T_1199; // @[Mux.scala 19:72:@1217.4]
  wire [1:0] _T_1201; // @[Mux.scala 19:72:@1218.4]
  wire [1:0] _T_1203; // @[Mux.scala 19:72:@1219.4]
  wire [1:0] _T_1205; // @[Mux.scala 19:72:@1220.4]
  wire [1:0] _T_1207; // @[Mux.scala 19:72:@1221.4]
  wire [1:0] _T_1209; // @[Mux.scala 19:72:@1222.4]
  wire [1:0] _T_1211; // @[Mux.scala 19:72:@1223.4]
  wire [1:0] _T_1213; // @[Mux.scala 19:72:@1224.4]
  wire [1:0] _T_1215; // @[Mux.scala 19:72:@1225.4]
  wire [1:0] _T_1217; // @[Mux.scala 19:72:@1226.4]
  wire [1:0] _T_1219; // @[Mux.scala 19:72:@1227.4]
  wire [1:0] _T_1221; // @[Mux.scala 19:72:@1228.4]
  wire [1:0] _T_1223; // @[Mux.scala 19:72:@1229.4]
  wire [1:0] _T_1225; // @[Mux.scala 19:72:@1230.4]
  wire [1:0] _T_1227; // @[Mux.scala 19:72:@1231.4]
  wire [1:0] _T_1229; // @[Mux.scala 19:72:@1232.4]
  wire [1:0] _T_1231; // @[Mux.scala 19:72:@1233.4]
  wire [1:0] _T_1233; // @[Mux.scala 19:72:@1234.4]
  wire [1:0] _T_1235; // @[Mux.scala 19:72:@1235.4]
  wire [1:0] _T_1237; // @[Mux.scala 19:72:@1236.4]
  wire [1:0] _T_1239; // @[Mux.scala 19:72:@1237.4]
  wire [1:0] _T_1241; // @[Mux.scala 19:72:@1238.4]
  wire [1:0] _T_1243; // @[Mux.scala 19:72:@1239.4]
  wire [1:0] _T_1245; // @[Mux.scala 19:72:@1240.4]
  wire [1:0] _T_1247; // @[Mux.scala 19:72:@1241.4]
  wire [1:0] _T_1249; // @[Mux.scala 19:72:@1242.4]
  wire [1:0] _T_1251; // @[Mux.scala 19:72:@1243.4]
  wire [1:0] _T_1253; // @[Mux.scala 19:72:@1244.4]
  wire [1:0] _T_1255; // @[Mux.scala 19:72:@1245.4]
  wire [1:0] _T_1257; // @[Mux.scala 19:72:@1246.4]
  wire [1:0] _T_1259; // @[Mux.scala 19:72:@1247.4]
  wire [1:0] _T_1261; // @[Mux.scala 19:72:@1248.4]
  wire [1:0] _T_1263; // @[Mux.scala 19:72:@1249.4]
  wire [1:0] _T_1265; // @[Mux.scala 19:72:@1250.4]
  wire [1:0] _T_1267; // @[Mux.scala 19:72:@1251.4]
  wire [1:0] _T_1269; // @[Mux.scala 19:72:@1252.4]
  wire [1:0] _T_1271; // @[Mux.scala 19:72:@1253.4]
  wire [1:0] _T_1273; // @[Mux.scala 19:72:@1254.4]
  wire [1:0] _T_1275; // @[Mux.scala 19:72:@1255.4]
  wire [1:0] _T_1277; // @[Mux.scala 19:72:@1256.4]
  wire [1:0] _T_1279; // @[Mux.scala 19:72:@1257.4]
  wire [1:0] _T_1281; // @[Mux.scala 19:72:@1258.4]
  wire [1:0] _T_1283; // @[Mux.scala 19:72:@1259.4]
  wire [1:0] _T_1285; // @[Mux.scala 19:72:@1260.4]
  wire [1:0] _T_1287; // @[Mux.scala 19:72:@1261.4]
  wire [1:0] _T_1289; // @[Mux.scala 19:72:@1262.4]
  wire [1:0] _T_1291; // @[Mux.scala 19:72:@1263.4]
  wire [1:0] _T_1293; // @[Mux.scala 19:72:@1264.4]
  wire [1:0] _T_1295; // @[Mux.scala 19:72:@1265.4]
  wire [1:0] _T_1296; // @[Mux.scala 19:72:@1266.4]
  wire [1:0] _T_1297; // @[Mux.scala 19:72:@1267.4]
  wire [1:0] _T_1298; // @[Mux.scala 19:72:@1268.4]
  wire [1:0] _T_1299; // @[Mux.scala 19:72:@1269.4]
  wire [1:0] _T_1300; // @[Mux.scala 19:72:@1270.4]
  wire [1:0] _T_1301; // @[Mux.scala 19:72:@1271.4]
  wire [1:0] _T_1302; // @[Mux.scala 19:72:@1272.4]
  wire [1:0] _T_1303; // @[Mux.scala 19:72:@1273.4]
  wire [1:0] _T_1304; // @[Mux.scala 19:72:@1274.4]
  wire [1:0] _T_1305; // @[Mux.scala 19:72:@1275.4]
  wire [1:0] _T_1306; // @[Mux.scala 19:72:@1276.4]
  wire [1:0] _T_1307; // @[Mux.scala 19:72:@1277.4]
  wire [1:0] _T_1308; // @[Mux.scala 19:72:@1278.4]
  wire [1:0] _T_1309; // @[Mux.scala 19:72:@1279.4]
  wire [1:0] _T_1310; // @[Mux.scala 19:72:@1280.4]
  wire [1:0] _T_1311; // @[Mux.scala 19:72:@1281.4]
  wire [1:0] _T_1312; // @[Mux.scala 19:72:@1282.4]
  wire [1:0] _T_1313; // @[Mux.scala 19:72:@1283.4]
  wire [1:0] _T_1314; // @[Mux.scala 19:72:@1284.4]
  wire [1:0] _T_1315; // @[Mux.scala 19:72:@1285.4]
  wire [1:0] _T_1316; // @[Mux.scala 19:72:@1286.4]
  wire [1:0] _T_1317; // @[Mux.scala 19:72:@1287.4]
  wire [1:0] _T_1318; // @[Mux.scala 19:72:@1288.4]
  wire [1:0] _T_1319; // @[Mux.scala 19:72:@1289.4]
  wire [1:0] _T_1320; // @[Mux.scala 19:72:@1290.4]
  wire [1:0] _T_1321; // @[Mux.scala 19:72:@1291.4]
  wire [1:0] _T_1322; // @[Mux.scala 19:72:@1292.4]
  wire [1:0] _T_1323; // @[Mux.scala 19:72:@1293.4]
  wire [1:0] _T_1324; // @[Mux.scala 19:72:@1294.4]
  wire [1:0] _T_1325; // @[Mux.scala 19:72:@1295.4]
  wire [1:0] _T_1326; // @[Mux.scala 19:72:@1296.4]
  wire [1:0] _T_1327; // @[Mux.scala 19:72:@1297.4]
  wire [1:0] _T_1328; // @[Mux.scala 19:72:@1298.4]
  wire [1:0] _T_1329; // @[Mux.scala 19:72:@1299.4]
  wire [1:0] _T_1330; // @[Mux.scala 19:72:@1300.4]
  wire [1:0] _T_1331; // @[Mux.scala 19:72:@1301.4]
  wire [1:0] _T_1332; // @[Mux.scala 19:72:@1302.4]
  wire [1:0] _T_1333; // @[Mux.scala 19:72:@1303.4]
  wire [1:0] _T_1334; // @[Mux.scala 19:72:@1304.4]
  wire [1:0] _T_1335; // @[Mux.scala 19:72:@1305.4]
  wire [1:0] _T_1336; // @[Mux.scala 19:72:@1306.4]
  wire [1:0] _T_1337; // @[Mux.scala 19:72:@1307.4]
  wire [1:0] _T_1338; // @[Mux.scala 19:72:@1308.4]
  wire [1:0] _T_1339; // @[Mux.scala 19:72:@1309.4]
  wire [1:0] _T_1340; // @[Mux.scala 19:72:@1310.4]
  wire [1:0] _T_1341; // @[Mux.scala 19:72:@1311.4]
  wire [1:0] _T_1342; // @[Mux.scala 19:72:@1312.4]
  wire [1:0] _T_1343; // @[Mux.scala 19:72:@1313.4]
  wire [1:0] _T_1344; // @[Mux.scala 19:72:@1314.4]
  wire [1:0] _T_1345; // @[Mux.scala 19:72:@1315.4]
  wire [1:0] _T_1346; // @[Mux.scala 19:72:@1316.4]
  wire [1:0] _T_1347; // @[Mux.scala 19:72:@1317.4]
  wire [1:0] _T_1348; // @[Mux.scala 19:72:@1318.4]
  wire [1:0] _T_1349; // @[Mux.scala 19:72:@1319.4]
  wire [1:0] _T_1350; // @[Mux.scala 19:72:@1320.4]
  wire [1:0] _T_1351; // @[Mux.scala 19:72:@1321.4]
  wire [1:0] _T_1352; // @[Mux.scala 19:72:@1322.4]
  wire [1:0] _T_1353; // @[Mux.scala 19:72:@1323.4]
  wire [1:0] _T_1354; // @[Mux.scala 19:72:@1324.4]
  wire [1:0] _T_1355; // @[Mux.scala 19:72:@1325.4]
  wire [1:0] _T_1356; // @[Mux.scala 19:72:@1326.4]
  wire [1:0] _T_1357; // @[Mux.scala 19:72:@1327.4]
  wire [1:0] predict_hcount; // @[Mux.scala 19:72:@1328.4]
  wire  _T_1362; // @[BTB.scala 76:35:@1332.4]
  wire  _T_1364; // @[BTB.scala 67:36:@1333.4]
  wire  _T_1365; // @[BTB.scala 67:67:@1334.4]
  wire  _T_1367; // @[BTB.scala 67:60:@1335.4]
  wire  _T_1368; // @[BTB.scala 67:57:@1336.4]
  wire  _T_1370; // @[BTB.scala 67:28:@1337.4]
  wire  _T_1372; // @[BTB.scala 67:82:@1338.4]
  wire  _T_1373; // @[BTB.scala 67:72:@1339.4]
  wire [31:0] _T_1374; // @[BTB.scala 67:27:@1340.4]
  reg  fb_reg_valid; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_256;
  reg  fb_reg_redirect; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_257;
  reg [5:0] fb_reg_lfsr; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_258;
  reg [31:0] fb_reg_pc; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_259;
  reg [31:0] fb_reg_target; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_260;
  reg [1:0] fb_reg_btype; // @[BTB.scala 78:23:@1350.4]
  reg [31:0] _RAND_261;
  wire  _T_1382; // @[BTB.scala 90:36:@1356.4]
  wire  _T_1383; // @[BTB.scala 90:46:@1357.4]
  wire  _T_1384; // @[BTB.scala 90:40:@1358.4]
  wire [4:0] _T_1385; // @[BTB.scala 90:55:@1359.4]
  wire [5:0] _T_1386; // @[Cat.scala 30:58:@1360.4]
  wire  _T_1388; // @[BTB.scala 114:42:@1363.4]
  wire  _T_1389; // @[BTB.scala 114:42:@1364.4]
  wire  _T_1390; // @[BTB.scala 114:42:@1365.4]
  wire  _T_1391; // @[BTB.scala 114:42:@1366.4]
  wire  _T_1392; // @[BTB.scala 114:42:@1367.4]
  wire  _T_1393; // @[BTB.scala 114:42:@1368.4]
  wire  _T_1394; // @[BTB.scala 114:42:@1369.4]
  wire  _T_1395; // @[BTB.scala 114:42:@1370.4]
  wire  _T_1396; // @[BTB.scala 114:42:@1371.4]
  wire  _T_1397; // @[BTB.scala 114:42:@1372.4]
  wire  _T_1398; // @[BTB.scala 114:42:@1373.4]
  wire  _T_1399; // @[BTB.scala 114:42:@1374.4]
  wire  _T_1400; // @[BTB.scala 114:42:@1375.4]
  wire  _T_1401; // @[BTB.scala 114:42:@1376.4]
  wire  _T_1402; // @[BTB.scala 114:42:@1377.4]
  wire  _T_1403; // @[BTB.scala 114:42:@1378.4]
  wire  _T_1404; // @[BTB.scala 114:42:@1379.4]
  wire  _T_1405; // @[BTB.scala 114:42:@1380.4]
  wire  _T_1406; // @[BTB.scala 114:42:@1381.4]
  wire  _T_1407; // @[BTB.scala 114:42:@1382.4]
  wire  _T_1408; // @[BTB.scala 114:42:@1383.4]
  wire  _T_1409; // @[BTB.scala 114:42:@1384.4]
  wire  _T_1410; // @[BTB.scala 114:42:@1385.4]
  wire  _T_1411; // @[BTB.scala 114:42:@1386.4]
  wire  _T_1412; // @[BTB.scala 114:42:@1387.4]
  wire  _T_1413; // @[BTB.scala 114:42:@1388.4]
  wire  _T_1414; // @[BTB.scala 114:42:@1389.4]
  wire  _T_1415; // @[BTB.scala 114:42:@1390.4]
  wire  _T_1416; // @[BTB.scala 114:42:@1391.4]
  wire  _T_1417; // @[BTB.scala 114:42:@1392.4]
  wire  _T_1418; // @[BTB.scala 114:42:@1393.4]
  wire  _T_1419; // @[BTB.scala 114:42:@1394.4]
  wire  _T_1420; // @[BTB.scala 114:42:@1395.4]
  wire  _T_1421; // @[BTB.scala 114:42:@1396.4]
  wire  _T_1422; // @[BTB.scala 114:42:@1397.4]
  wire  _T_1423; // @[BTB.scala 114:42:@1398.4]
  wire  _T_1424; // @[BTB.scala 114:42:@1399.4]
  wire  _T_1425; // @[BTB.scala 114:42:@1400.4]
  wire  _T_1426; // @[BTB.scala 114:42:@1401.4]
  wire  _T_1427; // @[BTB.scala 114:42:@1402.4]
  wire  _T_1428; // @[BTB.scala 114:42:@1403.4]
  wire  _T_1429; // @[BTB.scala 114:42:@1404.4]
  wire  _T_1430; // @[BTB.scala 114:42:@1405.4]
  wire  _T_1431; // @[BTB.scala 114:42:@1406.4]
  wire  _T_1432; // @[BTB.scala 114:42:@1407.4]
  wire  _T_1433; // @[BTB.scala 114:42:@1408.4]
  wire  _T_1434; // @[BTB.scala 114:42:@1409.4]
  wire  _T_1435; // @[BTB.scala 114:42:@1410.4]
  wire  _T_1436; // @[BTB.scala 114:42:@1411.4]
  wire  _T_1437; // @[BTB.scala 114:42:@1412.4]
  wire  _T_1438; // @[BTB.scala 114:42:@1413.4]
  wire  _T_1439; // @[BTB.scala 114:42:@1414.4]
  wire  _T_1440; // @[BTB.scala 114:42:@1415.4]
  wire  _T_1441; // @[BTB.scala 114:42:@1416.4]
  wire  _T_1442; // @[BTB.scala 114:42:@1417.4]
  wire  _T_1443; // @[BTB.scala 114:42:@1418.4]
  wire  _T_1444; // @[BTB.scala 114:42:@1419.4]
  wire  _T_1445; // @[BTB.scala 114:42:@1420.4]
  wire  _T_1446; // @[BTB.scala 114:42:@1421.4]
  wire  _T_1447; // @[BTB.scala 114:42:@1422.4]
  wire  _T_1448; // @[BTB.scala 114:42:@1423.4]
  wire  _T_1449; // @[BTB.scala 114:42:@1424.4]
  wire  _T_1450; // @[BTB.scala 114:42:@1425.4]
  wire  _T_1451; // @[BTB.scala 114:42:@1426.4]
  wire [7:0] _T_1528; // @[BTB.scala 114:58:@1498.4]
  wire [15:0] _T_1536; // @[BTB.scala 114:58:@1506.4]
  wire [7:0] _T_1543; // @[BTB.scala 114:58:@1513.4]
  wire [31:0] _T_1552; // @[BTB.scala 114:58:@1522.4]
  wire [7:0] _T_1559; // @[BTB.scala 114:58:@1529.4]
  wire [15:0] _T_1567; // @[BTB.scala 114:58:@1537.4]
  wire [7:0] _T_1574; // @[BTB.scala 114:58:@1544.4]
  wire [31:0] _T_1583; // @[BTB.scala 114:58:@1553.4]
  wire [63:0] _T_1584; // @[BTB.scala 114:58:@1554.4]
  wire [63:0] fb_wire_lookup; // @[BTB.scala 114:65:@1747.4]
  wire  _T_1847; // @[Mux.scala 21:36:@1749.4]
  wire  _T_1848; // @[Mux.scala 21:36:@1750.4]
  wire  _T_1849; // @[Mux.scala 21:36:@1751.4]
  wire  _T_1850; // @[Mux.scala 21:36:@1752.4]
  wire  _T_1851; // @[Mux.scala 21:36:@1753.4]
  wire  _T_1852; // @[Mux.scala 21:36:@1754.4]
  wire  _T_1853; // @[Mux.scala 21:36:@1755.4]
  wire  _T_1854; // @[Mux.scala 21:36:@1756.4]
  wire  _T_1855; // @[Mux.scala 21:36:@1757.4]
  wire  _T_1856; // @[Mux.scala 21:36:@1758.4]
  wire  _T_1857; // @[Mux.scala 21:36:@1759.4]
  wire  _T_1858; // @[Mux.scala 21:36:@1760.4]
  wire  _T_1859; // @[Mux.scala 21:36:@1761.4]
  wire  _T_1860; // @[Mux.scala 21:36:@1762.4]
  wire  _T_1861; // @[Mux.scala 21:36:@1763.4]
  wire  _T_1862; // @[Mux.scala 21:36:@1764.4]
  wire  _T_1863; // @[Mux.scala 21:36:@1765.4]
  wire  _T_1864; // @[Mux.scala 21:36:@1766.4]
  wire  _T_1865; // @[Mux.scala 21:36:@1767.4]
  wire  _T_1866; // @[Mux.scala 21:36:@1768.4]
  wire  _T_1867; // @[Mux.scala 21:36:@1769.4]
  wire  _T_1868; // @[Mux.scala 21:36:@1770.4]
  wire  _T_1869; // @[Mux.scala 21:36:@1771.4]
  wire  _T_1870; // @[Mux.scala 21:36:@1772.4]
  wire  _T_1871; // @[Mux.scala 21:36:@1773.4]
  wire  _T_1872; // @[Mux.scala 21:36:@1774.4]
  wire  _T_1873; // @[Mux.scala 21:36:@1775.4]
  wire  _T_1874; // @[Mux.scala 21:36:@1776.4]
  wire  _T_1875; // @[Mux.scala 21:36:@1777.4]
  wire  _T_1876; // @[Mux.scala 21:36:@1778.4]
  wire  _T_1877; // @[Mux.scala 21:36:@1779.4]
  wire  _T_1878; // @[Mux.scala 21:36:@1780.4]
  wire  _T_1879; // @[Mux.scala 21:36:@1781.4]
  wire  _T_1880; // @[Mux.scala 21:36:@1782.4]
  wire  _T_1881; // @[Mux.scala 21:36:@1783.4]
  wire  _T_1882; // @[Mux.scala 21:36:@1784.4]
  wire  _T_1883; // @[Mux.scala 21:36:@1785.4]
  wire  _T_1884; // @[Mux.scala 21:36:@1786.4]
  wire  _T_1885; // @[Mux.scala 21:36:@1787.4]
  wire  _T_1886; // @[Mux.scala 21:36:@1788.4]
  wire  _T_1887; // @[Mux.scala 21:36:@1789.4]
  wire  _T_1888; // @[Mux.scala 21:36:@1790.4]
  wire  _T_1889; // @[Mux.scala 21:36:@1791.4]
  wire  _T_1890; // @[Mux.scala 21:36:@1792.4]
  wire  _T_1891; // @[Mux.scala 21:36:@1793.4]
  wire  _T_1892; // @[Mux.scala 21:36:@1794.4]
  wire  _T_1893; // @[Mux.scala 21:36:@1795.4]
  wire  _T_1894; // @[Mux.scala 21:36:@1796.4]
  wire  _T_1895; // @[Mux.scala 21:36:@1797.4]
  wire  _T_1896; // @[Mux.scala 21:36:@1798.4]
  wire  _T_1897; // @[Mux.scala 21:36:@1799.4]
  wire  _T_1898; // @[Mux.scala 21:36:@1800.4]
  wire  _T_1899; // @[Mux.scala 21:36:@1801.4]
  wire  _T_1900; // @[Mux.scala 21:36:@1802.4]
  wire  _T_1901; // @[Mux.scala 21:36:@1803.4]
  wire  _T_1902; // @[Mux.scala 21:36:@1804.4]
  wire  _T_1903; // @[Mux.scala 21:36:@1805.4]
  wire  _T_1904; // @[Mux.scala 21:36:@1806.4]
  wire  _T_1905; // @[Mux.scala 21:36:@1807.4]
  wire  _T_1906; // @[Mux.scala 21:36:@1808.4]
  wire  _T_1907; // @[Mux.scala 21:36:@1809.4]
  wire  _T_1908; // @[Mux.scala 21:36:@1810.4]
  wire  _T_1909; // @[Mux.scala 21:36:@1811.4]
  wire  _T_1910; // @[Mux.scala 21:36:@1812.4]
  wire [1:0] _T_1913; // @[Mux.scala 19:72:@1813.4]
  wire [1:0] _T_1915; // @[Mux.scala 19:72:@1814.4]
  wire [1:0] _T_1917; // @[Mux.scala 19:72:@1815.4]
  wire [1:0] _T_1919; // @[Mux.scala 19:72:@1816.4]
  wire [1:0] _T_1921; // @[Mux.scala 19:72:@1817.4]
  wire [1:0] _T_1923; // @[Mux.scala 19:72:@1818.4]
  wire [1:0] _T_1925; // @[Mux.scala 19:72:@1819.4]
  wire [1:0] _T_1927; // @[Mux.scala 19:72:@1820.4]
  wire [1:0] _T_1929; // @[Mux.scala 19:72:@1821.4]
  wire [1:0] _T_1931; // @[Mux.scala 19:72:@1822.4]
  wire [1:0] _T_1933; // @[Mux.scala 19:72:@1823.4]
  wire [1:0] _T_1935; // @[Mux.scala 19:72:@1824.4]
  wire [1:0] _T_1937; // @[Mux.scala 19:72:@1825.4]
  wire [1:0] _T_1939; // @[Mux.scala 19:72:@1826.4]
  wire [1:0] _T_1941; // @[Mux.scala 19:72:@1827.4]
  wire [1:0] _T_1943; // @[Mux.scala 19:72:@1828.4]
  wire [1:0] _T_1945; // @[Mux.scala 19:72:@1829.4]
  wire [1:0] _T_1947; // @[Mux.scala 19:72:@1830.4]
  wire [1:0] _T_1949; // @[Mux.scala 19:72:@1831.4]
  wire [1:0] _T_1951; // @[Mux.scala 19:72:@1832.4]
  wire [1:0] _T_1953; // @[Mux.scala 19:72:@1833.4]
  wire [1:0] _T_1955; // @[Mux.scala 19:72:@1834.4]
  wire [1:0] _T_1957; // @[Mux.scala 19:72:@1835.4]
  wire [1:0] _T_1959; // @[Mux.scala 19:72:@1836.4]
  wire [1:0] _T_1961; // @[Mux.scala 19:72:@1837.4]
  wire [1:0] _T_1963; // @[Mux.scala 19:72:@1838.4]
  wire [1:0] _T_1965; // @[Mux.scala 19:72:@1839.4]
  wire [1:0] _T_1967; // @[Mux.scala 19:72:@1840.4]
  wire [1:0] _T_1969; // @[Mux.scala 19:72:@1841.4]
  wire [1:0] _T_1971; // @[Mux.scala 19:72:@1842.4]
  wire [1:0] _T_1973; // @[Mux.scala 19:72:@1843.4]
  wire [1:0] _T_1975; // @[Mux.scala 19:72:@1844.4]
  wire [1:0] _T_1977; // @[Mux.scala 19:72:@1845.4]
  wire [1:0] _T_1979; // @[Mux.scala 19:72:@1846.4]
  wire [1:0] _T_1981; // @[Mux.scala 19:72:@1847.4]
  wire [1:0] _T_1983; // @[Mux.scala 19:72:@1848.4]
  wire [1:0] _T_1985; // @[Mux.scala 19:72:@1849.4]
  wire [1:0] _T_1987; // @[Mux.scala 19:72:@1850.4]
  wire [1:0] _T_1989; // @[Mux.scala 19:72:@1851.4]
  wire [1:0] _T_1991; // @[Mux.scala 19:72:@1852.4]
  wire [1:0] _T_1993; // @[Mux.scala 19:72:@1853.4]
  wire [1:0] _T_1995; // @[Mux.scala 19:72:@1854.4]
  wire [1:0] _T_1997; // @[Mux.scala 19:72:@1855.4]
  wire [1:0] _T_1999; // @[Mux.scala 19:72:@1856.4]
  wire [1:0] _T_2001; // @[Mux.scala 19:72:@1857.4]
  wire [1:0] _T_2003; // @[Mux.scala 19:72:@1858.4]
  wire [1:0] _T_2005; // @[Mux.scala 19:72:@1859.4]
  wire [1:0] _T_2007; // @[Mux.scala 19:72:@1860.4]
  wire [1:0] _T_2009; // @[Mux.scala 19:72:@1861.4]
  wire [1:0] _T_2011; // @[Mux.scala 19:72:@1862.4]
  wire [1:0] _T_2013; // @[Mux.scala 19:72:@1863.4]
  wire [1:0] _T_2015; // @[Mux.scala 19:72:@1864.4]
  wire [1:0] _T_2017; // @[Mux.scala 19:72:@1865.4]
  wire [1:0] _T_2019; // @[Mux.scala 19:72:@1866.4]
  wire [1:0] _T_2021; // @[Mux.scala 19:72:@1867.4]
  wire [1:0] _T_2023; // @[Mux.scala 19:72:@1868.4]
  wire [1:0] _T_2025; // @[Mux.scala 19:72:@1869.4]
  wire [1:0] _T_2027; // @[Mux.scala 19:72:@1870.4]
  wire [1:0] _T_2029; // @[Mux.scala 19:72:@1871.4]
  wire [1:0] _T_2031; // @[Mux.scala 19:72:@1872.4]
  wire [1:0] _T_2033; // @[Mux.scala 19:72:@1873.4]
  wire [1:0] _T_2035; // @[Mux.scala 19:72:@1874.4]
  wire [1:0] _T_2037; // @[Mux.scala 19:72:@1875.4]
  wire [1:0] _T_2039; // @[Mux.scala 19:72:@1876.4]
  wire [1:0] _T_2040; // @[Mux.scala 19:72:@1877.4]
  wire [1:0] _T_2041; // @[Mux.scala 19:72:@1878.4]
  wire [1:0] _T_2042; // @[Mux.scala 19:72:@1879.4]
  wire [1:0] _T_2043; // @[Mux.scala 19:72:@1880.4]
  wire [1:0] _T_2044; // @[Mux.scala 19:72:@1881.4]
  wire [1:0] _T_2045; // @[Mux.scala 19:72:@1882.4]
  wire [1:0] _T_2046; // @[Mux.scala 19:72:@1883.4]
  wire [1:0] _T_2047; // @[Mux.scala 19:72:@1884.4]
  wire [1:0] _T_2048; // @[Mux.scala 19:72:@1885.4]
  wire [1:0] _T_2049; // @[Mux.scala 19:72:@1886.4]
  wire [1:0] _T_2050; // @[Mux.scala 19:72:@1887.4]
  wire [1:0] _T_2051; // @[Mux.scala 19:72:@1888.4]
  wire [1:0] _T_2052; // @[Mux.scala 19:72:@1889.4]
  wire [1:0] _T_2053; // @[Mux.scala 19:72:@1890.4]
  wire [1:0] _T_2054; // @[Mux.scala 19:72:@1891.4]
  wire [1:0] _T_2055; // @[Mux.scala 19:72:@1892.4]
  wire [1:0] _T_2056; // @[Mux.scala 19:72:@1893.4]
  wire [1:0] _T_2057; // @[Mux.scala 19:72:@1894.4]
  wire [1:0] _T_2058; // @[Mux.scala 19:72:@1895.4]
  wire [1:0] _T_2059; // @[Mux.scala 19:72:@1896.4]
  wire [1:0] _T_2060; // @[Mux.scala 19:72:@1897.4]
  wire [1:0] _T_2061; // @[Mux.scala 19:72:@1898.4]
  wire [1:0] _T_2062; // @[Mux.scala 19:72:@1899.4]
  wire [1:0] _T_2063; // @[Mux.scala 19:72:@1900.4]
  wire [1:0] _T_2064; // @[Mux.scala 19:72:@1901.4]
  wire [1:0] _T_2065; // @[Mux.scala 19:72:@1902.4]
  wire [1:0] _T_2066; // @[Mux.scala 19:72:@1903.4]
  wire [1:0] _T_2067; // @[Mux.scala 19:72:@1904.4]
  wire [1:0] _T_2068; // @[Mux.scala 19:72:@1905.4]
  wire [1:0] _T_2069; // @[Mux.scala 19:72:@1906.4]
  wire [1:0] _T_2070; // @[Mux.scala 19:72:@1907.4]
  wire [1:0] _T_2071; // @[Mux.scala 19:72:@1908.4]
  wire [1:0] _T_2072; // @[Mux.scala 19:72:@1909.4]
  wire [1:0] _T_2073; // @[Mux.scala 19:72:@1910.4]
  wire [1:0] _T_2074; // @[Mux.scala 19:72:@1911.4]
  wire [1:0] _T_2075; // @[Mux.scala 19:72:@1912.4]
  wire [1:0] _T_2076; // @[Mux.scala 19:72:@1913.4]
  wire [1:0] _T_2077; // @[Mux.scala 19:72:@1914.4]
  wire [1:0] _T_2078; // @[Mux.scala 19:72:@1915.4]
  wire [1:0] _T_2079; // @[Mux.scala 19:72:@1916.4]
  wire [1:0] _T_2080; // @[Mux.scala 19:72:@1917.4]
  wire [1:0] _T_2081; // @[Mux.scala 19:72:@1918.4]
  wire [1:0] _T_2082; // @[Mux.scala 19:72:@1919.4]
  wire [1:0] _T_2083; // @[Mux.scala 19:72:@1920.4]
  wire [1:0] _T_2084; // @[Mux.scala 19:72:@1921.4]
  wire [1:0] _T_2085; // @[Mux.scala 19:72:@1922.4]
  wire [1:0] _T_2086; // @[Mux.scala 19:72:@1923.4]
  wire [1:0] _T_2087; // @[Mux.scala 19:72:@1924.4]
  wire [1:0] _T_2088; // @[Mux.scala 19:72:@1925.4]
  wire [1:0] _T_2089; // @[Mux.scala 19:72:@1926.4]
  wire [1:0] _T_2090; // @[Mux.scala 19:72:@1927.4]
  wire [1:0] _T_2091; // @[Mux.scala 19:72:@1928.4]
  wire [1:0] _T_2092; // @[Mux.scala 19:72:@1929.4]
  wire [1:0] _T_2093; // @[Mux.scala 19:72:@1930.4]
  wire [1:0] _T_2094; // @[Mux.scala 19:72:@1931.4]
  wire [1:0] _T_2095; // @[Mux.scala 19:72:@1932.4]
  wire [1:0] _T_2096; // @[Mux.scala 19:72:@1933.4]
  wire [1:0] _T_2097; // @[Mux.scala 19:72:@1934.4]
  wire [1:0] _T_2098; // @[Mux.scala 19:72:@1935.4]
  wire [1:0] _T_2099; // @[Mux.scala 19:72:@1936.4]
  wire [1:0] _T_2100; // @[Mux.scala 19:72:@1937.4]
  wire [1:0] _T_2101; // @[Mux.scala 19:72:@1938.4]
  wire [1:0] fb_wire_hcount; // @[Mux.scala 19:72:@1939.4]
  wire  _T_2106; // @[BTB.scala 112:30:@1943.4]
  wire [31:0] _T_2107; // @[OneHot.scala 26:18:@1944.4]
  wire [31:0] _T_2108; // @[OneHot.scala 27:18:@1945.4]
  wire  _T_2110; // @[OneHot.scala 28:14:@1946.4]
  wire [31:0] _T_2111; // @[OneHot.scala 28:28:@1947.4]
  wire [15:0] _T_2112; // @[OneHot.scala 26:18:@1948.4]
  wire [15:0] _T_2113; // @[OneHot.scala 27:18:@1949.4]
  wire  _T_2115; // @[OneHot.scala 28:14:@1950.4]
  wire [15:0] _T_2116; // @[OneHot.scala 28:28:@1951.4]
  wire [7:0] _T_2117; // @[OneHot.scala 26:18:@1952.4]
  wire [7:0] _T_2118; // @[OneHot.scala 27:18:@1953.4]
  wire  _T_2120; // @[OneHot.scala 28:14:@1954.4]
  wire [7:0] _T_2121; // @[OneHot.scala 28:28:@1955.4]
  wire [3:0] _T_2122; // @[OneHot.scala 26:18:@1956.4]
  wire [3:0] _T_2123; // @[OneHot.scala 27:18:@1957.4]
  wire  _T_2125; // @[OneHot.scala 28:14:@1958.4]
  wire [3:0] _T_2126; // @[OneHot.scala 28:28:@1959.4]
  wire [1:0] _T_2127; // @[OneHot.scala 26:18:@1960.4]
  wire [1:0] _T_2128; // @[OneHot.scala 27:18:@1961.4]
  wire  _T_2130; // @[OneHot.scala 28:14:@1962.4]
  wire [1:0] _T_2131; // @[OneHot.scala 28:28:@1963.4]
  wire  _T_2132; // @[CircuitMath.scala 30:8:@1964.4]
  wire [5:0] _T_2137; // @[Cat.scala 30:58:@1969.4]
  wire [63:0] _T_2399; // @[BTB.scala 118:19:@2162.4]
  wire  _T_2401; // @[BTB.scala 118:19:@2163.4]
  wire  _T_2664; // @[OneHot.scala 39:40:@2357.4]
  wire  _T_2665; // @[OneHot.scala 39:40:@2358.4]
  wire  _T_2666; // @[OneHot.scala 39:40:@2359.4]
  wire  _T_2667; // @[OneHot.scala 39:40:@2360.4]
  wire  _T_2668; // @[OneHot.scala 39:40:@2361.4]
  wire  _T_2669; // @[OneHot.scala 39:40:@2362.4]
  wire  _T_2670; // @[OneHot.scala 39:40:@2363.4]
  wire  _T_2671; // @[OneHot.scala 39:40:@2364.4]
  wire  _T_2672; // @[OneHot.scala 39:40:@2365.4]
  wire  _T_2673; // @[OneHot.scala 39:40:@2366.4]
  wire  _T_2674; // @[OneHot.scala 39:40:@2367.4]
  wire  _T_2675; // @[OneHot.scala 39:40:@2368.4]
  wire  _T_2676; // @[OneHot.scala 39:40:@2369.4]
  wire  _T_2677; // @[OneHot.scala 39:40:@2370.4]
  wire  _T_2678; // @[OneHot.scala 39:40:@2371.4]
  wire  _T_2679; // @[OneHot.scala 39:40:@2372.4]
  wire  _T_2680; // @[OneHot.scala 39:40:@2373.4]
  wire  _T_2681; // @[OneHot.scala 39:40:@2374.4]
  wire  _T_2682; // @[OneHot.scala 39:40:@2375.4]
  wire  _T_2683; // @[OneHot.scala 39:40:@2376.4]
  wire  _T_2684; // @[OneHot.scala 39:40:@2377.4]
  wire  _T_2685; // @[OneHot.scala 39:40:@2378.4]
  wire  _T_2686; // @[OneHot.scala 39:40:@2379.4]
  wire  _T_2687; // @[OneHot.scala 39:40:@2380.4]
  wire  _T_2688; // @[OneHot.scala 39:40:@2381.4]
  wire  _T_2689; // @[OneHot.scala 39:40:@2382.4]
  wire  _T_2690; // @[OneHot.scala 39:40:@2383.4]
  wire  _T_2691; // @[OneHot.scala 39:40:@2384.4]
  wire  _T_2692; // @[OneHot.scala 39:40:@2385.4]
  wire  _T_2693; // @[OneHot.scala 39:40:@2386.4]
  wire  _T_2694; // @[OneHot.scala 39:40:@2387.4]
  wire  _T_2695; // @[OneHot.scala 39:40:@2388.4]
  wire  _T_2696; // @[OneHot.scala 39:40:@2389.4]
  wire  _T_2697; // @[OneHot.scala 39:40:@2390.4]
  wire  _T_2698; // @[OneHot.scala 39:40:@2391.4]
  wire  _T_2699; // @[OneHot.scala 39:40:@2392.4]
  wire  _T_2700; // @[OneHot.scala 39:40:@2393.4]
  wire  _T_2701; // @[OneHot.scala 39:40:@2394.4]
  wire  _T_2702; // @[OneHot.scala 39:40:@2395.4]
  wire  _T_2703; // @[OneHot.scala 39:40:@2396.4]
  wire  _T_2704; // @[OneHot.scala 39:40:@2397.4]
  wire  _T_2705; // @[OneHot.scala 39:40:@2398.4]
  wire  _T_2706; // @[OneHot.scala 39:40:@2399.4]
  wire  _T_2707; // @[OneHot.scala 39:40:@2400.4]
  wire  _T_2708; // @[OneHot.scala 39:40:@2401.4]
  wire  _T_2709; // @[OneHot.scala 39:40:@2402.4]
  wire  _T_2710; // @[OneHot.scala 39:40:@2403.4]
  wire  _T_2711; // @[OneHot.scala 39:40:@2404.4]
  wire  _T_2712; // @[OneHot.scala 39:40:@2405.4]
  wire  _T_2713; // @[OneHot.scala 39:40:@2406.4]
  wire  _T_2714; // @[OneHot.scala 39:40:@2407.4]
  wire  _T_2715; // @[OneHot.scala 39:40:@2408.4]
  wire  _T_2716; // @[OneHot.scala 39:40:@2409.4]
  wire  _T_2717; // @[OneHot.scala 39:40:@2410.4]
  wire  _T_2718; // @[OneHot.scala 39:40:@2411.4]
  wire  _T_2719; // @[OneHot.scala 39:40:@2412.4]
  wire  _T_2720; // @[OneHot.scala 39:40:@2413.4]
  wire  _T_2721; // @[OneHot.scala 39:40:@2414.4]
  wire  _T_2722; // @[OneHot.scala 39:40:@2415.4]
  wire  _T_2723; // @[OneHot.scala 39:40:@2416.4]
  wire  _T_2724; // @[OneHot.scala 39:40:@2417.4]
  wire  _T_2725; // @[OneHot.scala 39:40:@2418.4]
  wire  _T_2726; // @[OneHot.scala 39:40:@2419.4]
  wire [5:0] _T_2792; // @[Mux.scala 31:69:@2421.4]
  wire [5:0] _T_2793; // @[Mux.scala 31:69:@2422.4]
  wire [5:0] _T_2794; // @[Mux.scala 31:69:@2423.4]
  wire [5:0] _T_2795; // @[Mux.scala 31:69:@2424.4]
  wire [5:0] _T_2796; // @[Mux.scala 31:69:@2425.4]
  wire [5:0] _T_2797; // @[Mux.scala 31:69:@2426.4]
  wire [5:0] _T_2798; // @[Mux.scala 31:69:@2427.4]
  wire [5:0] _T_2799; // @[Mux.scala 31:69:@2428.4]
  wire [5:0] _T_2800; // @[Mux.scala 31:69:@2429.4]
  wire [5:0] _T_2801; // @[Mux.scala 31:69:@2430.4]
  wire [5:0] _T_2802; // @[Mux.scala 31:69:@2431.4]
  wire [5:0] _T_2803; // @[Mux.scala 31:69:@2432.4]
  wire [5:0] _T_2804; // @[Mux.scala 31:69:@2433.4]
  wire [5:0] _T_2805; // @[Mux.scala 31:69:@2434.4]
  wire [5:0] _T_2806; // @[Mux.scala 31:69:@2435.4]
  wire [5:0] _T_2807; // @[Mux.scala 31:69:@2436.4]
  wire [5:0] _T_2808; // @[Mux.scala 31:69:@2437.4]
  wire [5:0] _T_2809; // @[Mux.scala 31:69:@2438.4]
  wire [5:0] _T_2810; // @[Mux.scala 31:69:@2439.4]
  wire [5:0] _T_2811; // @[Mux.scala 31:69:@2440.4]
  wire [5:0] _T_2812; // @[Mux.scala 31:69:@2441.4]
  wire [5:0] _T_2813; // @[Mux.scala 31:69:@2442.4]
  wire [5:0] _T_2814; // @[Mux.scala 31:69:@2443.4]
  wire [5:0] _T_2815; // @[Mux.scala 31:69:@2444.4]
  wire [5:0] _T_2816; // @[Mux.scala 31:69:@2445.4]
  wire [5:0] _T_2817; // @[Mux.scala 31:69:@2446.4]
  wire [5:0] _T_2818; // @[Mux.scala 31:69:@2447.4]
  wire [5:0] _T_2819; // @[Mux.scala 31:69:@2448.4]
  wire [5:0] _T_2820; // @[Mux.scala 31:69:@2449.4]
  wire [5:0] _T_2821; // @[Mux.scala 31:69:@2450.4]
  wire [5:0] _T_2822; // @[Mux.scala 31:69:@2451.4]
  wire [5:0] _T_2823; // @[Mux.scala 31:69:@2452.4]
  wire [5:0] _T_2824; // @[Mux.scala 31:69:@2453.4]
  wire [5:0] _T_2825; // @[Mux.scala 31:69:@2454.4]
  wire [5:0] _T_2826; // @[Mux.scala 31:69:@2455.4]
  wire [5:0] _T_2827; // @[Mux.scala 31:69:@2456.4]
  wire [5:0] _T_2828; // @[Mux.scala 31:69:@2457.4]
  wire [5:0] _T_2829; // @[Mux.scala 31:69:@2458.4]
  wire [5:0] _T_2830; // @[Mux.scala 31:69:@2459.4]
  wire [5:0] _T_2831; // @[Mux.scala 31:69:@2460.4]
  wire [5:0] _T_2832; // @[Mux.scala 31:69:@2461.4]
  wire [5:0] _T_2833; // @[Mux.scala 31:69:@2462.4]
  wire [5:0] _T_2834; // @[Mux.scala 31:69:@2463.4]
  wire [5:0] _T_2835; // @[Mux.scala 31:69:@2464.4]
  wire [5:0] _T_2836; // @[Mux.scala 31:69:@2465.4]
  wire [5:0] _T_2837; // @[Mux.scala 31:69:@2466.4]
  wire [5:0] _T_2838; // @[Mux.scala 31:69:@2467.4]
  wire [5:0] _T_2839; // @[Mux.scala 31:69:@2468.4]
  wire [5:0] _T_2840; // @[Mux.scala 31:69:@2469.4]
  wire [5:0] _T_2841; // @[Mux.scala 31:69:@2470.4]
  wire [5:0] _T_2842; // @[Mux.scala 31:69:@2471.4]
  wire [5:0] _T_2843; // @[Mux.scala 31:69:@2472.4]
  wire [5:0] _T_2844; // @[Mux.scala 31:69:@2473.4]
  wire [5:0] _T_2845; // @[Mux.scala 31:69:@2474.4]
  wire [5:0] _T_2846; // @[Mux.scala 31:69:@2475.4]
  wire [5:0] _T_2847; // @[Mux.scala 31:69:@2476.4]
  wire [5:0] _T_2848; // @[Mux.scala 31:69:@2477.4]
  wire [5:0] _T_2849; // @[Mux.scala 31:69:@2478.4]
  wire [5:0] _T_2850; // @[Mux.scala 31:69:@2479.4]
  wire [5:0] _T_2851; // @[Mux.scala 31:69:@2480.4]
  wire [5:0] _T_2852; // @[Mux.scala 31:69:@2481.4]
  wire [5:0] _T_2853; // @[Mux.scala 31:69:@2482.4]
  wire [5:0] _T_2854; // @[Mux.scala 31:69:@2483.4]
  wire [5:0] _T_2855; // @[BTB.scala 118:8:@2484.4]
  wire [5:0] fb_wire_bindex; // @[BTB.scala 117:8:@2485.4]
  wire [31:0] _GEN_0; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_1; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_2; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_3; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_4; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_5; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_6; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_7; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_8; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_9; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_10; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_11; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_12; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_13; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_14; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_15; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_16; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_17; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_18; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_19; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_20; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_21; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_22; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_23; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_24; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_25; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_26; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_27; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_28; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_29; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_30; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_31; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_32; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_33; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_34; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_35; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_36; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_37; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_38; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_39; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_40; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_41; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_42; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_43; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_44; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_45; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_46; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_47; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_48; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_49; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_50; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_51; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_52; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_53; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_54; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_55; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_56; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_57; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_58; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_59; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_60; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_61; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_62; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_63; // @[BTB.scala 124:34:@2489.8]
  wire [31:0] _GEN_64; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_65; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_66; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_67; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_68; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_69; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_70; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_71; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_72; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_73; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_74; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_75; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_76; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_77; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_78; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_79; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_80; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_81; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_82; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_83; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_84; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_85; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_86; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_87; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_88; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_89; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_90; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_91; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_92; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_93; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_94; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_95; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_96; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_97; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_98; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_99; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_100; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_101; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_102; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_103; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_104; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_105; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_106; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_107; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_108; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_109; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_110; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_111; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_112; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_113; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_114; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_115; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_116; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_117; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_118; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_119; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_120; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_121; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_122; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_123; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_124; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_125; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_126; // @[BTB.scala 125:34:@2490.8]
  wire [31:0] _GEN_127; // @[BTB.scala 125:34:@2490.8]
  wire [1:0] _GEN_128; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_129; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_130; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_131; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_132; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_133; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_134; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_135; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_136; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_137; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_138; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_139; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_140; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_141; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_142; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_143; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_144; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_145; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_146; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_147; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_148; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_149; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_150; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_151; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_152; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_153; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_154; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_155; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_156; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_157; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_158; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_159; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_160; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_161; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_162; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_163; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_164; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_165; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_166; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_167; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_168; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_169; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_170; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_171; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_172; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_173; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_174; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_175; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_176; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_177; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_178; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_179; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_180; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_181; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_182; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_183; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_184; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_185; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_186; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_187; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_188; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_189; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_190; // @[BTB.scala 126:34:@2491.8]
  wire [1:0] _GEN_191; // @[BTB.scala 126:34:@2491.8]
  wire [31:0] _GEN_192; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_193; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_194; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_195; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_196; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_197; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_198; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_199; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_200; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_201; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_202; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_203; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_204; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_205; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_206; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_207; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_208; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_209; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_210; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_211; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_212; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_213; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_214; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_215; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_216; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_217; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_218; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_219; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_220; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_221; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_222; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_223; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_224; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_225; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_226; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_227; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_228; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_229; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_230; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_231; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_232; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_233; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_234; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_235; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_236; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_237; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_238; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_239; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_240; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_241; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_242; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_243; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_244; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_245; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_246; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_247; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_248; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_249; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_250; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_251; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_252; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_253; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_254; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_255; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_256; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_257; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_258; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_259; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_260; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_261; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_262; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_263; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_264; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_265; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_266; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_267; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_268; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_269; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_270; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_271; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_272; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_273; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_274; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_275; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_276; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_277; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_278; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_279; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_280; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_281; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_282; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_283; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_284; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_285; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_286; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_287; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_288; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_289; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_290; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_291; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_292; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_293; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_294; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_295; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_296; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_297; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_298; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_299; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_300; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_301; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_302; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_303; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_304; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_305; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_306; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_307; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_308; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_309; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_310; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_311; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_312; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_313; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_314; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_315; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_316; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_317; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_318; // @[BTB.scala 123:28:@2488.6]
  wire [31:0] _GEN_319; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_320; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_321; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_322; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_323; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_324; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_325; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_326; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_327; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_328; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_329; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_330; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_331; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_332; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_333; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_334; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_335; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_336; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_337; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_338; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_339; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_340; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_341; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_342; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_343; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_344; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_345; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_346; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_347; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_348; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_349; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_350; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_351; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_352; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_353; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_354; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_355; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_356; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_357; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_358; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_359; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_360; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_361; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_362; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_363; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_364; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_365; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_366; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_367; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_368; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_369; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_370; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_371; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_372; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_373; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_374; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_375; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_376; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_377; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_378; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_379; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_380; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_381; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_382; // @[BTB.scala 123:28:@2488.6]
  wire [1:0] _GEN_383; // @[BTB.scala 123:28:@2488.6]
  wire  _T_2858; // @[BTB.scala 128:24:@2493.6]
  wire  _T_2862; // @[BTB.scala 51:42:@2498.12]
  wire  _T_2863; // @[BTB.scala 51:49:@2499.12]
  wire  _T_2864; // @[BTB.scala 51:58:@2500.12]
  wire  _T_2866; // @[BTB.scala 51:56:@2501.12]
  wire  _T_2867; // @[BTB.scala 51:53:@2502.12]
  wire [1:0] _T_2868; // @[Cat.scala 30:58:@2503.12]
  wire [1:0] _GEN_384; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_385; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_386; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_387; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_388; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_389; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_390; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_391; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_392; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_393; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_394; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_395; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_396; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_397; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_398; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_399; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_400; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_401; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_402; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_403; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_404; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_405; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_406; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_407; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_408; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_409; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_410; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_411; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_412; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_413; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_414; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_415; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_416; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_417; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_418; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_419; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_420; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_421; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_422; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_423; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_424; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_425; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_426; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_427; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_428; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_429; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_430; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_431; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_432; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_433; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_434; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_435; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_436; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_437; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_438; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_439; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_440; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_441; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_442; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_443; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_444; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_445; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_446; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _GEN_447; // @[BTB.scala 131:38:@2504.12]
  wire [1:0] _T_2869; // @[BTB.scala 52:42:@2507.12]
  wire  _T_2871; // @[BTB.scala 52:42:@2508.12]
  wire  _T_2876; // @[BTB.scala 52:53:@2512.12]
  wire [1:0] _T_2877; // @[Cat.scala 30:58:@2513.12]
  wire [1:0] _GEN_448; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_449; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_450; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_451; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_452; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_453; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_454; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_455; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_456; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_457; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_458; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_459; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_460; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_461; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_462; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_463; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_464; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_465; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_466; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_467; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_468; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_469; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_470; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_471; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_472; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_473; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_474; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_475; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_476; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_477; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_478; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_479; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_480; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_481; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_482; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_483; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_484; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_485; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_486; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_487; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_488; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_489; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_490; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_491; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_492; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_493; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_494; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_495; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_496; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_497; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_498; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_499; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_500; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_501; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_502; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_503; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_504; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_505; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_506; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_507; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_508; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_509; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_510; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_511; // @[BTB.scala 133:38:@2514.12]
  wire [1:0] _GEN_512; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_513; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_514; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_515; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_516; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_517; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_518; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_519; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_520; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_521; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_522; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_523; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_524; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_525; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_526; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_527; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_528; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_529; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_530; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_531; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_532; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_533; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_534; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_535; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_536; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_537; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_538; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_539; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_540; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_541; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_542; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_543; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_544; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_545; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_546; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_547; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_548; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_549; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_550; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_551; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_552; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_553; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_554; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_555; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_556; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_557; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_558; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_559; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_560; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_561; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_562; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_563; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_564; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_565; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_566; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_567; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_568; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_569; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_570; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_571; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_572; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_573; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_574; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_575; // @[BTB.scala 130:32:@2497.10]
  wire [1:0] _GEN_576; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_577; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_578; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_579; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_580; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_581; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_582; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_583; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_584; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_585; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_586; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_587; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_588; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_589; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_590; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_591; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_592; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_593; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_594; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_595; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_596; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_597; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_598; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_599; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_600; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_601; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_602; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_603; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_604; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_605; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_606; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_607; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_608; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_609; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_610; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_611; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_612; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_613; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_614; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_615; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_616; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_617; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_618; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_619; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_620; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_621; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_622; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_623; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_624; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_625; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_626; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_627; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_628; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_629; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_630; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_631; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_632; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_633; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_634; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_635; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_636; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_637; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_638; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_639; // @[BTB.scala 136:36:@2519.12]
  wire [1:0] _GEN_640; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_641; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_642; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_643; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_644; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_645; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_646; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_647; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_648; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_649; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_650; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_651; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_652; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_653; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_654; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_655; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_656; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_657; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_658; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_659; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_660; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_661; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_662; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_663; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_664; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_665; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_666; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_667; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_668; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_669; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_670; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_671; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_672; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_673; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_674; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_675; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_676; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_677; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_678; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_679; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_680; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_681; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_682; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_683; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_684; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_685; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_686; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_687; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_688; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_689; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_690; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_691; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_692; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_693; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_694; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_695; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_696; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_697; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_698; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_699; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_700; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_701; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_702; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_703; // @[BTB.scala 135:35:@2518.10]
  wire [1:0] _GEN_704; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_705; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_706; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_707; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_708; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_709; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_710; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_711; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_712; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_713; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_714; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_715; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_716; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_717; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_718; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_719; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_720; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_721; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_722; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_723; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_724; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_725; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_726; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_727; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_728; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_729; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_730; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_731; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_732; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_733; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_734; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_735; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_736; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_737; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_738; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_739; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_740; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_741; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_742; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_743; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_744; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_745; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_746; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_747; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_748; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_749; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_750; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_751; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_752; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_753; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_754; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_755; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_756; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_757; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_758; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_759; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_760; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_761; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_762; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_763; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_764; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_765; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_766; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_767; // @[BTB.scala 129:28:@2496.8]
  wire [1:0] _GEN_768; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_769; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_770; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_771; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_772; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_773; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_774; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_775; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_776; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_777; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_778; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_779; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_780; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_781; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_782; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_783; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_784; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_785; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_786; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_787; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_788; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_789; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_790; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_791; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_792; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_793; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_794; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_795; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_796; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_797; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_798; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_799; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_800; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_801; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_802; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_803; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_804; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_805; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_806; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_807; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_808; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_809; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_810; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_811; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_812; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_813; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_814; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_815; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_816; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_817; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_818; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_819; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_820; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_821; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_822; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_823; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_824; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_825; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_826; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_827; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_828; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_829; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_830; // @[BTB.scala 128:46:@2494.6]
  wire [1:0] _GEN_831; // @[BTB.scala 128:46:@2494.6]
  wire [31:0] _GEN_832; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_833; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_834; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_835; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_836; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_837; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_838; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_839; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_840; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_841; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_842; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_843; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_844; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_845; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_846; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_847; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_848; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_849; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_850; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_851; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_852; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_853; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_854; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_855; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_856; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_857; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_858; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_859; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_860; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_861; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_862; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_863; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_864; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_865; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_866; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_867; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_868; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_869; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_870; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_871; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_872; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_873; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_874; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_875; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_876; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_877; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_878; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_879; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_880; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_881; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_882; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_883; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_884; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_885; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_886; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_887; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_888; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_889; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_890; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_891; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_892; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_893; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_894; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_895; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_896; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_897; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_898; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_899; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_900; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_901; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_902; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_903; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_904; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_905; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_906; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_907; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_908; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_909; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_910; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_911; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_912; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_913; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_914; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_915; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_916; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_917; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_918; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_919; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_920; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_921; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_922; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_923; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_924; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_925; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_926; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_927; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_928; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_929; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_930; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_931; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_932; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_933; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_934; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_935; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_936; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_937; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_938; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_939; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_940; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_941; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_942; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_943; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_944; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_945; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_946; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_947; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_948; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_949; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_950; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_951; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_952; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_953; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_954; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_955; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_956; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_957; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_958; // @[BTB.scala 122:23:@2487.4]
  wire [31:0] _GEN_959; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_960; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_961; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_962; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_963; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_964; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_965; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_966; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_967; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_968; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_969; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_970; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_971; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_972; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_973; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_974; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_975; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_976; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_977; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_978; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_979; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_980; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_981; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_982; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_983; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_984; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_985; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_986; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_987; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_988; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_989; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_990; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_991; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_992; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_993; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_994; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_995; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_996; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_997; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_998; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_999; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1000; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1001; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1002; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1003; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1004; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1005; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1006; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1007; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1008; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1009; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1010; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1011; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1012; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1013; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1014; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1015; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1016; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1017; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1018; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1019; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1020; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1021; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1022; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1023; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1024; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1025; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1026; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1027; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1028; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1029; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1030; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1031; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1032; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1033; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1034; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1035; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1036; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1037; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1038; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1039; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1040; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1041; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1042; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1043; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1044; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1045; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1046; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1047; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1048; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1049; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1050; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1051; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1052; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1053; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1054; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1055; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1056; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1057; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1058; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1059; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1060; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1061; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1062; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1063; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1064; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1065; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1066; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1067; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1068; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1069; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1070; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1071; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1072; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1073; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1074; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1075; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1076; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1077; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1078; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1079; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1080; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1081; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1082; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1083; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1084; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1085; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1086; // @[BTB.scala 122:23:@2487.4]
  wire [1:0] _GEN_1087; // @[BTB.scala 122:23:@2487.4]
  assign _T_125 = btb_pc_0 == io_if_pc; // @[BTB.scala 70:42:@361.4]
  assign _T_126 = btb_pc_1 == io_if_pc; // @[BTB.scala 70:42:@362.4]
  assign _T_127 = btb_pc_2 == io_if_pc; // @[BTB.scala 70:42:@363.4]
  assign _T_128 = btb_pc_3 == io_if_pc; // @[BTB.scala 70:42:@364.4]
  assign _T_129 = btb_pc_4 == io_if_pc; // @[BTB.scala 70:42:@365.4]
  assign _T_130 = btb_pc_5 == io_if_pc; // @[BTB.scala 70:42:@366.4]
  assign _T_131 = btb_pc_6 == io_if_pc; // @[BTB.scala 70:42:@367.4]
  assign _T_132 = btb_pc_7 == io_if_pc; // @[BTB.scala 70:42:@368.4]
  assign _T_133 = btb_pc_8 == io_if_pc; // @[BTB.scala 70:42:@369.4]
  assign _T_134 = btb_pc_9 == io_if_pc; // @[BTB.scala 70:42:@370.4]
  assign _T_135 = btb_pc_10 == io_if_pc; // @[BTB.scala 70:42:@371.4]
  assign _T_136 = btb_pc_11 == io_if_pc; // @[BTB.scala 70:42:@372.4]
  assign _T_137 = btb_pc_12 == io_if_pc; // @[BTB.scala 70:42:@373.4]
  assign _T_138 = btb_pc_13 == io_if_pc; // @[BTB.scala 70:42:@374.4]
  assign _T_139 = btb_pc_14 == io_if_pc; // @[BTB.scala 70:42:@375.4]
  assign _T_140 = btb_pc_15 == io_if_pc; // @[BTB.scala 70:42:@376.4]
  assign _T_141 = btb_pc_16 == io_if_pc; // @[BTB.scala 70:42:@377.4]
  assign _T_142 = btb_pc_17 == io_if_pc; // @[BTB.scala 70:42:@378.4]
  assign _T_143 = btb_pc_18 == io_if_pc; // @[BTB.scala 70:42:@379.4]
  assign _T_144 = btb_pc_19 == io_if_pc; // @[BTB.scala 70:42:@380.4]
  assign _T_145 = btb_pc_20 == io_if_pc; // @[BTB.scala 70:42:@381.4]
  assign _T_146 = btb_pc_21 == io_if_pc; // @[BTB.scala 70:42:@382.4]
  assign _T_147 = btb_pc_22 == io_if_pc; // @[BTB.scala 70:42:@383.4]
  assign _T_148 = btb_pc_23 == io_if_pc; // @[BTB.scala 70:42:@384.4]
  assign _T_149 = btb_pc_24 == io_if_pc; // @[BTB.scala 70:42:@385.4]
  assign _T_150 = btb_pc_25 == io_if_pc; // @[BTB.scala 70:42:@386.4]
  assign _T_151 = btb_pc_26 == io_if_pc; // @[BTB.scala 70:42:@387.4]
  assign _T_152 = btb_pc_27 == io_if_pc; // @[BTB.scala 70:42:@388.4]
  assign _T_153 = btb_pc_28 == io_if_pc; // @[BTB.scala 70:42:@389.4]
  assign _T_154 = btb_pc_29 == io_if_pc; // @[BTB.scala 70:42:@390.4]
  assign _T_155 = btb_pc_30 == io_if_pc; // @[BTB.scala 70:42:@391.4]
  assign _T_156 = btb_pc_31 == io_if_pc; // @[BTB.scala 70:42:@392.4]
  assign _T_157 = btb_pc_32 == io_if_pc; // @[BTB.scala 70:42:@393.4]
  assign _T_158 = btb_pc_33 == io_if_pc; // @[BTB.scala 70:42:@394.4]
  assign _T_159 = btb_pc_34 == io_if_pc; // @[BTB.scala 70:42:@395.4]
  assign _T_160 = btb_pc_35 == io_if_pc; // @[BTB.scala 70:42:@396.4]
  assign _T_161 = btb_pc_36 == io_if_pc; // @[BTB.scala 70:42:@397.4]
  assign _T_162 = btb_pc_37 == io_if_pc; // @[BTB.scala 70:42:@398.4]
  assign _T_163 = btb_pc_38 == io_if_pc; // @[BTB.scala 70:42:@399.4]
  assign _T_164 = btb_pc_39 == io_if_pc; // @[BTB.scala 70:42:@400.4]
  assign _T_165 = btb_pc_40 == io_if_pc; // @[BTB.scala 70:42:@401.4]
  assign _T_166 = btb_pc_41 == io_if_pc; // @[BTB.scala 70:42:@402.4]
  assign _T_167 = btb_pc_42 == io_if_pc; // @[BTB.scala 70:42:@403.4]
  assign _T_168 = btb_pc_43 == io_if_pc; // @[BTB.scala 70:42:@404.4]
  assign _T_169 = btb_pc_44 == io_if_pc; // @[BTB.scala 70:42:@405.4]
  assign _T_170 = btb_pc_45 == io_if_pc; // @[BTB.scala 70:42:@406.4]
  assign _T_171 = btb_pc_46 == io_if_pc; // @[BTB.scala 70:42:@407.4]
  assign _T_172 = btb_pc_47 == io_if_pc; // @[BTB.scala 70:42:@408.4]
  assign _T_173 = btb_pc_48 == io_if_pc; // @[BTB.scala 70:42:@409.4]
  assign _T_174 = btb_pc_49 == io_if_pc; // @[BTB.scala 70:42:@410.4]
  assign _T_175 = btb_pc_50 == io_if_pc; // @[BTB.scala 70:42:@411.4]
  assign _T_176 = btb_pc_51 == io_if_pc; // @[BTB.scala 70:42:@412.4]
  assign _T_177 = btb_pc_52 == io_if_pc; // @[BTB.scala 70:42:@413.4]
  assign _T_178 = btb_pc_53 == io_if_pc; // @[BTB.scala 70:42:@414.4]
  assign _T_179 = btb_pc_54 == io_if_pc; // @[BTB.scala 70:42:@415.4]
  assign _T_180 = btb_pc_55 == io_if_pc; // @[BTB.scala 70:42:@416.4]
  assign _T_181 = btb_pc_56 == io_if_pc; // @[BTB.scala 70:42:@417.4]
  assign _T_182 = btb_pc_57 == io_if_pc; // @[BTB.scala 70:42:@418.4]
  assign _T_183 = btb_pc_58 == io_if_pc; // @[BTB.scala 70:42:@419.4]
  assign _T_184 = btb_pc_59 == io_if_pc; // @[BTB.scala 70:42:@420.4]
  assign _T_185 = btb_pc_60 == io_if_pc; // @[BTB.scala 70:42:@421.4]
  assign _T_186 = btb_pc_61 == io_if_pc; // @[BTB.scala 70:42:@422.4]
  assign _T_187 = btb_pc_62 == io_if_pc; // @[BTB.scala 70:42:@423.4]
  assign _T_188 = btb_pc_63 == io_if_pc; // @[BTB.scala 70:42:@424.4]
  assign _T_265 = {_T_132,_T_131,_T_130,_T_129,_T_128,_T_127,_T_126,_T_125}; // @[BTB.scala 70:57:@496.4]
  assign _T_273 = {_T_140,_T_139,_T_138,_T_137,_T_136,_T_135,_T_134,_T_133,_T_265}; // @[BTB.scala 70:57:@504.4]
  assign _T_280 = {_T_148,_T_147,_T_146,_T_145,_T_144,_T_143,_T_142,_T_141}; // @[BTB.scala 70:57:@511.4]
  assign _T_289 = {_T_156,_T_155,_T_154,_T_153,_T_152,_T_151,_T_150,_T_149,_T_280,_T_273}; // @[BTB.scala 70:57:@520.4]
  assign _T_296 = {_T_164,_T_163,_T_162,_T_161,_T_160,_T_159,_T_158,_T_157}; // @[BTB.scala 70:57:@527.4]
  assign _T_304 = {_T_172,_T_171,_T_170,_T_169,_T_168,_T_167,_T_166,_T_165,_T_296}; // @[BTB.scala 70:57:@535.4]
  assign _T_311 = {_T_180,_T_179,_T_178,_T_177,_T_176,_T_175,_T_174,_T_173}; // @[BTB.scala 70:57:@542.4]
  assign _T_320 = {_T_188,_T_187,_T_186,_T_185,_T_184,_T_183,_T_182,_T_181,_T_311,_T_304}; // @[BTB.scala 70:57:@551.4]
  assign _T_321 = {_T_320,_T_289}; // @[BTB.scala 70:57:@552.4]
  assign _T_323 = btb_btype_0 != 2'h0; // @[BTB.scala 50:66:@553.4]
  assign _T_325 = btb_btype_1 != 2'h0; // @[BTB.scala 50:66:@554.4]
  assign _T_327 = btb_btype_2 != 2'h0; // @[BTB.scala 50:66:@555.4]
  assign _T_329 = btb_btype_3 != 2'h0; // @[BTB.scala 50:66:@556.4]
  assign _T_331 = btb_btype_4 != 2'h0; // @[BTB.scala 50:66:@557.4]
  assign _T_333 = btb_btype_5 != 2'h0; // @[BTB.scala 50:66:@558.4]
  assign _T_335 = btb_btype_6 != 2'h0; // @[BTB.scala 50:66:@559.4]
  assign _T_337 = btb_btype_7 != 2'h0; // @[BTB.scala 50:66:@560.4]
  assign _T_339 = btb_btype_8 != 2'h0; // @[BTB.scala 50:66:@561.4]
  assign _T_341 = btb_btype_9 != 2'h0; // @[BTB.scala 50:66:@562.4]
  assign _T_343 = btb_btype_10 != 2'h0; // @[BTB.scala 50:66:@563.4]
  assign _T_345 = btb_btype_11 != 2'h0; // @[BTB.scala 50:66:@564.4]
  assign _T_347 = btb_btype_12 != 2'h0; // @[BTB.scala 50:66:@565.4]
  assign _T_349 = btb_btype_13 != 2'h0; // @[BTB.scala 50:66:@566.4]
  assign _T_351 = btb_btype_14 != 2'h0; // @[BTB.scala 50:66:@567.4]
  assign _T_353 = btb_btype_15 != 2'h0; // @[BTB.scala 50:66:@568.4]
  assign _T_355 = btb_btype_16 != 2'h0; // @[BTB.scala 50:66:@569.4]
  assign _T_357 = btb_btype_17 != 2'h0; // @[BTB.scala 50:66:@570.4]
  assign _T_359 = btb_btype_18 != 2'h0; // @[BTB.scala 50:66:@571.4]
  assign _T_361 = btb_btype_19 != 2'h0; // @[BTB.scala 50:66:@572.4]
  assign _T_363 = btb_btype_20 != 2'h0; // @[BTB.scala 50:66:@573.4]
  assign _T_365 = btb_btype_21 != 2'h0; // @[BTB.scala 50:66:@574.4]
  assign _T_367 = btb_btype_22 != 2'h0; // @[BTB.scala 50:66:@575.4]
  assign _T_369 = btb_btype_23 != 2'h0; // @[BTB.scala 50:66:@576.4]
  assign _T_371 = btb_btype_24 != 2'h0; // @[BTB.scala 50:66:@577.4]
  assign _T_373 = btb_btype_25 != 2'h0; // @[BTB.scala 50:66:@578.4]
  assign _T_375 = btb_btype_26 != 2'h0; // @[BTB.scala 50:66:@579.4]
  assign _T_377 = btb_btype_27 != 2'h0; // @[BTB.scala 50:66:@580.4]
  assign _T_379 = btb_btype_28 != 2'h0; // @[BTB.scala 50:66:@581.4]
  assign _T_381 = btb_btype_29 != 2'h0; // @[BTB.scala 50:66:@582.4]
  assign _T_383 = btb_btype_30 != 2'h0; // @[BTB.scala 50:66:@583.4]
  assign _T_385 = btb_btype_31 != 2'h0; // @[BTB.scala 50:66:@584.4]
  assign _T_387 = btb_btype_32 != 2'h0; // @[BTB.scala 50:66:@585.4]
  assign _T_389 = btb_btype_33 != 2'h0; // @[BTB.scala 50:66:@586.4]
  assign _T_391 = btb_btype_34 != 2'h0; // @[BTB.scala 50:66:@587.4]
  assign _T_393 = btb_btype_35 != 2'h0; // @[BTB.scala 50:66:@588.4]
  assign _T_395 = btb_btype_36 != 2'h0; // @[BTB.scala 50:66:@589.4]
  assign _T_397 = btb_btype_37 != 2'h0; // @[BTB.scala 50:66:@590.4]
  assign _T_399 = btb_btype_38 != 2'h0; // @[BTB.scala 50:66:@591.4]
  assign _T_401 = btb_btype_39 != 2'h0; // @[BTB.scala 50:66:@592.4]
  assign _T_403 = btb_btype_40 != 2'h0; // @[BTB.scala 50:66:@593.4]
  assign _T_405 = btb_btype_41 != 2'h0; // @[BTB.scala 50:66:@594.4]
  assign _T_407 = btb_btype_42 != 2'h0; // @[BTB.scala 50:66:@595.4]
  assign _T_409 = btb_btype_43 != 2'h0; // @[BTB.scala 50:66:@596.4]
  assign _T_411 = btb_btype_44 != 2'h0; // @[BTB.scala 50:66:@597.4]
  assign _T_413 = btb_btype_45 != 2'h0; // @[BTB.scala 50:66:@598.4]
  assign _T_415 = btb_btype_46 != 2'h0; // @[BTB.scala 50:66:@599.4]
  assign _T_417 = btb_btype_47 != 2'h0; // @[BTB.scala 50:66:@600.4]
  assign _T_419 = btb_btype_48 != 2'h0; // @[BTB.scala 50:66:@601.4]
  assign _T_421 = btb_btype_49 != 2'h0; // @[BTB.scala 50:66:@602.4]
  assign _T_423 = btb_btype_50 != 2'h0; // @[BTB.scala 50:66:@603.4]
  assign _T_425 = btb_btype_51 != 2'h0; // @[BTB.scala 50:66:@604.4]
  assign _T_427 = btb_btype_52 != 2'h0; // @[BTB.scala 50:66:@605.4]
  assign _T_429 = btb_btype_53 != 2'h0; // @[BTB.scala 50:66:@606.4]
  assign _T_431 = btb_btype_54 != 2'h0; // @[BTB.scala 50:66:@607.4]
  assign _T_433 = btb_btype_55 != 2'h0; // @[BTB.scala 50:66:@608.4]
  assign _T_435 = btb_btype_56 != 2'h0; // @[BTB.scala 50:66:@609.4]
  assign _T_437 = btb_btype_57 != 2'h0; // @[BTB.scala 50:66:@610.4]
  assign _T_439 = btb_btype_58 != 2'h0; // @[BTB.scala 50:66:@611.4]
  assign _T_441 = btb_btype_59 != 2'h0; // @[BTB.scala 50:66:@612.4]
  assign _T_443 = btb_btype_60 != 2'h0; // @[BTB.scala 50:66:@613.4]
  assign _T_445 = btb_btype_61 != 2'h0; // @[BTB.scala 50:66:@614.4]
  assign _T_447 = btb_btype_62 != 2'h0; // @[BTB.scala 50:66:@615.4]
  assign _T_449 = btb_btype_63 != 2'h0; // @[BTB.scala 50:66:@616.4]
  assign _T_526 = {_T_337,_T_335,_T_333,_T_331,_T_329,_T_327,_T_325,_T_323}; // @[BTB.scala 50:72:@688.4]
  assign _T_534 = {_T_353,_T_351,_T_349,_T_347,_T_345,_T_343,_T_341,_T_339,_T_526}; // @[BTB.scala 50:72:@696.4]
  assign _T_541 = {_T_369,_T_367,_T_365,_T_363,_T_361,_T_359,_T_357,_T_355}; // @[BTB.scala 50:72:@703.4]
  assign _T_550 = {_T_385,_T_383,_T_381,_T_379,_T_377,_T_375,_T_373,_T_371,_T_541,_T_534}; // @[BTB.scala 50:72:@712.4]
  assign _T_557 = {_T_401,_T_399,_T_397,_T_395,_T_393,_T_391,_T_389,_T_387}; // @[BTB.scala 50:72:@719.4]
  assign _T_565 = {_T_417,_T_415,_T_413,_T_411,_T_409,_T_407,_T_405,_T_403,_T_557}; // @[BTB.scala 50:72:@727.4]
  assign _T_572 = {_T_433,_T_431,_T_429,_T_427,_T_425,_T_423,_T_421,_T_419}; // @[BTB.scala 50:72:@734.4]
  assign _T_581 = {_T_449,_T_447,_T_445,_T_443,_T_441,_T_439,_T_437,_T_435,_T_572,_T_565}; // @[BTB.scala 50:72:@743.4]
  assign _T_582 = {_T_581,_T_550}; // @[BTB.scala 50:72:@744.4]
  assign predict_lookup = _T_321 & _T_582; // @[BTB.scala 70:64:@745.4]
  assign _T_585 = io_if_pc + 32'h4; // @[BTB.scala 71:32:@747.4]
  assign predict_cont_tgt = io_if_pc + 32'h4; // @[BTB.scala 71:32:@748.4]
  assign _T_587 = predict_lookup[0]; // @[Mux.scala 21:36:@750.4]
  assign _T_588 = predict_lookup[1]; // @[Mux.scala 21:36:@751.4]
  assign _T_589 = predict_lookup[2]; // @[Mux.scala 21:36:@752.4]
  assign _T_590 = predict_lookup[3]; // @[Mux.scala 21:36:@753.4]
  assign _T_591 = predict_lookup[4]; // @[Mux.scala 21:36:@754.4]
  assign _T_592 = predict_lookup[5]; // @[Mux.scala 21:36:@755.4]
  assign _T_593 = predict_lookup[6]; // @[Mux.scala 21:36:@756.4]
  assign _T_594 = predict_lookup[7]; // @[Mux.scala 21:36:@757.4]
  assign _T_595 = predict_lookup[8]; // @[Mux.scala 21:36:@758.4]
  assign _T_596 = predict_lookup[9]; // @[Mux.scala 21:36:@759.4]
  assign _T_597 = predict_lookup[10]; // @[Mux.scala 21:36:@760.4]
  assign _T_598 = predict_lookup[11]; // @[Mux.scala 21:36:@761.4]
  assign _T_599 = predict_lookup[12]; // @[Mux.scala 21:36:@762.4]
  assign _T_600 = predict_lookup[13]; // @[Mux.scala 21:36:@763.4]
  assign _T_601 = predict_lookup[14]; // @[Mux.scala 21:36:@764.4]
  assign _T_602 = predict_lookup[15]; // @[Mux.scala 21:36:@765.4]
  assign _T_603 = predict_lookup[16]; // @[Mux.scala 21:36:@766.4]
  assign _T_604 = predict_lookup[17]; // @[Mux.scala 21:36:@767.4]
  assign _T_605 = predict_lookup[18]; // @[Mux.scala 21:36:@768.4]
  assign _T_606 = predict_lookup[19]; // @[Mux.scala 21:36:@769.4]
  assign _T_607 = predict_lookup[20]; // @[Mux.scala 21:36:@770.4]
  assign _T_608 = predict_lookup[21]; // @[Mux.scala 21:36:@771.4]
  assign _T_609 = predict_lookup[22]; // @[Mux.scala 21:36:@772.4]
  assign _T_610 = predict_lookup[23]; // @[Mux.scala 21:36:@773.4]
  assign _T_611 = predict_lookup[24]; // @[Mux.scala 21:36:@774.4]
  assign _T_612 = predict_lookup[25]; // @[Mux.scala 21:36:@775.4]
  assign _T_613 = predict_lookup[26]; // @[Mux.scala 21:36:@776.4]
  assign _T_614 = predict_lookup[27]; // @[Mux.scala 21:36:@777.4]
  assign _T_615 = predict_lookup[28]; // @[Mux.scala 21:36:@778.4]
  assign _T_616 = predict_lookup[29]; // @[Mux.scala 21:36:@779.4]
  assign _T_617 = predict_lookup[30]; // @[Mux.scala 21:36:@780.4]
  assign _T_618 = predict_lookup[31]; // @[Mux.scala 21:36:@781.4]
  assign _T_619 = predict_lookup[32]; // @[Mux.scala 21:36:@782.4]
  assign _T_620 = predict_lookup[33]; // @[Mux.scala 21:36:@783.4]
  assign _T_621 = predict_lookup[34]; // @[Mux.scala 21:36:@784.4]
  assign _T_622 = predict_lookup[35]; // @[Mux.scala 21:36:@785.4]
  assign _T_623 = predict_lookup[36]; // @[Mux.scala 21:36:@786.4]
  assign _T_624 = predict_lookup[37]; // @[Mux.scala 21:36:@787.4]
  assign _T_625 = predict_lookup[38]; // @[Mux.scala 21:36:@788.4]
  assign _T_626 = predict_lookup[39]; // @[Mux.scala 21:36:@789.4]
  assign _T_627 = predict_lookup[40]; // @[Mux.scala 21:36:@790.4]
  assign _T_628 = predict_lookup[41]; // @[Mux.scala 21:36:@791.4]
  assign _T_629 = predict_lookup[42]; // @[Mux.scala 21:36:@792.4]
  assign _T_630 = predict_lookup[43]; // @[Mux.scala 21:36:@793.4]
  assign _T_631 = predict_lookup[44]; // @[Mux.scala 21:36:@794.4]
  assign _T_632 = predict_lookup[45]; // @[Mux.scala 21:36:@795.4]
  assign _T_633 = predict_lookup[46]; // @[Mux.scala 21:36:@796.4]
  assign _T_634 = predict_lookup[47]; // @[Mux.scala 21:36:@797.4]
  assign _T_635 = predict_lookup[48]; // @[Mux.scala 21:36:@798.4]
  assign _T_636 = predict_lookup[49]; // @[Mux.scala 21:36:@799.4]
  assign _T_637 = predict_lookup[50]; // @[Mux.scala 21:36:@800.4]
  assign _T_638 = predict_lookup[51]; // @[Mux.scala 21:36:@801.4]
  assign _T_639 = predict_lookup[52]; // @[Mux.scala 21:36:@802.4]
  assign _T_640 = predict_lookup[53]; // @[Mux.scala 21:36:@803.4]
  assign _T_641 = predict_lookup[54]; // @[Mux.scala 21:36:@804.4]
  assign _T_642 = predict_lookup[55]; // @[Mux.scala 21:36:@805.4]
  assign _T_643 = predict_lookup[56]; // @[Mux.scala 21:36:@806.4]
  assign _T_644 = predict_lookup[57]; // @[Mux.scala 21:36:@807.4]
  assign _T_645 = predict_lookup[58]; // @[Mux.scala 21:36:@808.4]
  assign _T_646 = predict_lookup[59]; // @[Mux.scala 21:36:@809.4]
  assign _T_647 = predict_lookup[60]; // @[Mux.scala 21:36:@810.4]
  assign _T_648 = predict_lookup[61]; // @[Mux.scala 21:36:@811.4]
  assign _T_649 = predict_lookup[62]; // @[Mux.scala 21:36:@812.4]
  assign _T_650 = predict_lookup[63]; // @[Mux.scala 21:36:@813.4]
  assign _T_653 = _T_587 ? btb_target_0 : 32'h0; // @[Mux.scala 19:72:@814.4]
  assign _T_655 = _T_588 ? btb_target_1 : 32'h0; // @[Mux.scala 19:72:@815.4]
  assign _T_657 = _T_589 ? btb_target_2 : 32'h0; // @[Mux.scala 19:72:@816.4]
  assign _T_659 = _T_590 ? btb_target_3 : 32'h0; // @[Mux.scala 19:72:@817.4]
  assign _T_661 = _T_591 ? btb_target_4 : 32'h0; // @[Mux.scala 19:72:@818.4]
  assign _T_663 = _T_592 ? btb_target_5 : 32'h0; // @[Mux.scala 19:72:@819.4]
  assign _T_665 = _T_593 ? btb_target_6 : 32'h0; // @[Mux.scala 19:72:@820.4]
  assign _T_667 = _T_594 ? btb_target_7 : 32'h0; // @[Mux.scala 19:72:@821.4]
  assign _T_669 = _T_595 ? btb_target_8 : 32'h0; // @[Mux.scala 19:72:@822.4]
  assign _T_671 = _T_596 ? btb_target_9 : 32'h0; // @[Mux.scala 19:72:@823.4]
  assign _T_673 = _T_597 ? btb_target_10 : 32'h0; // @[Mux.scala 19:72:@824.4]
  assign _T_675 = _T_598 ? btb_target_11 : 32'h0; // @[Mux.scala 19:72:@825.4]
  assign _T_677 = _T_599 ? btb_target_12 : 32'h0; // @[Mux.scala 19:72:@826.4]
  assign _T_679 = _T_600 ? btb_target_13 : 32'h0; // @[Mux.scala 19:72:@827.4]
  assign _T_681 = _T_601 ? btb_target_14 : 32'h0; // @[Mux.scala 19:72:@828.4]
  assign _T_683 = _T_602 ? btb_target_15 : 32'h0; // @[Mux.scala 19:72:@829.4]
  assign _T_685 = _T_603 ? btb_target_16 : 32'h0; // @[Mux.scala 19:72:@830.4]
  assign _T_687 = _T_604 ? btb_target_17 : 32'h0; // @[Mux.scala 19:72:@831.4]
  assign _T_689 = _T_605 ? btb_target_18 : 32'h0; // @[Mux.scala 19:72:@832.4]
  assign _T_691 = _T_606 ? btb_target_19 : 32'h0; // @[Mux.scala 19:72:@833.4]
  assign _T_693 = _T_607 ? btb_target_20 : 32'h0; // @[Mux.scala 19:72:@834.4]
  assign _T_695 = _T_608 ? btb_target_21 : 32'h0; // @[Mux.scala 19:72:@835.4]
  assign _T_697 = _T_609 ? btb_target_22 : 32'h0; // @[Mux.scala 19:72:@836.4]
  assign _T_699 = _T_610 ? btb_target_23 : 32'h0; // @[Mux.scala 19:72:@837.4]
  assign _T_701 = _T_611 ? btb_target_24 : 32'h0; // @[Mux.scala 19:72:@838.4]
  assign _T_703 = _T_612 ? btb_target_25 : 32'h0; // @[Mux.scala 19:72:@839.4]
  assign _T_705 = _T_613 ? btb_target_26 : 32'h0; // @[Mux.scala 19:72:@840.4]
  assign _T_707 = _T_614 ? btb_target_27 : 32'h0; // @[Mux.scala 19:72:@841.4]
  assign _T_709 = _T_615 ? btb_target_28 : 32'h0; // @[Mux.scala 19:72:@842.4]
  assign _T_711 = _T_616 ? btb_target_29 : 32'h0; // @[Mux.scala 19:72:@843.4]
  assign _T_713 = _T_617 ? btb_target_30 : 32'h0; // @[Mux.scala 19:72:@844.4]
  assign _T_715 = _T_618 ? btb_target_31 : 32'h0; // @[Mux.scala 19:72:@845.4]
  assign _T_717 = _T_619 ? btb_target_32 : 32'h0; // @[Mux.scala 19:72:@846.4]
  assign _T_719 = _T_620 ? btb_target_33 : 32'h0; // @[Mux.scala 19:72:@847.4]
  assign _T_721 = _T_621 ? btb_target_34 : 32'h0; // @[Mux.scala 19:72:@848.4]
  assign _T_723 = _T_622 ? btb_target_35 : 32'h0; // @[Mux.scala 19:72:@849.4]
  assign _T_725 = _T_623 ? btb_target_36 : 32'h0; // @[Mux.scala 19:72:@850.4]
  assign _T_727 = _T_624 ? btb_target_37 : 32'h0; // @[Mux.scala 19:72:@851.4]
  assign _T_729 = _T_625 ? btb_target_38 : 32'h0; // @[Mux.scala 19:72:@852.4]
  assign _T_731 = _T_626 ? btb_target_39 : 32'h0; // @[Mux.scala 19:72:@853.4]
  assign _T_733 = _T_627 ? btb_target_40 : 32'h0; // @[Mux.scala 19:72:@854.4]
  assign _T_735 = _T_628 ? btb_target_41 : 32'h0; // @[Mux.scala 19:72:@855.4]
  assign _T_737 = _T_629 ? btb_target_42 : 32'h0; // @[Mux.scala 19:72:@856.4]
  assign _T_739 = _T_630 ? btb_target_43 : 32'h0; // @[Mux.scala 19:72:@857.4]
  assign _T_741 = _T_631 ? btb_target_44 : 32'h0; // @[Mux.scala 19:72:@858.4]
  assign _T_743 = _T_632 ? btb_target_45 : 32'h0; // @[Mux.scala 19:72:@859.4]
  assign _T_745 = _T_633 ? btb_target_46 : 32'h0; // @[Mux.scala 19:72:@860.4]
  assign _T_747 = _T_634 ? btb_target_47 : 32'h0; // @[Mux.scala 19:72:@861.4]
  assign _T_749 = _T_635 ? btb_target_48 : 32'h0; // @[Mux.scala 19:72:@862.4]
  assign _T_751 = _T_636 ? btb_target_49 : 32'h0; // @[Mux.scala 19:72:@863.4]
  assign _T_753 = _T_637 ? btb_target_50 : 32'h0; // @[Mux.scala 19:72:@864.4]
  assign _T_755 = _T_638 ? btb_target_51 : 32'h0; // @[Mux.scala 19:72:@865.4]
  assign _T_757 = _T_639 ? btb_target_52 : 32'h0; // @[Mux.scala 19:72:@866.4]
  assign _T_759 = _T_640 ? btb_target_53 : 32'h0; // @[Mux.scala 19:72:@867.4]
  assign _T_761 = _T_641 ? btb_target_54 : 32'h0; // @[Mux.scala 19:72:@868.4]
  assign _T_763 = _T_642 ? btb_target_55 : 32'h0; // @[Mux.scala 19:72:@869.4]
  assign _T_765 = _T_643 ? btb_target_56 : 32'h0; // @[Mux.scala 19:72:@870.4]
  assign _T_767 = _T_644 ? btb_target_57 : 32'h0; // @[Mux.scala 19:72:@871.4]
  assign _T_769 = _T_645 ? btb_target_58 : 32'h0; // @[Mux.scala 19:72:@872.4]
  assign _T_771 = _T_646 ? btb_target_59 : 32'h0; // @[Mux.scala 19:72:@873.4]
  assign _T_773 = _T_647 ? btb_target_60 : 32'h0; // @[Mux.scala 19:72:@874.4]
  assign _T_775 = _T_648 ? btb_target_61 : 32'h0; // @[Mux.scala 19:72:@875.4]
  assign _T_777 = _T_649 ? btb_target_62 : 32'h0; // @[Mux.scala 19:72:@876.4]
  assign _T_779 = _T_650 ? btb_target_63 : 32'h0; // @[Mux.scala 19:72:@877.4]
  assign _T_780 = _T_653 | _T_655; // @[Mux.scala 19:72:@878.4]
  assign _T_781 = _T_780 | _T_657; // @[Mux.scala 19:72:@879.4]
  assign _T_782 = _T_781 | _T_659; // @[Mux.scala 19:72:@880.4]
  assign _T_783 = _T_782 | _T_661; // @[Mux.scala 19:72:@881.4]
  assign _T_784 = _T_783 | _T_663; // @[Mux.scala 19:72:@882.4]
  assign _T_785 = _T_784 | _T_665; // @[Mux.scala 19:72:@883.4]
  assign _T_786 = _T_785 | _T_667; // @[Mux.scala 19:72:@884.4]
  assign _T_787 = _T_786 | _T_669; // @[Mux.scala 19:72:@885.4]
  assign _T_788 = _T_787 | _T_671; // @[Mux.scala 19:72:@886.4]
  assign _T_789 = _T_788 | _T_673; // @[Mux.scala 19:72:@887.4]
  assign _T_790 = _T_789 | _T_675; // @[Mux.scala 19:72:@888.4]
  assign _T_791 = _T_790 | _T_677; // @[Mux.scala 19:72:@889.4]
  assign _T_792 = _T_791 | _T_679; // @[Mux.scala 19:72:@890.4]
  assign _T_793 = _T_792 | _T_681; // @[Mux.scala 19:72:@891.4]
  assign _T_794 = _T_793 | _T_683; // @[Mux.scala 19:72:@892.4]
  assign _T_795 = _T_794 | _T_685; // @[Mux.scala 19:72:@893.4]
  assign _T_796 = _T_795 | _T_687; // @[Mux.scala 19:72:@894.4]
  assign _T_797 = _T_796 | _T_689; // @[Mux.scala 19:72:@895.4]
  assign _T_798 = _T_797 | _T_691; // @[Mux.scala 19:72:@896.4]
  assign _T_799 = _T_798 | _T_693; // @[Mux.scala 19:72:@897.4]
  assign _T_800 = _T_799 | _T_695; // @[Mux.scala 19:72:@898.4]
  assign _T_801 = _T_800 | _T_697; // @[Mux.scala 19:72:@899.4]
  assign _T_802 = _T_801 | _T_699; // @[Mux.scala 19:72:@900.4]
  assign _T_803 = _T_802 | _T_701; // @[Mux.scala 19:72:@901.4]
  assign _T_804 = _T_803 | _T_703; // @[Mux.scala 19:72:@902.4]
  assign _T_805 = _T_804 | _T_705; // @[Mux.scala 19:72:@903.4]
  assign _T_806 = _T_805 | _T_707; // @[Mux.scala 19:72:@904.4]
  assign _T_807 = _T_806 | _T_709; // @[Mux.scala 19:72:@905.4]
  assign _T_808 = _T_807 | _T_711; // @[Mux.scala 19:72:@906.4]
  assign _T_809 = _T_808 | _T_713; // @[Mux.scala 19:72:@907.4]
  assign _T_810 = _T_809 | _T_715; // @[Mux.scala 19:72:@908.4]
  assign _T_811 = _T_810 | _T_717; // @[Mux.scala 19:72:@909.4]
  assign _T_812 = _T_811 | _T_719; // @[Mux.scala 19:72:@910.4]
  assign _T_813 = _T_812 | _T_721; // @[Mux.scala 19:72:@911.4]
  assign _T_814 = _T_813 | _T_723; // @[Mux.scala 19:72:@912.4]
  assign _T_815 = _T_814 | _T_725; // @[Mux.scala 19:72:@913.4]
  assign _T_816 = _T_815 | _T_727; // @[Mux.scala 19:72:@914.4]
  assign _T_817 = _T_816 | _T_729; // @[Mux.scala 19:72:@915.4]
  assign _T_818 = _T_817 | _T_731; // @[Mux.scala 19:72:@916.4]
  assign _T_819 = _T_818 | _T_733; // @[Mux.scala 19:72:@917.4]
  assign _T_820 = _T_819 | _T_735; // @[Mux.scala 19:72:@918.4]
  assign _T_821 = _T_820 | _T_737; // @[Mux.scala 19:72:@919.4]
  assign _T_822 = _T_821 | _T_739; // @[Mux.scala 19:72:@920.4]
  assign _T_823 = _T_822 | _T_741; // @[Mux.scala 19:72:@921.4]
  assign _T_824 = _T_823 | _T_743; // @[Mux.scala 19:72:@922.4]
  assign _T_825 = _T_824 | _T_745; // @[Mux.scala 19:72:@923.4]
  assign _T_826 = _T_825 | _T_747; // @[Mux.scala 19:72:@924.4]
  assign _T_827 = _T_826 | _T_749; // @[Mux.scala 19:72:@925.4]
  assign _T_828 = _T_827 | _T_751; // @[Mux.scala 19:72:@926.4]
  assign _T_829 = _T_828 | _T_753; // @[Mux.scala 19:72:@927.4]
  assign _T_830 = _T_829 | _T_755; // @[Mux.scala 19:72:@928.4]
  assign _T_831 = _T_830 | _T_757; // @[Mux.scala 19:72:@929.4]
  assign _T_832 = _T_831 | _T_759; // @[Mux.scala 19:72:@930.4]
  assign _T_833 = _T_832 | _T_761; // @[Mux.scala 19:72:@931.4]
  assign _T_834 = _T_833 | _T_763; // @[Mux.scala 19:72:@932.4]
  assign _T_835 = _T_834 | _T_765; // @[Mux.scala 19:72:@933.4]
  assign _T_836 = _T_835 | _T_767; // @[Mux.scala 19:72:@934.4]
  assign _T_837 = _T_836 | _T_769; // @[Mux.scala 19:72:@935.4]
  assign _T_838 = _T_837 | _T_771; // @[Mux.scala 19:72:@936.4]
  assign _T_839 = _T_838 | _T_773; // @[Mux.scala 19:72:@937.4]
  assign _T_840 = _T_839 | _T_775; // @[Mux.scala 19:72:@938.4]
  assign _T_841 = _T_840 | _T_777; // @[Mux.scala 19:72:@939.4]
  assign predict_jump_tgt = _T_841 | _T_779; // @[Mux.scala 19:72:@940.4]
  assign _T_911 = _T_587 ? btb_btype_0 : 2'h0; // @[Mux.scala 19:72:@1008.4]
  assign _T_913 = _T_588 ? btb_btype_1 : 2'h0; // @[Mux.scala 19:72:@1009.4]
  assign _T_915 = _T_589 ? btb_btype_2 : 2'h0; // @[Mux.scala 19:72:@1010.4]
  assign _T_917 = _T_590 ? btb_btype_3 : 2'h0; // @[Mux.scala 19:72:@1011.4]
  assign _T_919 = _T_591 ? btb_btype_4 : 2'h0; // @[Mux.scala 19:72:@1012.4]
  assign _T_921 = _T_592 ? btb_btype_5 : 2'h0; // @[Mux.scala 19:72:@1013.4]
  assign _T_923 = _T_593 ? btb_btype_6 : 2'h0; // @[Mux.scala 19:72:@1014.4]
  assign _T_925 = _T_594 ? btb_btype_7 : 2'h0; // @[Mux.scala 19:72:@1015.4]
  assign _T_927 = _T_595 ? btb_btype_8 : 2'h0; // @[Mux.scala 19:72:@1016.4]
  assign _T_929 = _T_596 ? btb_btype_9 : 2'h0; // @[Mux.scala 19:72:@1017.4]
  assign _T_931 = _T_597 ? btb_btype_10 : 2'h0; // @[Mux.scala 19:72:@1018.4]
  assign _T_933 = _T_598 ? btb_btype_11 : 2'h0; // @[Mux.scala 19:72:@1019.4]
  assign _T_935 = _T_599 ? btb_btype_12 : 2'h0; // @[Mux.scala 19:72:@1020.4]
  assign _T_937 = _T_600 ? btb_btype_13 : 2'h0; // @[Mux.scala 19:72:@1021.4]
  assign _T_939 = _T_601 ? btb_btype_14 : 2'h0; // @[Mux.scala 19:72:@1022.4]
  assign _T_941 = _T_602 ? btb_btype_15 : 2'h0; // @[Mux.scala 19:72:@1023.4]
  assign _T_943 = _T_603 ? btb_btype_16 : 2'h0; // @[Mux.scala 19:72:@1024.4]
  assign _T_945 = _T_604 ? btb_btype_17 : 2'h0; // @[Mux.scala 19:72:@1025.4]
  assign _T_947 = _T_605 ? btb_btype_18 : 2'h0; // @[Mux.scala 19:72:@1026.4]
  assign _T_949 = _T_606 ? btb_btype_19 : 2'h0; // @[Mux.scala 19:72:@1027.4]
  assign _T_951 = _T_607 ? btb_btype_20 : 2'h0; // @[Mux.scala 19:72:@1028.4]
  assign _T_953 = _T_608 ? btb_btype_21 : 2'h0; // @[Mux.scala 19:72:@1029.4]
  assign _T_955 = _T_609 ? btb_btype_22 : 2'h0; // @[Mux.scala 19:72:@1030.4]
  assign _T_957 = _T_610 ? btb_btype_23 : 2'h0; // @[Mux.scala 19:72:@1031.4]
  assign _T_959 = _T_611 ? btb_btype_24 : 2'h0; // @[Mux.scala 19:72:@1032.4]
  assign _T_961 = _T_612 ? btb_btype_25 : 2'h0; // @[Mux.scala 19:72:@1033.4]
  assign _T_963 = _T_613 ? btb_btype_26 : 2'h0; // @[Mux.scala 19:72:@1034.4]
  assign _T_965 = _T_614 ? btb_btype_27 : 2'h0; // @[Mux.scala 19:72:@1035.4]
  assign _T_967 = _T_615 ? btb_btype_28 : 2'h0; // @[Mux.scala 19:72:@1036.4]
  assign _T_969 = _T_616 ? btb_btype_29 : 2'h0; // @[Mux.scala 19:72:@1037.4]
  assign _T_971 = _T_617 ? btb_btype_30 : 2'h0; // @[Mux.scala 19:72:@1038.4]
  assign _T_973 = _T_618 ? btb_btype_31 : 2'h0; // @[Mux.scala 19:72:@1039.4]
  assign _T_975 = _T_619 ? btb_btype_32 : 2'h0; // @[Mux.scala 19:72:@1040.4]
  assign _T_977 = _T_620 ? btb_btype_33 : 2'h0; // @[Mux.scala 19:72:@1041.4]
  assign _T_979 = _T_621 ? btb_btype_34 : 2'h0; // @[Mux.scala 19:72:@1042.4]
  assign _T_981 = _T_622 ? btb_btype_35 : 2'h0; // @[Mux.scala 19:72:@1043.4]
  assign _T_983 = _T_623 ? btb_btype_36 : 2'h0; // @[Mux.scala 19:72:@1044.4]
  assign _T_985 = _T_624 ? btb_btype_37 : 2'h0; // @[Mux.scala 19:72:@1045.4]
  assign _T_987 = _T_625 ? btb_btype_38 : 2'h0; // @[Mux.scala 19:72:@1046.4]
  assign _T_989 = _T_626 ? btb_btype_39 : 2'h0; // @[Mux.scala 19:72:@1047.4]
  assign _T_991 = _T_627 ? btb_btype_40 : 2'h0; // @[Mux.scala 19:72:@1048.4]
  assign _T_993 = _T_628 ? btb_btype_41 : 2'h0; // @[Mux.scala 19:72:@1049.4]
  assign _T_995 = _T_629 ? btb_btype_42 : 2'h0; // @[Mux.scala 19:72:@1050.4]
  assign _T_997 = _T_630 ? btb_btype_43 : 2'h0; // @[Mux.scala 19:72:@1051.4]
  assign _T_999 = _T_631 ? btb_btype_44 : 2'h0; // @[Mux.scala 19:72:@1052.4]
  assign _T_1001 = _T_632 ? btb_btype_45 : 2'h0; // @[Mux.scala 19:72:@1053.4]
  assign _T_1003 = _T_633 ? btb_btype_46 : 2'h0; // @[Mux.scala 19:72:@1054.4]
  assign _T_1005 = _T_634 ? btb_btype_47 : 2'h0; // @[Mux.scala 19:72:@1055.4]
  assign _T_1007 = _T_635 ? btb_btype_48 : 2'h0; // @[Mux.scala 19:72:@1056.4]
  assign _T_1009 = _T_636 ? btb_btype_49 : 2'h0; // @[Mux.scala 19:72:@1057.4]
  assign _T_1011 = _T_637 ? btb_btype_50 : 2'h0; // @[Mux.scala 19:72:@1058.4]
  assign _T_1013 = _T_638 ? btb_btype_51 : 2'h0; // @[Mux.scala 19:72:@1059.4]
  assign _T_1015 = _T_639 ? btb_btype_52 : 2'h0; // @[Mux.scala 19:72:@1060.4]
  assign _T_1017 = _T_640 ? btb_btype_53 : 2'h0; // @[Mux.scala 19:72:@1061.4]
  assign _T_1019 = _T_641 ? btb_btype_54 : 2'h0; // @[Mux.scala 19:72:@1062.4]
  assign _T_1021 = _T_642 ? btb_btype_55 : 2'h0; // @[Mux.scala 19:72:@1063.4]
  assign _T_1023 = _T_643 ? btb_btype_56 : 2'h0; // @[Mux.scala 19:72:@1064.4]
  assign _T_1025 = _T_644 ? btb_btype_57 : 2'h0; // @[Mux.scala 19:72:@1065.4]
  assign _T_1027 = _T_645 ? btb_btype_58 : 2'h0; // @[Mux.scala 19:72:@1066.4]
  assign _T_1029 = _T_646 ? btb_btype_59 : 2'h0; // @[Mux.scala 19:72:@1067.4]
  assign _T_1031 = _T_647 ? btb_btype_60 : 2'h0; // @[Mux.scala 19:72:@1068.4]
  assign _T_1033 = _T_648 ? btb_btype_61 : 2'h0; // @[Mux.scala 19:72:@1069.4]
  assign _T_1035 = _T_649 ? btb_btype_62 : 2'h0; // @[Mux.scala 19:72:@1070.4]
  assign _T_1037 = _T_650 ? btb_btype_63 : 2'h0; // @[Mux.scala 19:72:@1071.4]
  assign _T_1038 = _T_911 | _T_913; // @[Mux.scala 19:72:@1072.4]
  assign _T_1039 = _T_1038 | _T_915; // @[Mux.scala 19:72:@1073.4]
  assign _T_1040 = _T_1039 | _T_917; // @[Mux.scala 19:72:@1074.4]
  assign _T_1041 = _T_1040 | _T_919; // @[Mux.scala 19:72:@1075.4]
  assign _T_1042 = _T_1041 | _T_921; // @[Mux.scala 19:72:@1076.4]
  assign _T_1043 = _T_1042 | _T_923; // @[Mux.scala 19:72:@1077.4]
  assign _T_1044 = _T_1043 | _T_925; // @[Mux.scala 19:72:@1078.4]
  assign _T_1045 = _T_1044 | _T_927; // @[Mux.scala 19:72:@1079.4]
  assign _T_1046 = _T_1045 | _T_929; // @[Mux.scala 19:72:@1080.4]
  assign _T_1047 = _T_1046 | _T_931; // @[Mux.scala 19:72:@1081.4]
  assign _T_1048 = _T_1047 | _T_933; // @[Mux.scala 19:72:@1082.4]
  assign _T_1049 = _T_1048 | _T_935; // @[Mux.scala 19:72:@1083.4]
  assign _T_1050 = _T_1049 | _T_937; // @[Mux.scala 19:72:@1084.4]
  assign _T_1051 = _T_1050 | _T_939; // @[Mux.scala 19:72:@1085.4]
  assign _T_1052 = _T_1051 | _T_941; // @[Mux.scala 19:72:@1086.4]
  assign _T_1053 = _T_1052 | _T_943; // @[Mux.scala 19:72:@1087.4]
  assign _T_1054 = _T_1053 | _T_945; // @[Mux.scala 19:72:@1088.4]
  assign _T_1055 = _T_1054 | _T_947; // @[Mux.scala 19:72:@1089.4]
  assign _T_1056 = _T_1055 | _T_949; // @[Mux.scala 19:72:@1090.4]
  assign _T_1057 = _T_1056 | _T_951; // @[Mux.scala 19:72:@1091.4]
  assign _T_1058 = _T_1057 | _T_953; // @[Mux.scala 19:72:@1092.4]
  assign _T_1059 = _T_1058 | _T_955; // @[Mux.scala 19:72:@1093.4]
  assign _T_1060 = _T_1059 | _T_957; // @[Mux.scala 19:72:@1094.4]
  assign _T_1061 = _T_1060 | _T_959; // @[Mux.scala 19:72:@1095.4]
  assign _T_1062 = _T_1061 | _T_961; // @[Mux.scala 19:72:@1096.4]
  assign _T_1063 = _T_1062 | _T_963; // @[Mux.scala 19:72:@1097.4]
  assign _T_1064 = _T_1063 | _T_965; // @[Mux.scala 19:72:@1098.4]
  assign _T_1065 = _T_1064 | _T_967; // @[Mux.scala 19:72:@1099.4]
  assign _T_1066 = _T_1065 | _T_969; // @[Mux.scala 19:72:@1100.4]
  assign _T_1067 = _T_1066 | _T_971; // @[Mux.scala 19:72:@1101.4]
  assign _T_1068 = _T_1067 | _T_973; // @[Mux.scala 19:72:@1102.4]
  assign _T_1069 = _T_1068 | _T_975; // @[Mux.scala 19:72:@1103.4]
  assign _T_1070 = _T_1069 | _T_977; // @[Mux.scala 19:72:@1104.4]
  assign _T_1071 = _T_1070 | _T_979; // @[Mux.scala 19:72:@1105.4]
  assign _T_1072 = _T_1071 | _T_981; // @[Mux.scala 19:72:@1106.4]
  assign _T_1073 = _T_1072 | _T_983; // @[Mux.scala 19:72:@1107.4]
  assign _T_1074 = _T_1073 | _T_985; // @[Mux.scala 19:72:@1108.4]
  assign _T_1075 = _T_1074 | _T_987; // @[Mux.scala 19:72:@1109.4]
  assign _T_1076 = _T_1075 | _T_989; // @[Mux.scala 19:72:@1110.4]
  assign _T_1077 = _T_1076 | _T_991; // @[Mux.scala 19:72:@1111.4]
  assign _T_1078 = _T_1077 | _T_993; // @[Mux.scala 19:72:@1112.4]
  assign _T_1079 = _T_1078 | _T_995; // @[Mux.scala 19:72:@1113.4]
  assign _T_1080 = _T_1079 | _T_997; // @[Mux.scala 19:72:@1114.4]
  assign _T_1081 = _T_1080 | _T_999; // @[Mux.scala 19:72:@1115.4]
  assign _T_1082 = _T_1081 | _T_1001; // @[Mux.scala 19:72:@1116.4]
  assign _T_1083 = _T_1082 | _T_1003; // @[Mux.scala 19:72:@1117.4]
  assign _T_1084 = _T_1083 | _T_1005; // @[Mux.scala 19:72:@1118.4]
  assign _T_1085 = _T_1084 | _T_1007; // @[Mux.scala 19:72:@1119.4]
  assign _T_1086 = _T_1085 | _T_1009; // @[Mux.scala 19:72:@1120.4]
  assign _T_1087 = _T_1086 | _T_1011; // @[Mux.scala 19:72:@1121.4]
  assign _T_1088 = _T_1087 | _T_1013; // @[Mux.scala 19:72:@1122.4]
  assign _T_1089 = _T_1088 | _T_1015; // @[Mux.scala 19:72:@1123.4]
  assign _T_1090 = _T_1089 | _T_1017; // @[Mux.scala 19:72:@1124.4]
  assign _T_1091 = _T_1090 | _T_1019; // @[Mux.scala 19:72:@1125.4]
  assign _T_1092 = _T_1091 | _T_1021; // @[Mux.scala 19:72:@1126.4]
  assign _T_1093 = _T_1092 | _T_1023; // @[Mux.scala 19:72:@1127.4]
  assign _T_1094 = _T_1093 | _T_1025; // @[Mux.scala 19:72:@1128.4]
  assign _T_1095 = _T_1094 | _T_1027; // @[Mux.scala 19:72:@1129.4]
  assign _T_1096 = _T_1095 | _T_1029; // @[Mux.scala 19:72:@1130.4]
  assign _T_1097 = _T_1096 | _T_1031; // @[Mux.scala 19:72:@1131.4]
  assign _T_1098 = _T_1097 | _T_1033; // @[Mux.scala 19:72:@1132.4]
  assign _T_1099 = _T_1098 | _T_1035; // @[Mux.scala 19:72:@1133.4]
  assign predict_btype = _T_1099 | _T_1037; // @[Mux.scala 19:72:@1134.4]
  assign _T_1169 = _T_587 ? btb_hcount_0 : 2'h0; // @[Mux.scala 19:72:@1202.4]
  assign _T_1171 = _T_588 ? btb_hcount_1 : 2'h0; // @[Mux.scala 19:72:@1203.4]
  assign _T_1173 = _T_589 ? btb_hcount_2 : 2'h0; // @[Mux.scala 19:72:@1204.4]
  assign _T_1175 = _T_590 ? btb_hcount_3 : 2'h0; // @[Mux.scala 19:72:@1205.4]
  assign _T_1177 = _T_591 ? btb_hcount_4 : 2'h0; // @[Mux.scala 19:72:@1206.4]
  assign _T_1179 = _T_592 ? btb_hcount_5 : 2'h0; // @[Mux.scala 19:72:@1207.4]
  assign _T_1181 = _T_593 ? btb_hcount_6 : 2'h0; // @[Mux.scala 19:72:@1208.4]
  assign _T_1183 = _T_594 ? btb_hcount_7 : 2'h0; // @[Mux.scala 19:72:@1209.4]
  assign _T_1185 = _T_595 ? btb_hcount_8 : 2'h0; // @[Mux.scala 19:72:@1210.4]
  assign _T_1187 = _T_596 ? btb_hcount_9 : 2'h0; // @[Mux.scala 19:72:@1211.4]
  assign _T_1189 = _T_597 ? btb_hcount_10 : 2'h0; // @[Mux.scala 19:72:@1212.4]
  assign _T_1191 = _T_598 ? btb_hcount_11 : 2'h0; // @[Mux.scala 19:72:@1213.4]
  assign _T_1193 = _T_599 ? btb_hcount_12 : 2'h0; // @[Mux.scala 19:72:@1214.4]
  assign _T_1195 = _T_600 ? btb_hcount_13 : 2'h0; // @[Mux.scala 19:72:@1215.4]
  assign _T_1197 = _T_601 ? btb_hcount_14 : 2'h0; // @[Mux.scala 19:72:@1216.4]
  assign _T_1199 = _T_602 ? btb_hcount_15 : 2'h0; // @[Mux.scala 19:72:@1217.4]
  assign _T_1201 = _T_603 ? btb_hcount_16 : 2'h0; // @[Mux.scala 19:72:@1218.4]
  assign _T_1203 = _T_604 ? btb_hcount_17 : 2'h0; // @[Mux.scala 19:72:@1219.4]
  assign _T_1205 = _T_605 ? btb_hcount_18 : 2'h0; // @[Mux.scala 19:72:@1220.4]
  assign _T_1207 = _T_606 ? btb_hcount_19 : 2'h0; // @[Mux.scala 19:72:@1221.4]
  assign _T_1209 = _T_607 ? btb_hcount_20 : 2'h0; // @[Mux.scala 19:72:@1222.4]
  assign _T_1211 = _T_608 ? btb_hcount_21 : 2'h0; // @[Mux.scala 19:72:@1223.4]
  assign _T_1213 = _T_609 ? btb_hcount_22 : 2'h0; // @[Mux.scala 19:72:@1224.4]
  assign _T_1215 = _T_610 ? btb_hcount_23 : 2'h0; // @[Mux.scala 19:72:@1225.4]
  assign _T_1217 = _T_611 ? btb_hcount_24 : 2'h0; // @[Mux.scala 19:72:@1226.4]
  assign _T_1219 = _T_612 ? btb_hcount_25 : 2'h0; // @[Mux.scala 19:72:@1227.4]
  assign _T_1221 = _T_613 ? btb_hcount_26 : 2'h0; // @[Mux.scala 19:72:@1228.4]
  assign _T_1223 = _T_614 ? btb_hcount_27 : 2'h0; // @[Mux.scala 19:72:@1229.4]
  assign _T_1225 = _T_615 ? btb_hcount_28 : 2'h0; // @[Mux.scala 19:72:@1230.4]
  assign _T_1227 = _T_616 ? btb_hcount_29 : 2'h0; // @[Mux.scala 19:72:@1231.4]
  assign _T_1229 = _T_617 ? btb_hcount_30 : 2'h0; // @[Mux.scala 19:72:@1232.4]
  assign _T_1231 = _T_618 ? btb_hcount_31 : 2'h0; // @[Mux.scala 19:72:@1233.4]
  assign _T_1233 = _T_619 ? btb_hcount_32 : 2'h0; // @[Mux.scala 19:72:@1234.4]
  assign _T_1235 = _T_620 ? btb_hcount_33 : 2'h0; // @[Mux.scala 19:72:@1235.4]
  assign _T_1237 = _T_621 ? btb_hcount_34 : 2'h0; // @[Mux.scala 19:72:@1236.4]
  assign _T_1239 = _T_622 ? btb_hcount_35 : 2'h0; // @[Mux.scala 19:72:@1237.4]
  assign _T_1241 = _T_623 ? btb_hcount_36 : 2'h0; // @[Mux.scala 19:72:@1238.4]
  assign _T_1243 = _T_624 ? btb_hcount_37 : 2'h0; // @[Mux.scala 19:72:@1239.4]
  assign _T_1245 = _T_625 ? btb_hcount_38 : 2'h0; // @[Mux.scala 19:72:@1240.4]
  assign _T_1247 = _T_626 ? btb_hcount_39 : 2'h0; // @[Mux.scala 19:72:@1241.4]
  assign _T_1249 = _T_627 ? btb_hcount_40 : 2'h0; // @[Mux.scala 19:72:@1242.4]
  assign _T_1251 = _T_628 ? btb_hcount_41 : 2'h0; // @[Mux.scala 19:72:@1243.4]
  assign _T_1253 = _T_629 ? btb_hcount_42 : 2'h0; // @[Mux.scala 19:72:@1244.4]
  assign _T_1255 = _T_630 ? btb_hcount_43 : 2'h0; // @[Mux.scala 19:72:@1245.4]
  assign _T_1257 = _T_631 ? btb_hcount_44 : 2'h0; // @[Mux.scala 19:72:@1246.4]
  assign _T_1259 = _T_632 ? btb_hcount_45 : 2'h0; // @[Mux.scala 19:72:@1247.4]
  assign _T_1261 = _T_633 ? btb_hcount_46 : 2'h0; // @[Mux.scala 19:72:@1248.4]
  assign _T_1263 = _T_634 ? btb_hcount_47 : 2'h0; // @[Mux.scala 19:72:@1249.4]
  assign _T_1265 = _T_635 ? btb_hcount_48 : 2'h0; // @[Mux.scala 19:72:@1250.4]
  assign _T_1267 = _T_636 ? btb_hcount_49 : 2'h0; // @[Mux.scala 19:72:@1251.4]
  assign _T_1269 = _T_637 ? btb_hcount_50 : 2'h0; // @[Mux.scala 19:72:@1252.4]
  assign _T_1271 = _T_638 ? btb_hcount_51 : 2'h0; // @[Mux.scala 19:72:@1253.4]
  assign _T_1273 = _T_639 ? btb_hcount_52 : 2'h0; // @[Mux.scala 19:72:@1254.4]
  assign _T_1275 = _T_640 ? btb_hcount_53 : 2'h0; // @[Mux.scala 19:72:@1255.4]
  assign _T_1277 = _T_641 ? btb_hcount_54 : 2'h0; // @[Mux.scala 19:72:@1256.4]
  assign _T_1279 = _T_642 ? btb_hcount_55 : 2'h0; // @[Mux.scala 19:72:@1257.4]
  assign _T_1281 = _T_643 ? btb_hcount_56 : 2'h0; // @[Mux.scala 19:72:@1258.4]
  assign _T_1283 = _T_644 ? btb_hcount_57 : 2'h0; // @[Mux.scala 19:72:@1259.4]
  assign _T_1285 = _T_645 ? btb_hcount_58 : 2'h0; // @[Mux.scala 19:72:@1260.4]
  assign _T_1287 = _T_646 ? btb_hcount_59 : 2'h0; // @[Mux.scala 19:72:@1261.4]
  assign _T_1289 = _T_647 ? btb_hcount_60 : 2'h0; // @[Mux.scala 19:72:@1262.4]
  assign _T_1291 = _T_648 ? btb_hcount_61 : 2'h0; // @[Mux.scala 19:72:@1263.4]
  assign _T_1293 = _T_649 ? btb_hcount_62 : 2'h0; // @[Mux.scala 19:72:@1264.4]
  assign _T_1295 = _T_650 ? btb_hcount_63 : 2'h0; // @[Mux.scala 19:72:@1265.4]
  assign _T_1296 = _T_1169 | _T_1171; // @[Mux.scala 19:72:@1266.4]
  assign _T_1297 = _T_1296 | _T_1173; // @[Mux.scala 19:72:@1267.4]
  assign _T_1298 = _T_1297 | _T_1175; // @[Mux.scala 19:72:@1268.4]
  assign _T_1299 = _T_1298 | _T_1177; // @[Mux.scala 19:72:@1269.4]
  assign _T_1300 = _T_1299 | _T_1179; // @[Mux.scala 19:72:@1270.4]
  assign _T_1301 = _T_1300 | _T_1181; // @[Mux.scala 19:72:@1271.4]
  assign _T_1302 = _T_1301 | _T_1183; // @[Mux.scala 19:72:@1272.4]
  assign _T_1303 = _T_1302 | _T_1185; // @[Mux.scala 19:72:@1273.4]
  assign _T_1304 = _T_1303 | _T_1187; // @[Mux.scala 19:72:@1274.4]
  assign _T_1305 = _T_1304 | _T_1189; // @[Mux.scala 19:72:@1275.4]
  assign _T_1306 = _T_1305 | _T_1191; // @[Mux.scala 19:72:@1276.4]
  assign _T_1307 = _T_1306 | _T_1193; // @[Mux.scala 19:72:@1277.4]
  assign _T_1308 = _T_1307 | _T_1195; // @[Mux.scala 19:72:@1278.4]
  assign _T_1309 = _T_1308 | _T_1197; // @[Mux.scala 19:72:@1279.4]
  assign _T_1310 = _T_1309 | _T_1199; // @[Mux.scala 19:72:@1280.4]
  assign _T_1311 = _T_1310 | _T_1201; // @[Mux.scala 19:72:@1281.4]
  assign _T_1312 = _T_1311 | _T_1203; // @[Mux.scala 19:72:@1282.4]
  assign _T_1313 = _T_1312 | _T_1205; // @[Mux.scala 19:72:@1283.4]
  assign _T_1314 = _T_1313 | _T_1207; // @[Mux.scala 19:72:@1284.4]
  assign _T_1315 = _T_1314 | _T_1209; // @[Mux.scala 19:72:@1285.4]
  assign _T_1316 = _T_1315 | _T_1211; // @[Mux.scala 19:72:@1286.4]
  assign _T_1317 = _T_1316 | _T_1213; // @[Mux.scala 19:72:@1287.4]
  assign _T_1318 = _T_1317 | _T_1215; // @[Mux.scala 19:72:@1288.4]
  assign _T_1319 = _T_1318 | _T_1217; // @[Mux.scala 19:72:@1289.4]
  assign _T_1320 = _T_1319 | _T_1219; // @[Mux.scala 19:72:@1290.4]
  assign _T_1321 = _T_1320 | _T_1221; // @[Mux.scala 19:72:@1291.4]
  assign _T_1322 = _T_1321 | _T_1223; // @[Mux.scala 19:72:@1292.4]
  assign _T_1323 = _T_1322 | _T_1225; // @[Mux.scala 19:72:@1293.4]
  assign _T_1324 = _T_1323 | _T_1227; // @[Mux.scala 19:72:@1294.4]
  assign _T_1325 = _T_1324 | _T_1229; // @[Mux.scala 19:72:@1295.4]
  assign _T_1326 = _T_1325 | _T_1231; // @[Mux.scala 19:72:@1296.4]
  assign _T_1327 = _T_1326 | _T_1233; // @[Mux.scala 19:72:@1297.4]
  assign _T_1328 = _T_1327 | _T_1235; // @[Mux.scala 19:72:@1298.4]
  assign _T_1329 = _T_1328 | _T_1237; // @[Mux.scala 19:72:@1299.4]
  assign _T_1330 = _T_1329 | _T_1239; // @[Mux.scala 19:72:@1300.4]
  assign _T_1331 = _T_1330 | _T_1241; // @[Mux.scala 19:72:@1301.4]
  assign _T_1332 = _T_1331 | _T_1243; // @[Mux.scala 19:72:@1302.4]
  assign _T_1333 = _T_1332 | _T_1245; // @[Mux.scala 19:72:@1303.4]
  assign _T_1334 = _T_1333 | _T_1247; // @[Mux.scala 19:72:@1304.4]
  assign _T_1335 = _T_1334 | _T_1249; // @[Mux.scala 19:72:@1305.4]
  assign _T_1336 = _T_1335 | _T_1251; // @[Mux.scala 19:72:@1306.4]
  assign _T_1337 = _T_1336 | _T_1253; // @[Mux.scala 19:72:@1307.4]
  assign _T_1338 = _T_1337 | _T_1255; // @[Mux.scala 19:72:@1308.4]
  assign _T_1339 = _T_1338 | _T_1257; // @[Mux.scala 19:72:@1309.4]
  assign _T_1340 = _T_1339 | _T_1259; // @[Mux.scala 19:72:@1310.4]
  assign _T_1341 = _T_1340 | _T_1261; // @[Mux.scala 19:72:@1311.4]
  assign _T_1342 = _T_1341 | _T_1263; // @[Mux.scala 19:72:@1312.4]
  assign _T_1343 = _T_1342 | _T_1265; // @[Mux.scala 19:72:@1313.4]
  assign _T_1344 = _T_1343 | _T_1267; // @[Mux.scala 19:72:@1314.4]
  assign _T_1345 = _T_1344 | _T_1269; // @[Mux.scala 19:72:@1315.4]
  assign _T_1346 = _T_1345 | _T_1271; // @[Mux.scala 19:72:@1316.4]
  assign _T_1347 = _T_1346 | _T_1273; // @[Mux.scala 19:72:@1317.4]
  assign _T_1348 = _T_1347 | _T_1275; // @[Mux.scala 19:72:@1318.4]
  assign _T_1349 = _T_1348 | _T_1277; // @[Mux.scala 19:72:@1319.4]
  assign _T_1350 = _T_1349 | _T_1279; // @[Mux.scala 19:72:@1320.4]
  assign _T_1351 = _T_1350 | _T_1281; // @[Mux.scala 19:72:@1321.4]
  assign _T_1352 = _T_1351 | _T_1283; // @[Mux.scala 19:72:@1322.4]
  assign _T_1353 = _T_1352 | _T_1285; // @[Mux.scala 19:72:@1323.4]
  assign _T_1354 = _T_1353 | _T_1287; // @[Mux.scala 19:72:@1324.4]
  assign _T_1355 = _T_1354 | _T_1289; // @[Mux.scala 19:72:@1325.4]
  assign _T_1356 = _T_1355 | _T_1291; // @[Mux.scala 19:72:@1326.4]
  assign _T_1357 = _T_1356 | _T_1293; // @[Mux.scala 19:72:@1327.4]
  assign predict_hcount = _T_1357 | _T_1295; // @[Mux.scala 19:72:@1328.4]
  assign _T_1362 = predict_btype == 2'h1; // @[BTB.scala 76:35:@1332.4]
  assign _T_1364 = predict_btype == 2'h2; // @[BTB.scala 67:36:@1333.4]
  assign _T_1365 = predict_hcount[1]; // @[BTB.scala 67:67:@1334.4]
  assign _T_1367 = _T_1365 == 1'h0; // @[BTB.scala 67:60:@1335.4]
  assign _T_1368 = _T_1364 & _T_1367; // @[BTB.scala 67:57:@1336.4]
  assign _T_1370 = _T_1368 == 1'h0; // @[BTB.scala 67:28:@1337.4]
  assign _T_1372 = predict_lookup != 64'h0; // @[BTB.scala 67:82:@1338.4]
  assign _T_1373 = _T_1370 & _T_1372; // @[BTB.scala 67:72:@1339.4]
  assign _T_1374 = _T_1373 ? predict_jump_tgt : predict_cont_tgt; // @[BTB.scala 67:27:@1340.4]
  assign _T_1382 = fb_reg_lfsr[0]; // @[BTB.scala 90:36:@1356.4]
  assign _T_1383 = fb_reg_lfsr[1]; // @[BTB.scala 90:46:@1357.4]
  assign _T_1384 = _T_1382 ^ _T_1383; // @[BTB.scala 90:40:@1358.4]
  assign _T_1385 = fb_reg_lfsr[5:1]; // @[BTB.scala 90:55:@1359.4]
  assign _T_1386 = {_T_1384,_T_1385}; // @[Cat.scala 30:58:@1360.4]
  assign _T_1388 = btb_pc_0 == fb_reg_pc; // @[BTB.scala 114:42:@1363.4]
  assign _T_1389 = btb_pc_1 == fb_reg_pc; // @[BTB.scala 114:42:@1364.4]
  assign _T_1390 = btb_pc_2 == fb_reg_pc; // @[BTB.scala 114:42:@1365.4]
  assign _T_1391 = btb_pc_3 == fb_reg_pc; // @[BTB.scala 114:42:@1366.4]
  assign _T_1392 = btb_pc_4 == fb_reg_pc; // @[BTB.scala 114:42:@1367.4]
  assign _T_1393 = btb_pc_5 == fb_reg_pc; // @[BTB.scala 114:42:@1368.4]
  assign _T_1394 = btb_pc_6 == fb_reg_pc; // @[BTB.scala 114:42:@1369.4]
  assign _T_1395 = btb_pc_7 == fb_reg_pc; // @[BTB.scala 114:42:@1370.4]
  assign _T_1396 = btb_pc_8 == fb_reg_pc; // @[BTB.scala 114:42:@1371.4]
  assign _T_1397 = btb_pc_9 == fb_reg_pc; // @[BTB.scala 114:42:@1372.4]
  assign _T_1398 = btb_pc_10 == fb_reg_pc; // @[BTB.scala 114:42:@1373.4]
  assign _T_1399 = btb_pc_11 == fb_reg_pc; // @[BTB.scala 114:42:@1374.4]
  assign _T_1400 = btb_pc_12 == fb_reg_pc; // @[BTB.scala 114:42:@1375.4]
  assign _T_1401 = btb_pc_13 == fb_reg_pc; // @[BTB.scala 114:42:@1376.4]
  assign _T_1402 = btb_pc_14 == fb_reg_pc; // @[BTB.scala 114:42:@1377.4]
  assign _T_1403 = btb_pc_15 == fb_reg_pc; // @[BTB.scala 114:42:@1378.4]
  assign _T_1404 = btb_pc_16 == fb_reg_pc; // @[BTB.scala 114:42:@1379.4]
  assign _T_1405 = btb_pc_17 == fb_reg_pc; // @[BTB.scala 114:42:@1380.4]
  assign _T_1406 = btb_pc_18 == fb_reg_pc; // @[BTB.scala 114:42:@1381.4]
  assign _T_1407 = btb_pc_19 == fb_reg_pc; // @[BTB.scala 114:42:@1382.4]
  assign _T_1408 = btb_pc_20 == fb_reg_pc; // @[BTB.scala 114:42:@1383.4]
  assign _T_1409 = btb_pc_21 == fb_reg_pc; // @[BTB.scala 114:42:@1384.4]
  assign _T_1410 = btb_pc_22 == fb_reg_pc; // @[BTB.scala 114:42:@1385.4]
  assign _T_1411 = btb_pc_23 == fb_reg_pc; // @[BTB.scala 114:42:@1386.4]
  assign _T_1412 = btb_pc_24 == fb_reg_pc; // @[BTB.scala 114:42:@1387.4]
  assign _T_1413 = btb_pc_25 == fb_reg_pc; // @[BTB.scala 114:42:@1388.4]
  assign _T_1414 = btb_pc_26 == fb_reg_pc; // @[BTB.scala 114:42:@1389.4]
  assign _T_1415 = btb_pc_27 == fb_reg_pc; // @[BTB.scala 114:42:@1390.4]
  assign _T_1416 = btb_pc_28 == fb_reg_pc; // @[BTB.scala 114:42:@1391.4]
  assign _T_1417 = btb_pc_29 == fb_reg_pc; // @[BTB.scala 114:42:@1392.4]
  assign _T_1418 = btb_pc_30 == fb_reg_pc; // @[BTB.scala 114:42:@1393.4]
  assign _T_1419 = btb_pc_31 == fb_reg_pc; // @[BTB.scala 114:42:@1394.4]
  assign _T_1420 = btb_pc_32 == fb_reg_pc; // @[BTB.scala 114:42:@1395.4]
  assign _T_1421 = btb_pc_33 == fb_reg_pc; // @[BTB.scala 114:42:@1396.4]
  assign _T_1422 = btb_pc_34 == fb_reg_pc; // @[BTB.scala 114:42:@1397.4]
  assign _T_1423 = btb_pc_35 == fb_reg_pc; // @[BTB.scala 114:42:@1398.4]
  assign _T_1424 = btb_pc_36 == fb_reg_pc; // @[BTB.scala 114:42:@1399.4]
  assign _T_1425 = btb_pc_37 == fb_reg_pc; // @[BTB.scala 114:42:@1400.4]
  assign _T_1426 = btb_pc_38 == fb_reg_pc; // @[BTB.scala 114:42:@1401.4]
  assign _T_1427 = btb_pc_39 == fb_reg_pc; // @[BTB.scala 114:42:@1402.4]
  assign _T_1428 = btb_pc_40 == fb_reg_pc; // @[BTB.scala 114:42:@1403.4]
  assign _T_1429 = btb_pc_41 == fb_reg_pc; // @[BTB.scala 114:42:@1404.4]
  assign _T_1430 = btb_pc_42 == fb_reg_pc; // @[BTB.scala 114:42:@1405.4]
  assign _T_1431 = btb_pc_43 == fb_reg_pc; // @[BTB.scala 114:42:@1406.4]
  assign _T_1432 = btb_pc_44 == fb_reg_pc; // @[BTB.scala 114:42:@1407.4]
  assign _T_1433 = btb_pc_45 == fb_reg_pc; // @[BTB.scala 114:42:@1408.4]
  assign _T_1434 = btb_pc_46 == fb_reg_pc; // @[BTB.scala 114:42:@1409.4]
  assign _T_1435 = btb_pc_47 == fb_reg_pc; // @[BTB.scala 114:42:@1410.4]
  assign _T_1436 = btb_pc_48 == fb_reg_pc; // @[BTB.scala 114:42:@1411.4]
  assign _T_1437 = btb_pc_49 == fb_reg_pc; // @[BTB.scala 114:42:@1412.4]
  assign _T_1438 = btb_pc_50 == fb_reg_pc; // @[BTB.scala 114:42:@1413.4]
  assign _T_1439 = btb_pc_51 == fb_reg_pc; // @[BTB.scala 114:42:@1414.4]
  assign _T_1440 = btb_pc_52 == fb_reg_pc; // @[BTB.scala 114:42:@1415.4]
  assign _T_1441 = btb_pc_53 == fb_reg_pc; // @[BTB.scala 114:42:@1416.4]
  assign _T_1442 = btb_pc_54 == fb_reg_pc; // @[BTB.scala 114:42:@1417.4]
  assign _T_1443 = btb_pc_55 == fb_reg_pc; // @[BTB.scala 114:42:@1418.4]
  assign _T_1444 = btb_pc_56 == fb_reg_pc; // @[BTB.scala 114:42:@1419.4]
  assign _T_1445 = btb_pc_57 == fb_reg_pc; // @[BTB.scala 114:42:@1420.4]
  assign _T_1446 = btb_pc_58 == fb_reg_pc; // @[BTB.scala 114:42:@1421.4]
  assign _T_1447 = btb_pc_59 == fb_reg_pc; // @[BTB.scala 114:42:@1422.4]
  assign _T_1448 = btb_pc_60 == fb_reg_pc; // @[BTB.scala 114:42:@1423.4]
  assign _T_1449 = btb_pc_61 == fb_reg_pc; // @[BTB.scala 114:42:@1424.4]
  assign _T_1450 = btb_pc_62 == fb_reg_pc; // @[BTB.scala 114:42:@1425.4]
  assign _T_1451 = btb_pc_63 == fb_reg_pc; // @[BTB.scala 114:42:@1426.4]
  assign _T_1528 = {_T_1395,_T_1394,_T_1393,_T_1392,_T_1391,_T_1390,_T_1389,_T_1388}; // @[BTB.scala 114:58:@1498.4]
  assign _T_1536 = {_T_1403,_T_1402,_T_1401,_T_1400,_T_1399,_T_1398,_T_1397,_T_1396,_T_1528}; // @[BTB.scala 114:58:@1506.4]
  assign _T_1543 = {_T_1411,_T_1410,_T_1409,_T_1408,_T_1407,_T_1406,_T_1405,_T_1404}; // @[BTB.scala 114:58:@1513.4]
  assign _T_1552 = {_T_1419,_T_1418,_T_1417,_T_1416,_T_1415,_T_1414,_T_1413,_T_1412,_T_1543,_T_1536}; // @[BTB.scala 114:58:@1522.4]
  assign _T_1559 = {_T_1427,_T_1426,_T_1425,_T_1424,_T_1423,_T_1422,_T_1421,_T_1420}; // @[BTB.scala 114:58:@1529.4]
  assign _T_1567 = {_T_1435,_T_1434,_T_1433,_T_1432,_T_1431,_T_1430,_T_1429,_T_1428,_T_1559}; // @[BTB.scala 114:58:@1537.4]
  assign _T_1574 = {_T_1443,_T_1442,_T_1441,_T_1440,_T_1439,_T_1438,_T_1437,_T_1436}; // @[BTB.scala 114:58:@1544.4]
  assign _T_1583 = {_T_1451,_T_1450,_T_1449,_T_1448,_T_1447,_T_1446,_T_1445,_T_1444,_T_1574,_T_1567}; // @[BTB.scala 114:58:@1553.4]
  assign _T_1584 = {_T_1583,_T_1552}; // @[BTB.scala 114:58:@1554.4]
  assign fb_wire_lookup = _T_1584 & _T_582; // @[BTB.scala 114:65:@1747.4]
  assign _T_1847 = fb_wire_lookup[0]; // @[Mux.scala 21:36:@1749.4]
  assign _T_1848 = fb_wire_lookup[1]; // @[Mux.scala 21:36:@1750.4]
  assign _T_1849 = fb_wire_lookup[2]; // @[Mux.scala 21:36:@1751.4]
  assign _T_1850 = fb_wire_lookup[3]; // @[Mux.scala 21:36:@1752.4]
  assign _T_1851 = fb_wire_lookup[4]; // @[Mux.scala 21:36:@1753.4]
  assign _T_1852 = fb_wire_lookup[5]; // @[Mux.scala 21:36:@1754.4]
  assign _T_1853 = fb_wire_lookup[6]; // @[Mux.scala 21:36:@1755.4]
  assign _T_1854 = fb_wire_lookup[7]; // @[Mux.scala 21:36:@1756.4]
  assign _T_1855 = fb_wire_lookup[8]; // @[Mux.scala 21:36:@1757.4]
  assign _T_1856 = fb_wire_lookup[9]; // @[Mux.scala 21:36:@1758.4]
  assign _T_1857 = fb_wire_lookup[10]; // @[Mux.scala 21:36:@1759.4]
  assign _T_1858 = fb_wire_lookup[11]; // @[Mux.scala 21:36:@1760.4]
  assign _T_1859 = fb_wire_lookup[12]; // @[Mux.scala 21:36:@1761.4]
  assign _T_1860 = fb_wire_lookup[13]; // @[Mux.scala 21:36:@1762.4]
  assign _T_1861 = fb_wire_lookup[14]; // @[Mux.scala 21:36:@1763.4]
  assign _T_1862 = fb_wire_lookup[15]; // @[Mux.scala 21:36:@1764.4]
  assign _T_1863 = fb_wire_lookup[16]; // @[Mux.scala 21:36:@1765.4]
  assign _T_1864 = fb_wire_lookup[17]; // @[Mux.scala 21:36:@1766.4]
  assign _T_1865 = fb_wire_lookup[18]; // @[Mux.scala 21:36:@1767.4]
  assign _T_1866 = fb_wire_lookup[19]; // @[Mux.scala 21:36:@1768.4]
  assign _T_1867 = fb_wire_lookup[20]; // @[Mux.scala 21:36:@1769.4]
  assign _T_1868 = fb_wire_lookup[21]; // @[Mux.scala 21:36:@1770.4]
  assign _T_1869 = fb_wire_lookup[22]; // @[Mux.scala 21:36:@1771.4]
  assign _T_1870 = fb_wire_lookup[23]; // @[Mux.scala 21:36:@1772.4]
  assign _T_1871 = fb_wire_lookup[24]; // @[Mux.scala 21:36:@1773.4]
  assign _T_1872 = fb_wire_lookup[25]; // @[Mux.scala 21:36:@1774.4]
  assign _T_1873 = fb_wire_lookup[26]; // @[Mux.scala 21:36:@1775.4]
  assign _T_1874 = fb_wire_lookup[27]; // @[Mux.scala 21:36:@1776.4]
  assign _T_1875 = fb_wire_lookup[28]; // @[Mux.scala 21:36:@1777.4]
  assign _T_1876 = fb_wire_lookup[29]; // @[Mux.scala 21:36:@1778.4]
  assign _T_1877 = fb_wire_lookup[30]; // @[Mux.scala 21:36:@1779.4]
  assign _T_1878 = fb_wire_lookup[31]; // @[Mux.scala 21:36:@1780.4]
  assign _T_1879 = fb_wire_lookup[32]; // @[Mux.scala 21:36:@1781.4]
  assign _T_1880 = fb_wire_lookup[33]; // @[Mux.scala 21:36:@1782.4]
  assign _T_1881 = fb_wire_lookup[34]; // @[Mux.scala 21:36:@1783.4]
  assign _T_1882 = fb_wire_lookup[35]; // @[Mux.scala 21:36:@1784.4]
  assign _T_1883 = fb_wire_lookup[36]; // @[Mux.scala 21:36:@1785.4]
  assign _T_1884 = fb_wire_lookup[37]; // @[Mux.scala 21:36:@1786.4]
  assign _T_1885 = fb_wire_lookup[38]; // @[Mux.scala 21:36:@1787.4]
  assign _T_1886 = fb_wire_lookup[39]; // @[Mux.scala 21:36:@1788.4]
  assign _T_1887 = fb_wire_lookup[40]; // @[Mux.scala 21:36:@1789.4]
  assign _T_1888 = fb_wire_lookup[41]; // @[Mux.scala 21:36:@1790.4]
  assign _T_1889 = fb_wire_lookup[42]; // @[Mux.scala 21:36:@1791.4]
  assign _T_1890 = fb_wire_lookup[43]; // @[Mux.scala 21:36:@1792.4]
  assign _T_1891 = fb_wire_lookup[44]; // @[Mux.scala 21:36:@1793.4]
  assign _T_1892 = fb_wire_lookup[45]; // @[Mux.scala 21:36:@1794.4]
  assign _T_1893 = fb_wire_lookup[46]; // @[Mux.scala 21:36:@1795.4]
  assign _T_1894 = fb_wire_lookup[47]; // @[Mux.scala 21:36:@1796.4]
  assign _T_1895 = fb_wire_lookup[48]; // @[Mux.scala 21:36:@1797.4]
  assign _T_1896 = fb_wire_lookup[49]; // @[Mux.scala 21:36:@1798.4]
  assign _T_1897 = fb_wire_lookup[50]; // @[Mux.scala 21:36:@1799.4]
  assign _T_1898 = fb_wire_lookup[51]; // @[Mux.scala 21:36:@1800.4]
  assign _T_1899 = fb_wire_lookup[52]; // @[Mux.scala 21:36:@1801.4]
  assign _T_1900 = fb_wire_lookup[53]; // @[Mux.scala 21:36:@1802.4]
  assign _T_1901 = fb_wire_lookup[54]; // @[Mux.scala 21:36:@1803.4]
  assign _T_1902 = fb_wire_lookup[55]; // @[Mux.scala 21:36:@1804.4]
  assign _T_1903 = fb_wire_lookup[56]; // @[Mux.scala 21:36:@1805.4]
  assign _T_1904 = fb_wire_lookup[57]; // @[Mux.scala 21:36:@1806.4]
  assign _T_1905 = fb_wire_lookup[58]; // @[Mux.scala 21:36:@1807.4]
  assign _T_1906 = fb_wire_lookup[59]; // @[Mux.scala 21:36:@1808.4]
  assign _T_1907 = fb_wire_lookup[60]; // @[Mux.scala 21:36:@1809.4]
  assign _T_1908 = fb_wire_lookup[61]; // @[Mux.scala 21:36:@1810.4]
  assign _T_1909 = fb_wire_lookup[62]; // @[Mux.scala 21:36:@1811.4]
  assign _T_1910 = fb_wire_lookup[63]; // @[Mux.scala 21:36:@1812.4]
  assign _T_1913 = _T_1847 ? btb_hcount_0 : 2'h0; // @[Mux.scala 19:72:@1813.4]
  assign _T_1915 = _T_1848 ? btb_hcount_1 : 2'h0; // @[Mux.scala 19:72:@1814.4]
  assign _T_1917 = _T_1849 ? btb_hcount_2 : 2'h0; // @[Mux.scala 19:72:@1815.4]
  assign _T_1919 = _T_1850 ? btb_hcount_3 : 2'h0; // @[Mux.scala 19:72:@1816.4]
  assign _T_1921 = _T_1851 ? btb_hcount_4 : 2'h0; // @[Mux.scala 19:72:@1817.4]
  assign _T_1923 = _T_1852 ? btb_hcount_5 : 2'h0; // @[Mux.scala 19:72:@1818.4]
  assign _T_1925 = _T_1853 ? btb_hcount_6 : 2'h0; // @[Mux.scala 19:72:@1819.4]
  assign _T_1927 = _T_1854 ? btb_hcount_7 : 2'h0; // @[Mux.scala 19:72:@1820.4]
  assign _T_1929 = _T_1855 ? btb_hcount_8 : 2'h0; // @[Mux.scala 19:72:@1821.4]
  assign _T_1931 = _T_1856 ? btb_hcount_9 : 2'h0; // @[Mux.scala 19:72:@1822.4]
  assign _T_1933 = _T_1857 ? btb_hcount_10 : 2'h0; // @[Mux.scala 19:72:@1823.4]
  assign _T_1935 = _T_1858 ? btb_hcount_11 : 2'h0; // @[Mux.scala 19:72:@1824.4]
  assign _T_1937 = _T_1859 ? btb_hcount_12 : 2'h0; // @[Mux.scala 19:72:@1825.4]
  assign _T_1939 = _T_1860 ? btb_hcount_13 : 2'h0; // @[Mux.scala 19:72:@1826.4]
  assign _T_1941 = _T_1861 ? btb_hcount_14 : 2'h0; // @[Mux.scala 19:72:@1827.4]
  assign _T_1943 = _T_1862 ? btb_hcount_15 : 2'h0; // @[Mux.scala 19:72:@1828.4]
  assign _T_1945 = _T_1863 ? btb_hcount_16 : 2'h0; // @[Mux.scala 19:72:@1829.4]
  assign _T_1947 = _T_1864 ? btb_hcount_17 : 2'h0; // @[Mux.scala 19:72:@1830.4]
  assign _T_1949 = _T_1865 ? btb_hcount_18 : 2'h0; // @[Mux.scala 19:72:@1831.4]
  assign _T_1951 = _T_1866 ? btb_hcount_19 : 2'h0; // @[Mux.scala 19:72:@1832.4]
  assign _T_1953 = _T_1867 ? btb_hcount_20 : 2'h0; // @[Mux.scala 19:72:@1833.4]
  assign _T_1955 = _T_1868 ? btb_hcount_21 : 2'h0; // @[Mux.scala 19:72:@1834.4]
  assign _T_1957 = _T_1869 ? btb_hcount_22 : 2'h0; // @[Mux.scala 19:72:@1835.4]
  assign _T_1959 = _T_1870 ? btb_hcount_23 : 2'h0; // @[Mux.scala 19:72:@1836.4]
  assign _T_1961 = _T_1871 ? btb_hcount_24 : 2'h0; // @[Mux.scala 19:72:@1837.4]
  assign _T_1963 = _T_1872 ? btb_hcount_25 : 2'h0; // @[Mux.scala 19:72:@1838.4]
  assign _T_1965 = _T_1873 ? btb_hcount_26 : 2'h0; // @[Mux.scala 19:72:@1839.4]
  assign _T_1967 = _T_1874 ? btb_hcount_27 : 2'h0; // @[Mux.scala 19:72:@1840.4]
  assign _T_1969 = _T_1875 ? btb_hcount_28 : 2'h0; // @[Mux.scala 19:72:@1841.4]
  assign _T_1971 = _T_1876 ? btb_hcount_29 : 2'h0; // @[Mux.scala 19:72:@1842.4]
  assign _T_1973 = _T_1877 ? btb_hcount_30 : 2'h0; // @[Mux.scala 19:72:@1843.4]
  assign _T_1975 = _T_1878 ? btb_hcount_31 : 2'h0; // @[Mux.scala 19:72:@1844.4]
  assign _T_1977 = _T_1879 ? btb_hcount_32 : 2'h0; // @[Mux.scala 19:72:@1845.4]
  assign _T_1979 = _T_1880 ? btb_hcount_33 : 2'h0; // @[Mux.scala 19:72:@1846.4]
  assign _T_1981 = _T_1881 ? btb_hcount_34 : 2'h0; // @[Mux.scala 19:72:@1847.4]
  assign _T_1983 = _T_1882 ? btb_hcount_35 : 2'h0; // @[Mux.scala 19:72:@1848.4]
  assign _T_1985 = _T_1883 ? btb_hcount_36 : 2'h0; // @[Mux.scala 19:72:@1849.4]
  assign _T_1987 = _T_1884 ? btb_hcount_37 : 2'h0; // @[Mux.scala 19:72:@1850.4]
  assign _T_1989 = _T_1885 ? btb_hcount_38 : 2'h0; // @[Mux.scala 19:72:@1851.4]
  assign _T_1991 = _T_1886 ? btb_hcount_39 : 2'h0; // @[Mux.scala 19:72:@1852.4]
  assign _T_1993 = _T_1887 ? btb_hcount_40 : 2'h0; // @[Mux.scala 19:72:@1853.4]
  assign _T_1995 = _T_1888 ? btb_hcount_41 : 2'h0; // @[Mux.scala 19:72:@1854.4]
  assign _T_1997 = _T_1889 ? btb_hcount_42 : 2'h0; // @[Mux.scala 19:72:@1855.4]
  assign _T_1999 = _T_1890 ? btb_hcount_43 : 2'h0; // @[Mux.scala 19:72:@1856.4]
  assign _T_2001 = _T_1891 ? btb_hcount_44 : 2'h0; // @[Mux.scala 19:72:@1857.4]
  assign _T_2003 = _T_1892 ? btb_hcount_45 : 2'h0; // @[Mux.scala 19:72:@1858.4]
  assign _T_2005 = _T_1893 ? btb_hcount_46 : 2'h0; // @[Mux.scala 19:72:@1859.4]
  assign _T_2007 = _T_1894 ? btb_hcount_47 : 2'h0; // @[Mux.scala 19:72:@1860.4]
  assign _T_2009 = _T_1895 ? btb_hcount_48 : 2'h0; // @[Mux.scala 19:72:@1861.4]
  assign _T_2011 = _T_1896 ? btb_hcount_49 : 2'h0; // @[Mux.scala 19:72:@1862.4]
  assign _T_2013 = _T_1897 ? btb_hcount_50 : 2'h0; // @[Mux.scala 19:72:@1863.4]
  assign _T_2015 = _T_1898 ? btb_hcount_51 : 2'h0; // @[Mux.scala 19:72:@1864.4]
  assign _T_2017 = _T_1899 ? btb_hcount_52 : 2'h0; // @[Mux.scala 19:72:@1865.4]
  assign _T_2019 = _T_1900 ? btb_hcount_53 : 2'h0; // @[Mux.scala 19:72:@1866.4]
  assign _T_2021 = _T_1901 ? btb_hcount_54 : 2'h0; // @[Mux.scala 19:72:@1867.4]
  assign _T_2023 = _T_1902 ? btb_hcount_55 : 2'h0; // @[Mux.scala 19:72:@1868.4]
  assign _T_2025 = _T_1903 ? btb_hcount_56 : 2'h0; // @[Mux.scala 19:72:@1869.4]
  assign _T_2027 = _T_1904 ? btb_hcount_57 : 2'h0; // @[Mux.scala 19:72:@1870.4]
  assign _T_2029 = _T_1905 ? btb_hcount_58 : 2'h0; // @[Mux.scala 19:72:@1871.4]
  assign _T_2031 = _T_1906 ? btb_hcount_59 : 2'h0; // @[Mux.scala 19:72:@1872.4]
  assign _T_2033 = _T_1907 ? btb_hcount_60 : 2'h0; // @[Mux.scala 19:72:@1873.4]
  assign _T_2035 = _T_1908 ? btb_hcount_61 : 2'h0; // @[Mux.scala 19:72:@1874.4]
  assign _T_2037 = _T_1909 ? btb_hcount_62 : 2'h0; // @[Mux.scala 19:72:@1875.4]
  assign _T_2039 = _T_1910 ? btb_hcount_63 : 2'h0; // @[Mux.scala 19:72:@1876.4]
  assign _T_2040 = _T_1913 | _T_1915; // @[Mux.scala 19:72:@1877.4]
  assign _T_2041 = _T_2040 | _T_1917; // @[Mux.scala 19:72:@1878.4]
  assign _T_2042 = _T_2041 | _T_1919; // @[Mux.scala 19:72:@1879.4]
  assign _T_2043 = _T_2042 | _T_1921; // @[Mux.scala 19:72:@1880.4]
  assign _T_2044 = _T_2043 | _T_1923; // @[Mux.scala 19:72:@1881.4]
  assign _T_2045 = _T_2044 | _T_1925; // @[Mux.scala 19:72:@1882.4]
  assign _T_2046 = _T_2045 | _T_1927; // @[Mux.scala 19:72:@1883.4]
  assign _T_2047 = _T_2046 | _T_1929; // @[Mux.scala 19:72:@1884.4]
  assign _T_2048 = _T_2047 | _T_1931; // @[Mux.scala 19:72:@1885.4]
  assign _T_2049 = _T_2048 | _T_1933; // @[Mux.scala 19:72:@1886.4]
  assign _T_2050 = _T_2049 | _T_1935; // @[Mux.scala 19:72:@1887.4]
  assign _T_2051 = _T_2050 | _T_1937; // @[Mux.scala 19:72:@1888.4]
  assign _T_2052 = _T_2051 | _T_1939; // @[Mux.scala 19:72:@1889.4]
  assign _T_2053 = _T_2052 | _T_1941; // @[Mux.scala 19:72:@1890.4]
  assign _T_2054 = _T_2053 | _T_1943; // @[Mux.scala 19:72:@1891.4]
  assign _T_2055 = _T_2054 | _T_1945; // @[Mux.scala 19:72:@1892.4]
  assign _T_2056 = _T_2055 | _T_1947; // @[Mux.scala 19:72:@1893.4]
  assign _T_2057 = _T_2056 | _T_1949; // @[Mux.scala 19:72:@1894.4]
  assign _T_2058 = _T_2057 | _T_1951; // @[Mux.scala 19:72:@1895.4]
  assign _T_2059 = _T_2058 | _T_1953; // @[Mux.scala 19:72:@1896.4]
  assign _T_2060 = _T_2059 | _T_1955; // @[Mux.scala 19:72:@1897.4]
  assign _T_2061 = _T_2060 | _T_1957; // @[Mux.scala 19:72:@1898.4]
  assign _T_2062 = _T_2061 | _T_1959; // @[Mux.scala 19:72:@1899.4]
  assign _T_2063 = _T_2062 | _T_1961; // @[Mux.scala 19:72:@1900.4]
  assign _T_2064 = _T_2063 | _T_1963; // @[Mux.scala 19:72:@1901.4]
  assign _T_2065 = _T_2064 | _T_1965; // @[Mux.scala 19:72:@1902.4]
  assign _T_2066 = _T_2065 | _T_1967; // @[Mux.scala 19:72:@1903.4]
  assign _T_2067 = _T_2066 | _T_1969; // @[Mux.scala 19:72:@1904.4]
  assign _T_2068 = _T_2067 | _T_1971; // @[Mux.scala 19:72:@1905.4]
  assign _T_2069 = _T_2068 | _T_1973; // @[Mux.scala 19:72:@1906.4]
  assign _T_2070 = _T_2069 | _T_1975; // @[Mux.scala 19:72:@1907.4]
  assign _T_2071 = _T_2070 | _T_1977; // @[Mux.scala 19:72:@1908.4]
  assign _T_2072 = _T_2071 | _T_1979; // @[Mux.scala 19:72:@1909.4]
  assign _T_2073 = _T_2072 | _T_1981; // @[Mux.scala 19:72:@1910.4]
  assign _T_2074 = _T_2073 | _T_1983; // @[Mux.scala 19:72:@1911.4]
  assign _T_2075 = _T_2074 | _T_1985; // @[Mux.scala 19:72:@1912.4]
  assign _T_2076 = _T_2075 | _T_1987; // @[Mux.scala 19:72:@1913.4]
  assign _T_2077 = _T_2076 | _T_1989; // @[Mux.scala 19:72:@1914.4]
  assign _T_2078 = _T_2077 | _T_1991; // @[Mux.scala 19:72:@1915.4]
  assign _T_2079 = _T_2078 | _T_1993; // @[Mux.scala 19:72:@1916.4]
  assign _T_2080 = _T_2079 | _T_1995; // @[Mux.scala 19:72:@1917.4]
  assign _T_2081 = _T_2080 | _T_1997; // @[Mux.scala 19:72:@1918.4]
  assign _T_2082 = _T_2081 | _T_1999; // @[Mux.scala 19:72:@1919.4]
  assign _T_2083 = _T_2082 | _T_2001; // @[Mux.scala 19:72:@1920.4]
  assign _T_2084 = _T_2083 | _T_2003; // @[Mux.scala 19:72:@1921.4]
  assign _T_2085 = _T_2084 | _T_2005; // @[Mux.scala 19:72:@1922.4]
  assign _T_2086 = _T_2085 | _T_2007; // @[Mux.scala 19:72:@1923.4]
  assign _T_2087 = _T_2086 | _T_2009; // @[Mux.scala 19:72:@1924.4]
  assign _T_2088 = _T_2087 | _T_2011; // @[Mux.scala 19:72:@1925.4]
  assign _T_2089 = _T_2088 | _T_2013; // @[Mux.scala 19:72:@1926.4]
  assign _T_2090 = _T_2089 | _T_2015; // @[Mux.scala 19:72:@1927.4]
  assign _T_2091 = _T_2090 | _T_2017; // @[Mux.scala 19:72:@1928.4]
  assign _T_2092 = _T_2091 | _T_2019; // @[Mux.scala 19:72:@1929.4]
  assign _T_2093 = _T_2092 | _T_2021; // @[Mux.scala 19:72:@1930.4]
  assign _T_2094 = _T_2093 | _T_2023; // @[Mux.scala 19:72:@1931.4]
  assign _T_2095 = _T_2094 | _T_2025; // @[Mux.scala 19:72:@1932.4]
  assign _T_2096 = _T_2095 | _T_2027; // @[Mux.scala 19:72:@1933.4]
  assign _T_2097 = _T_2096 | _T_2029; // @[Mux.scala 19:72:@1934.4]
  assign _T_2098 = _T_2097 | _T_2031; // @[Mux.scala 19:72:@1935.4]
  assign _T_2099 = _T_2098 | _T_2033; // @[Mux.scala 19:72:@1936.4]
  assign _T_2100 = _T_2099 | _T_2035; // @[Mux.scala 19:72:@1937.4]
  assign _T_2101 = _T_2100 | _T_2037; // @[Mux.scala 19:72:@1938.4]
  assign fb_wire_hcount = _T_2101 | _T_2039; // @[Mux.scala 19:72:@1939.4]
  assign _T_2106 = fb_wire_lookup != 64'h0; // @[BTB.scala 112:30:@1943.4]
  assign _T_2107 = fb_wire_lookup[63:32]; // @[OneHot.scala 26:18:@1944.4]
  assign _T_2108 = fb_wire_lookup[31:0]; // @[OneHot.scala 27:18:@1945.4]
  assign _T_2110 = _T_2107 != 32'h0; // @[OneHot.scala 28:14:@1946.4]
  assign _T_2111 = _T_2107 | _T_2108; // @[OneHot.scala 28:28:@1947.4]
  assign _T_2112 = _T_2111[31:16]; // @[OneHot.scala 26:18:@1948.4]
  assign _T_2113 = _T_2111[15:0]; // @[OneHot.scala 27:18:@1949.4]
  assign _T_2115 = _T_2112 != 16'h0; // @[OneHot.scala 28:14:@1950.4]
  assign _T_2116 = _T_2112 | _T_2113; // @[OneHot.scala 28:28:@1951.4]
  assign _T_2117 = _T_2116[15:8]; // @[OneHot.scala 26:18:@1952.4]
  assign _T_2118 = _T_2116[7:0]; // @[OneHot.scala 27:18:@1953.4]
  assign _T_2120 = _T_2117 != 8'h0; // @[OneHot.scala 28:14:@1954.4]
  assign _T_2121 = _T_2117 | _T_2118; // @[OneHot.scala 28:28:@1955.4]
  assign _T_2122 = _T_2121[7:4]; // @[OneHot.scala 26:18:@1956.4]
  assign _T_2123 = _T_2121[3:0]; // @[OneHot.scala 27:18:@1957.4]
  assign _T_2125 = _T_2122 != 4'h0; // @[OneHot.scala 28:14:@1958.4]
  assign _T_2126 = _T_2122 | _T_2123; // @[OneHot.scala 28:28:@1959.4]
  assign _T_2127 = _T_2126[3:2]; // @[OneHot.scala 26:18:@1960.4]
  assign _T_2128 = _T_2126[1:0]; // @[OneHot.scala 27:18:@1961.4]
  assign _T_2130 = _T_2127 != 2'h0; // @[OneHot.scala 28:14:@1962.4]
  assign _T_2131 = _T_2127 | _T_2128; // @[OneHot.scala 28:28:@1963.4]
  assign _T_2132 = _T_2131[1]; // @[CircuitMath.scala 30:8:@1964.4]
  assign _T_2137 = {_T_2110,_T_2115,_T_2120,_T_2125,_T_2130,_T_2132}; // @[Cat.scala 30:58:@1969.4]
  assign _T_2399 = ~ _T_582; // @[BTB.scala 118:19:@2162.4]
  assign _T_2401 = _T_2399 == 64'h0; // @[BTB.scala 118:19:@2163.4]
  assign _T_2664 = _T_2399[0]; // @[OneHot.scala 39:40:@2357.4]
  assign _T_2665 = _T_2399[1]; // @[OneHot.scala 39:40:@2358.4]
  assign _T_2666 = _T_2399[2]; // @[OneHot.scala 39:40:@2359.4]
  assign _T_2667 = _T_2399[3]; // @[OneHot.scala 39:40:@2360.4]
  assign _T_2668 = _T_2399[4]; // @[OneHot.scala 39:40:@2361.4]
  assign _T_2669 = _T_2399[5]; // @[OneHot.scala 39:40:@2362.4]
  assign _T_2670 = _T_2399[6]; // @[OneHot.scala 39:40:@2363.4]
  assign _T_2671 = _T_2399[7]; // @[OneHot.scala 39:40:@2364.4]
  assign _T_2672 = _T_2399[8]; // @[OneHot.scala 39:40:@2365.4]
  assign _T_2673 = _T_2399[9]; // @[OneHot.scala 39:40:@2366.4]
  assign _T_2674 = _T_2399[10]; // @[OneHot.scala 39:40:@2367.4]
  assign _T_2675 = _T_2399[11]; // @[OneHot.scala 39:40:@2368.4]
  assign _T_2676 = _T_2399[12]; // @[OneHot.scala 39:40:@2369.4]
  assign _T_2677 = _T_2399[13]; // @[OneHot.scala 39:40:@2370.4]
  assign _T_2678 = _T_2399[14]; // @[OneHot.scala 39:40:@2371.4]
  assign _T_2679 = _T_2399[15]; // @[OneHot.scala 39:40:@2372.4]
  assign _T_2680 = _T_2399[16]; // @[OneHot.scala 39:40:@2373.4]
  assign _T_2681 = _T_2399[17]; // @[OneHot.scala 39:40:@2374.4]
  assign _T_2682 = _T_2399[18]; // @[OneHot.scala 39:40:@2375.4]
  assign _T_2683 = _T_2399[19]; // @[OneHot.scala 39:40:@2376.4]
  assign _T_2684 = _T_2399[20]; // @[OneHot.scala 39:40:@2377.4]
  assign _T_2685 = _T_2399[21]; // @[OneHot.scala 39:40:@2378.4]
  assign _T_2686 = _T_2399[22]; // @[OneHot.scala 39:40:@2379.4]
  assign _T_2687 = _T_2399[23]; // @[OneHot.scala 39:40:@2380.4]
  assign _T_2688 = _T_2399[24]; // @[OneHot.scala 39:40:@2381.4]
  assign _T_2689 = _T_2399[25]; // @[OneHot.scala 39:40:@2382.4]
  assign _T_2690 = _T_2399[26]; // @[OneHot.scala 39:40:@2383.4]
  assign _T_2691 = _T_2399[27]; // @[OneHot.scala 39:40:@2384.4]
  assign _T_2692 = _T_2399[28]; // @[OneHot.scala 39:40:@2385.4]
  assign _T_2693 = _T_2399[29]; // @[OneHot.scala 39:40:@2386.4]
  assign _T_2694 = _T_2399[30]; // @[OneHot.scala 39:40:@2387.4]
  assign _T_2695 = _T_2399[31]; // @[OneHot.scala 39:40:@2388.4]
  assign _T_2696 = _T_2399[32]; // @[OneHot.scala 39:40:@2389.4]
  assign _T_2697 = _T_2399[33]; // @[OneHot.scala 39:40:@2390.4]
  assign _T_2698 = _T_2399[34]; // @[OneHot.scala 39:40:@2391.4]
  assign _T_2699 = _T_2399[35]; // @[OneHot.scala 39:40:@2392.4]
  assign _T_2700 = _T_2399[36]; // @[OneHot.scala 39:40:@2393.4]
  assign _T_2701 = _T_2399[37]; // @[OneHot.scala 39:40:@2394.4]
  assign _T_2702 = _T_2399[38]; // @[OneHot.scala 39:40:@2395.4]
  assign _T_2703 = _T_2399[39]; // @[OneHot.scala 39:40:@2396.4]
  assign _T_2704 = _T_2399[40]; // @[OneHot.scala 39:40:@2397.4]
  assign _T_2705 = _T_2399[41]; // @[OneHot.scala 39:40:@2398.4]
  assign _T_2706 = _T_2399[42]; // @[OneHot.scala 39:40:@2399.4]
  assign _T_2707 = _T_2399[43]; // @[OneHot.scala 39:40:@2400.4]
  assign _T_2708 = _T_2399[44]; // @[OneHot.scala 39:40:@2401.4]
  assign _T_2709 = _T_2399[45]; // @[OneHot.scala 39:40:@2402.4]
  assign _T_2710 = _T_2399[46]; // @[OneHot.scala 39:40:@2403.4]
  assign _T_2711 = _T_2399[47]; // @[OneHot.scala 39:40:@2404.4]
  assign _T_2712 = _T_2399[48]; // @[OneHot.scala 39:40:@2405.4]
  assign _T_2713 = _T_2399[49]; // @[OneHot.scala 39:40:@2406.4]
  assign _T_2714 = _T_2399[50]; // @[OneHot.scala 39:40:@2407.4]
  assign _T_2715 = _T_2399[51]; // @[OneHot.scala 39:40:@2408.4]
  assign _T_2716 = _T_2399[52]; // @[OneHot.scala 39:40:@2409.4]
  assign _T_2717 = _T_2399[53]; // @[OneHot.scala 39:40:@2410.4]
  assign _T_2718 = _T_2399[54]; // @[OneHot.scala 39:40:@2411.4]
  assign _T_2719 = _T_2399[55]; // @[OneHot.scala 39:40:@2412.4]
  assign _T_2720 = _T_2399[56]; // @[OneHot.scala 39:40:@2413.4]
  assign _T_2721 = _T_2399[57]; // @[OneHot.scala 39:40:@2414.4]
  assign _T_2722 = _T_2399[58]; // @[OneHot.scala 39:40:@2415.4]
  assign _T_2723 = _T_2399[59]; // @[OneHot.scala 39:40:@2416.4]
  assign _T_2724 = _T_2399[60]; // @[OneHot.scala 39:40:@2417.4]
  assign _T_2725 = _T_2399[61]; // @[OneHot.scala 39:40:@2418.4]
  assign _T_2726 = _T_2399[62]; // @[OneHot.scala 39:40:@2419.4]
  assign _T_2792 = _T_2726 ? 6'h3e : 6'h3f; // @[Mux.scala 31:69:@2421.4]
  assign _T_2793 = _T_2725 ? 6'h3d : _T_2792; // @[Mux.scala 31:69:@2422.4]
  assign _T_2794 = _T_2724 ? 6'h3c : _T_2793; // @[Mux.scala 31:69:@2423.4]
  assign _T_2795 = _T_2723 ? 6'h3b : _T_2794; // @[Mux.scala 31:69:@2424.4]
  assign _T_2796 = _T_2722 ? 6'h3a : _T_2795; // @[Mux.scala 31:69:@2425.4]
  assign _T_2797 = _T_2721 ? 6'h39 : _T_2796; // @[Mux.scala 31:69:@2426.4]
  assign _T_2798 = _T_2720 ? 6'h38 : _T_2797; // @[Mux.scala 31:69:@2427.4]
  assign _T_2799 = _T_2719 ? 6'h37 : _T_2798; // @[Mux.scala 31:69:@2428.4]
  assign _T_2800 = _T_2718 ? 6'h36 : _T_2799; // @[Mux.scala 31:69:@2429.4]
  assign _T_2801 = _T_2717 ? 6'h35 : _T_2800; // @[Mux.scala 31:69:@2430.4]
  assign _T_2802 = _T_2716 ? 6'h34 : _T_2801; // @[Mux.scala 31:69:@2431.4]
  assign _T_2803 = _T_2715 ? 6'h33 : _T_2802; // @[Mux.scala 31:69:@2432.4]
  assign _T_2804 = _T_2714 ? 6'h32 : _T_2803; // @[Mux.scala 31:69:@2433.4]
  assign _T_2805 = _T_2713 ? 6'h31 : _T_2804; // @[Mux.scala 31:69:@2434.4]
  assign _T_2806 = _T_2712 ? 6'h30 : _T_2805; // @[Mux.scala 31:69:@2435.4]
  assign _T_2807 = _T_2711 ? 6'h2f : _T_2806; // @[Mux.scala 31:69:@2436.4]
  assign _T_2808 = _T_2710 ? 6'h2e : _T_2807; // @[Mux.scala 31:69:@2437.4]
  assign _T_2809 = _T_2709 ? 6'h2d : _T_2808; // @[Mux.scala 31:69:@2438.4]
  assign _T_2810 = _T_2708 ? 6'h2c : _T_2809; // @[Mux.scala 31:69:@2439.4]
  assign _T_2811 = _T_2707 ? 6'h2b : _T_2810; // @[Mux.scala 31:69:@2440.4]
  assign _T_2812 = _T_2706 ? 6'h2a : _T_2811; // @[Mux.scala 31:69:@2441.4]
  assign _T_2813 = _T_2705 ? 6'h29 : _T_2812; // @[Mux.scala 31:69:@2442.4]
  assign _T_2814 = _T_2704 ? 6'h28 : _T_2813; // @[Mux.scala 31:69:@2443.4]
  assign _T_2815 = _T_2703 ? 6'h27 : _T_2814; // @[Mux.scala 31:69:@2444.4]
  assign _T_2816 = _T_2702 ? 6'h26 : _T_2815; // @[Mux.scala 31:69:@2445.4]
  assign _T_2817 = _T_2701 ? 6'h25 : _T_2816; // @[Mux.scala 31:69:@2446.4]
  assign _T_2818 = _T_2700 ? 6'h24 : _T_2817; // @[Mux.scala 31:69:@2447.4]
  assign _T_2819 = _T_2699 ? 6'h23 : _T_2818; // @[Mux.scala 31:69:@2448.4]
  assign _T_2820 = _T_2698 ? 6'h22 : _T_2819; // @[Mux.scala 31:69:@2449.4]
  assign _T_2821 = _T_2697 ? 6'h21 : _T_2820; // @[Mux.scala 31:69:@2450.4]
  assign _T_2822 = _T_2696 ? 6'h20 : _T_2821; // @[Mux.scala 31:69:@2451.4]
  assign _T_2823 = _T_2695 ? 6'h1f : _T_2822; // @[Mux.scala 31:69:@2452.4]
  assign _T_2824 = _T_2694 ? 6'h1e : _T_2823; // @[Mux.scala 31:69:@2453.4]
  assign _T_2825 = _T_2693 ? 6'h1d : _T_2824; // @[Mux.scala 31:69:@2454.4]
  assign _T_2826 = _T_2692 ? 6'h1c : _T_2825; // @[Mux.scala 31:69:@2455.4]
  assign _T_2827 = _T_2691 ? 6'h1b : _T_2826; // @[Mux.scala 31:69:@2456.4]
  assign _T_2828 = _T_2690 ? 6'h1a : _T_2827; // @[Mux.scala 31:69:@2457.4]
  assign _T_2829 = _T_2689 ? 6'h19 : _T_2828; // @[Mux.scala 31:69:@2458.4]
  assign _T_2830 = _T_2688 ? 6'h18 : _T_2829; // @[Mux.scala 31:69:@2459.4]
  assign _T_2831 = _T_2687 ? 6'h17 : _T_2830; // @[Mux.scala 31:69:@2460.4]
  assign _T_2832 = _T_2686 ? 6'h16 : _T_2831; // @[Mux.scala 31:69:@2461.4]
  assign _T_2833 = _T_2685 ? 6'h15 : _T_2832; // @[Mux.scala 31:69:@2462.4]
  assign _T_2834 = _T_2684 ? 6'h14 : _T_2833; // @[Mux.scala 31:69:@2463.4]
  assign _T_2835 = _T_2683 ? 6'h13 : _T_2834; // @[Mux.scala 31:69:@2464.4]
  assign _T_2836 = _T_2682 ? 6'h12 : _T_2835; // @[Mux.scala 31:69:@2465.4]
  assign _T_2837 = _T_2681 ? 6'h11 : _T_2836; // @[Mux.scala 31:69:@2466.4]
  assign _T_2838 = _T_2680 ? 6'h10 : _T_2837; // @[Mux.scala 31:69:@2467.4]
  assign _T_2839 = _T_2679 ? 6'hf : _T_2838; // @[Mux.scala 31:69:@2468.4]
  assign _T_2840 = _T_2678 ? 6'he : _T_2839; // @[Mux.scala 31:69:@2469.4]
  assign _T_2841 = _T_2677 ? 6'hd : _T_2840; // @[Mux.scala 31:69:@2470.4]
  assign _T_2842 = _T_2676 ? 6'hc : _T_2841; // @[Mux.scala 31:69:@2471.4]
  assign _T_2843 = _T_2675 ? 6'hb : _T_2842; // @[Mux.scala 31:69:@2472.4]
  assign _T_2844 = _T_2674 ? 6'ha : _T_2843; // @[Mux.scala 31:69:@2473.4]
  assign _T_2845 = _T_2673 ? 6'h9 : _T_2844; // @[Mux.scala 31:69:@2474.4]
  assign _T_2846 = _T_2672 ? 6'h8 : _T_2845; // @[Mux.scala 31:69:@2475.4]
  assign _T_2847 = _T_2671 ? 6'h7 : _T_2846; // @[Mux.scala 31:69:@2476.4]
  assign _T_2848 = _T_2670 ? 6'h6 : _T_2847; // @[Mux.scala 31:69:@2477.4]
  assign _T_2849 = _T_2669 ? 6'h5 : _T_2848; // @[Mux.scala 31:69:@2478.4]
  assign _T_2850 = _T_2668 ? 6'h4 : _T_2849; // @[Mux.scala 31:69:@2479.4]
  assign _T_2851 = _T_2667 ? 6'h3 : _T_2850; // @[Mux.scala 31:69:@2480.4]
  assign _T_2852 = _T_2666 ? 6'h2 : _T_2851; // @[Mux.scala 31:69:@2481.4]
  assign _T_2853 = _T_2665 ? 6'h1 : _T_2852; // @[Mux.scala 31:69:@2482.4]
  assign _T_2854 = _T_2664 ? 6'h0 : _T_2853; // @[Mux.scala 31:69:@2483.4]
  assign _T_2855 = _T_2401 ? fb_reg_lfsr : _T_2854; // @[BTB.scala 118:8:@2484.4]
  assign fb_wire_bindex = _T_2106 ? _T_2137 : _T_2855; // @[BTB.scala 117:8:@2485.4]
  assign _GEN_0 = 6'h0 == fb_wire_bindex ? fb_reg_pc : btb_pc_0; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_1 = 6'h1 == fb_wire_bindex ? fb_reg_pc : btb_pc_1; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_2 = 6'h2 == fb_wire_bindex ? fb_reg_pc : btb_pc_2; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_3 = 6'h3 == fb_wire_bindex ? fb_reg_pc : btb_pc_3; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_4 = 6'h4 == fb_wire_bindex ? fb_reg_pc : btb_pc_4; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_5 = 6'h5 == fb_wire_bindex ? fb_reg_pc : btb_pc_5; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_6 = 6'h6 == fb_wire_bindex ? fb_reg_pc : btb_pc_6; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_7 = 6'h7 == fb_wire_bindex ? fb_reg_pc : btb_pc_7; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_8 = 6'h8 == fb_wire_bindex ? fb_reg_pc : btb_pc_8; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_9 = 6'h9 == fb_wire_bindex ? fb_reg_pc : btb_pc_9; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_10 = 6'ha == fb_wire_bindex ? fb_reg_pc : btb_pc_10; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_11 = 6'hb == fb_wire_bindex ? fb_reg_pc : btb_pc_11; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_12 = 6'hc == fb_wire_bindex ? fb_reg_pc : btb_pc_12; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_13 = 6'hd == fb_wire_bindex ? fb_reg_pc : btb_pc_13; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_14 = 6'he == fb_wire_bindex ? fb_reg_pc : btb_pc_14; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_15 = 6'hf == fb_wire_bindex ? fb_reg_pc : btb_pc_15; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_16 = 6'h10 == fb_wire_bindex ? fb_reg_pc : btb_pc_16; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_17 = 6'h11 == fb_wire_bindex ? fb_reg_pc : btb_pc_17; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_18 = 6'h12 == fb_wire_bindex ? fb_reg_pc : btb_pc_18; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_19 = 6'h13 == fb_wire_bindex ? fb_reg_pc : btb_pc_19; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_20 = 6'h14 == fb_wire_bindex ? fb_reg_pc : btb_pc_20; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_21 = 6'h15 == fb_wire_bindex ? fb_reg_pc : btb_pc_21; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_22 = 6'h16 == fb_wire_bindex ? fb_reg_pc : btb_pc_22; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_23 = 6'h17 == fb_wire_bindex ? fb_reg_pc : btb_pc_23; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_24 = 6'h18 == fb_wire_bindex ? fb_reg_pc : btb_pc_24; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_25 = 6'h19 == fb_wire_bindex ? fb_reg_pc : btb_pc_25; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_26 = 6'h1a == fb_wire_bindex ? fb_reg_pc : btb_pc_26; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_27 = 6'h1b == fb_wire_bindex ? fb_reg_pc : btb_pc_27; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_28 = 6'h1c == fb_wire_bindex ? fb_reg_pc : btb_pc_28; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_29 = 6'h1d == fb_wire_bindex ? fb_reg_pc : btb_pc_29; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_30 = 6'h1e == fb_wire_bindex ? fb_reg_pc : btb_pc_30; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_31 = 6'h1f == fb_wire_bindex ? fb_reg_pc : btb_pc_31; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_32 = 6'h20 == fb_wire_bindex ? fb_reg_pc : btb_pc_32; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_33 = 6'h21 == fb_wire_bindex ? fb_reg_pc : btb_pc_33; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_34 = 6'h22 == fb_wire_bindex ? fb_reg_pc : btb_pc_34; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_35 = 6'h23 == fb_wire_bindex ? fb_reg_pc : btb_pc_35; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_36 = 6'h24 == fb_wire_bindex ? fb_reg_pc : btb_pc_36; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_37 = 6'h25 == fb_wire_bindex ? fb_reg_pc : btb_pc_37; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_38 = 6'h26 == fb_wire_bindex ? fb_reg_pc : btb_pc_38; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_39 = 6'h27 == fb_wire_bindex ? fb_reg_pc : btb_pc_39; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_40 = 6'h28 == fb_wire_bindex ? fb_reg_pc : btb_pc_40; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_41 = 6'h29 == fb_wire_bindex ? fb_reg_pc : btb_pc_41; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_42 = 6'h2a == fb_wire_bindex ? fb_reg_pc : btb_pc_42; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_43 = 6'h2b == fb_wire_bindex ? fb_reg_pc : btb_pc_43; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_44 = 6'h2c == fb_wire_bindex ? fb_reg_pc : btb_pc_44; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_45 = 6'h2d == fb_wire_bindex ? fb_reg_pc : btb_pc_45; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_46 = 6'h2e == fb_wire_bindex ? fb_reg_pc : btb_pc_46; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_47 = 6'h2f == fb_wire_bindex ? fb_reg_pc : btb_pc_47; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_48 = 6'h30 == fb_wire_bindex ? fb_reg_pc : btb_pc_48; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_49 = 6'h31 == fb_wire_bindex ? fb_reg_pc : btb_pc_49; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_50 = 6'h32 == fb_wire_bindex ? fb_reg_pc : btb_pc_50; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_51 = 6'h33 == fb_wire_bindex ? fb_reg_pc : btb_pc_51; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_52 = 6'h34 == fb_wire_bindex ? fb_reg_pc : btb_pc_52; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_53 = 6'h35 == fb_wire_bindex ? fb_reg_pc : btb_pc_53; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_54 = 6'h36 == fb_wire_bindex ? fb_reg_pc : btb_pc_54; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_55 = 6'h37 == fb_wire_bindex ? fb_reg_pc : btb_pc_55; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_56 = 6'h38 == fb_wire_bindex ? fb_reg_pc : btb_pc_56; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_57 = 6'h39 == fb_wire_bindex ? fb_reg_pc : btb_pc_57; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_58 = 6'h3a == fb_wire_bindex ? fb_reg_pc : btb_pc_58; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_59 = 6'h3b == fb_wire_bindex ? fb_reg_pc : btb_pc_59; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_60 = 6'h3c == fb_wire_bindex ? fb_reg_pc : btb_pc_60; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_61 = 6'h3d == fb_wire_bindex ? fb_reg_pc : btb_pc_61; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_62 = 6'h3e == fb_wire_bindex ? fb_reg_pc : btb_pc_62; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_63 = 6'h3f == fb_wire_bindex ? fb_reg_pc : btb_pc_63; // @[BTB.scala 124:34:@2489.8]
  assign _GEN_64 = 6'h0 == fb_wire_bindex ? fb_reg_target : btb_target_0; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_65 = 6'h1 == fb_wire_bindex ? fb_reg_target : btb_target_1; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_66 = 6'h2 == fb_wire_bindex ? fb_reg_target : btb_target_2; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_67 = 6'h3 == fb_wire_bindex ? fb_reg_target : btb_target_3; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_68 = 6'h4 == fb_wire_bindex ? fb_reg_target : btb_target_4; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_69 = 6'h5 == fb_wire_bindex ? fb_reg_target : btb_target_5; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_70 = 6'h6 == fb_wire_bindex ? fb_reg_target : btb_target_6; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_71 = 6'h7 == fb_wire_bindex ? fb_reg_target : btb_target_7; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_72 = 6'h8 == fb_wire_bindex ? fb_reg_target : btb_target_8; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_73 = 6'h9 == fb_wire_bindex ? fb_reg_target : btb_target_9; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_74 = 6'ha == fb_wire_bindex ? fb_reg_target : btb_target_10; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_75 = 6'hb == fb_wire_bindex ? fb_reg_target : btb_target_11; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_76 = 6'hc == fb_wire_bindex ? fb_reg_target : btb_target_12; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_77 = 6'hd == fb_wire_bindex ? fb_reg_target : btb_target_13; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_78 = 6'he == fb_wire_bindex ? fb_reg_target : btb_target_14; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_79 = 6'hf == fb_wire_bindex ? fb_reg_target : btb_target_15; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_80 = 6'h10 == fb_wire_bindex ? fb_reg_target : btb_target_16; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_81 = 6'h11 == fb_wire_bindex ? fb_reg_target : btb_target_17; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_82 = 6'h12 == fb_wire_bindex ? fb_reg_target : btb_target_18; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_83 = 6'h13 == fb_wire_bindex ? fb_reg_target : btb_target_19; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_84 = 6'h14 == fb_wire_bindex ? fb_reg_target : btb_target_20; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_85 = 6'h15 == fb_wire_bindex ? fb_reg_target : btb_target_21; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_86 = 6'h16 == fb_wire_bindex ? fb_reg_target : btb_target_22; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_87 = 6'h17 == fb_wire_bindex ? fb_reg_target : btb_target_23; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_88 = 6'h18 == fb_wire_bindex ? fb_reg_target : btb_target_24; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_89 = 6'h19 == fb_wire_bindex ? fb_reg_target : btb_target_25; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_90 = 6'h1a == fb_wire_bindex ? fb_reg_target : btb_target_26; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_91 = 6'h1b == fb_wire_bindex ? fb_reg_target : btb_target_27; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_92 = 6'h1c == fb_wire_bindex ? fb_reg_target : btb_target_28; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_93 = 6'h1d == fb_wire_bindex ? fb_reg_target : btb_target_29; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_94 = 6'h1e == fb_wire_bindex ? fb_reg_target : btb_target_30; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_95 = 6'h1f == fb_wire_bindex ? fb_reg_target : btb_target_31; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_96 = 6'h20 == fb_wire_bindex ? fb_reg_target : btb_target_32; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_97 = 6'h21 == fb_wire_bindex ? fb_reg_target : btb_target_33; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_98 = 6'h22 == fb_wire_bindex ? fb_reg_target : btb_target_34; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_99 = 6'h23 == fb_wire_bindex ? fb_reg_target : btb_target_35; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_100 = 6'h24 == fb_wire_bindex ? fb_reg_target : btb_target_36; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_101 = 6'h25 == fb_wire_bindex ? fb_reg_target : btb_target_37; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_102 = 6'h26 == fb_wire_bindex ? fb_reg_target : btb_target_38; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_103 = 6'h27 == fb_wire_bindex ? fb_reg_target : btb_target_39; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_104 = 6'h28 == fb_wire_bindex ? fb_reg_target : btb_target_40; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_105 = 6'h29 == fb_wire_bindex ? fb_reg_target : btb_target_41; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_106 = 6'h2a == fb_wire_bindex ? fb_reg_target : btb_target_42; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_107 = 6'h2b == fb_wire_bindex ? fb_reg_target : btb_target_43; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_108 = 6'h2c == fb_wire_bindex ? fb_reg_target : btb_target_44; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_109 = 6'h2d == fb_wire_bindex ? fb_reg_target : btb_target_45; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_110 = 6'h2e == fb_wire_bindex ? fb_reg_target : btb_target_46; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_111 = 6'h2f == fb_wire_bindex ? fb_reg_target : btb_target_47; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_112 = 6'h30 == fb_wire_bindex ? fb_reg_target : btb_target_48; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_113 = 6'h31 == fb_wire_bindex ? fb_reg_target : btb_target_49; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_114 = 6'h32 == fb_wire_bindex ? fb_reg_target : btb_target_50; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_115 = 6'h33 == fb_wire_bindex ? fb_reg_target : btb_target_51; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_116 = 6'h34 == fb_wire_bindex ? fb_reg_target : btb_target_52; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_117 = 6'h35 == fb_wire_bindex ? fb_reg_target : btb_target_53; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_118 = 6'h36 == fb_wire_bindex ? fb_reg_target : btb_target_54; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_119 = 6'h37 == fb_wire_bindex ? fb_reg_target : btb_target_55; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_120 = 6'h38 == fb_wire_bindex ? fb_reg_target : btb_target_56; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_121 = 6'h39 == fb_wire_bindex ? fb_reg_target : btb_target_57; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_122 = 6'h3a == fb_wire_bindex ? fb_reg_target : btb_target_58; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_123 = 6'h3b == fb_wire_bindex ? fb_reg_target : btb_target_59; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_124 = 6'h3c == fb_wire_bindex ? fb_reg_target : btb_target_60; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_125 = 6'h3d == fb_wire_bindex ? fb_reg_target : btb_target_61; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_126 = 6'h3e == fb_wire_bindex ? fb_reg_target : btb_target_62; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_127 = 6'h3f == fb_wire_bindex ? fb_reg_target : btb_target_63; // @[BTB.scala 125:34:@2490.8]
  assign _GEN_128 = 6'h0 == fb_wire_bindex ? fb_reg_btype : btb_btype_0; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_129 = 6'h1 == fb_wire_bindex ? fb_reg_btype : btb_btype_1; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_130 = 6'h2 == fb_wire_bindex ? fb_reg_btype : btb_btype_2; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_131 = 6'h3 == fb_wire_bindex ? fb_reg_btype : btb_btype_3; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_132 = 6'h4 == fb_wire_bindex ? fb_reg_btype : btb_btype_4; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_133 = 6'h5 == fb_wire_bindex ? fb_reg_btype : btb_btype_5; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_134 = 6'h6 == fb_wire_bindex ? fb_reg_btype : btb_btype_6; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_135 = 6'h7 == fb_wire_bindex ? fb_reg_btype : btb_btype_7; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_136 = 6'h8 == fb_wire_bindex ? fb_reg_btype : btb_btype_8; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_137 = 6'h9 == fb_wire_bindex ? fb_reg_btype : btb_btype_9; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_138 = 6'ha == fb_wire_bindex ? fb_reg_btype : btb_btype_10; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_139 = 6'hb == fb_wire_bindex ? fb_reg_btype : btb_btype_11; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_140 = 6'hc == fb_wire_bindex ? fb_reg_btype : btb_btype_12; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_141 = 6'hd == fb_wire_bindex ? fb_reg_btype : btb_btype_13; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_142 = 6'he == fb_wire_bindex ? fb_reg_btype : btb_btype_14; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_143 = 6'hf == fb_wire_bindex ? fb_reg_btype : btb_btype_15; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_144 = 6'h10 == fb_wire_bindex ? fb_reg_btype : btb_btype_16; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_145 = 6'h11 == fb_wire_bindex ? fb_reg_btype : btb_btype_17; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_146 = 6'h12 == fb_wire_bindex ? fb_reg_btype : btb_btype_18; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_147 = 6'h13 == fb_wire_bindex ? fb_reg_btype : btb_btype_19; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_148 = 6'h14 == fb_wire_bindex ? fb_reg_btype : btb_btype_20; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_149 = 6'h15 == fb_wire_bindex ? fb_reg_btype : btb_btype_21; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_150 = 6'h16 == fb_wire_bindex ? fb_reg_btype : btb_btype_22; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_151 = 6'h17 == fb_wire_bindex ? fb_reg_btype : btb_btype_23; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_152 = 6'h18 == fb_wire_bindex ? fb_reg_btype : btb_btype_24; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_153 = 6'h19 == fb_wire_bindex ? fb_reg_btype : btb_btype_25; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_154 = 6'h1a == fb_wire_bindex ? fb_reg_btype : btb_btype_26; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_155 = 6'h1b == fb_wire_bindex ? fb_reg_btype : btb_btype_27; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_156 = 6'h1c == fb_wire_bindex ? fb_reg_btype : btb_btype_28; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_157 = 6'h1d == fb_wire_bindex ? fb_reg_btype : btb_btype_29; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_158 = 6'h1e == fb_wire_bindex ? fb_reg_btype : btb_btype_30; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_159 = 6'h1f == fb_wire_bindex ? fb_reg_btype : btb_btype_31; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_160 = 6'h20 == fb_wire_bindex ? fb_reg_btype : btb_btype_32; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_161 = 6'h21 == fb_wire_bindex ? fb_reg_btype : btb_btype_33; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_162 = 6'h22 == fb_wire_bindex ? fb_reg_btype : btb_btype_34; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_163 = 6'h23 == fb_wire_bindex ? fb_reg_btype : btb_btype_35; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_164 = 6'h24 == fb_wire_bindex ? fb_reg_btype : btb_btype_36; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_165 = 6'h25 == fb_wire_bindex ? fb_reg_btype : btb_btype_37; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_166 = 6'h26 == fb_wire_bindex ? fb_reg_btype : btb_btype_38; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_167 = 6'h27 == fb_wire_bindex ? fb_reg_btype : btb_btype_39; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_168 = 6'h28 == fb_wire_bindex ? fb_reg_btype : btb_btype_40; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_169 = 6'h29 == fb_wire_bindex ? fb_reg_btype : btb_btype_41; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_170 = 6'h2a == fb_wire_bindex ? fb_reg_btype : btb_btype_42; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_171 = 6'h2b == fb_wire_bindex ? fb_reg_btype : btb_btype_43; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_172 = 6'h2c == fb_wire_bindex ? fb_reg_btype : btb_btype_44; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_173 = 6'h2d == fb_wire_bindex ? fb_reg_btype : btb_btype_45; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_174 = 6'h2e == fb_wire_bindex ? fb_reg_btype : btb_btype_46; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_175 = 6'h2f == fb_wire_bindex ? fb_reg_btype : btb_btype_47; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_176 = 6'h30 == fb_wire_bindex ? fb_reg_btype : btb_btype_48; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_177 = 6'h31 == fb_wire_bindex ? fb_reg_btype : btb_btype_49; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_178 = 6'h32 == fb_wire_bindex ? fb_reg_btype : btb_btype_50; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_179 = 6'h33 == fb_wire_bindex ? fb_reg_btype : btb_btype_51; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_180 = 6'h34 == fb_wire_bindex ? fb_reg_btype : btb_btype_52; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_181 = 6'h35 == fb_wire_bindex ? fb_reg_btype : btb_btype_53; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_182 = 6'h36 == fb_wire_bindex ? fb_reg_btype : btb_btype_54; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_183 = 6'h37 == fb_wire_bindex ? fb_reg_btype : btb_btype_55; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_184 = 6'h38 == fb_wire_bindex ? fb_reg_btype : btb_btype_56; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_185 = 6'h39 == fb_wire_bindex ? fb_reg_btype : btb_btype_57; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_186 = 6'h3a == fb_wire_bindex ? fb_reg_btype : btb_btype_58; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_187 = 6'h3b == fb_wire_bindex ? fb_reg_btype : btb_btype_59; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_188 = 6'h3c == fb_wire_bindex ? fb_reg_btype : btb_btype_60; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_189 = 6'h3d == fb_wire_bindex ? fb_reg_btype : btb_btype_61; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_190 = 6'h3e == fb_wire_bindex ? fb_reg_btype : btb_btype_62; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_191 = 6'h3f == fb_wire_bindex ? fb_reg_btype : btb_btype_63; // @[BTB.scala 126:34:@2491.8]
  assign _GEN_192 = fb_reg_redirect ? _GEN_0 : btb_pc_0; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_193 = fb_reg_redirect ? _GEN_1 : btb_pc_1; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_194 = fb_reg_redirect ? _GEN_2 : btb_pc_2; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_195 = fb_reg_redirect ? _GEN_3 : btb_pc_3; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_196 = fb_reg_redirect ? _GEN_4 : btb_pc_4; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_197 = fb_reg_redirect ? _GEN_5 : btb_pc_5; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_198 = fb_reg_redirect ? _GEN_6 : btb_pc_6; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_199 = fb_reg_redirect ? _GEN_7 : btb_pc_7; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_200 = fb_reg_redirect ? _GEN_8 : btb_pc_8; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_201 = fb_reg_redirect ? _GEN_9 : btb_pc_9; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_202 = fb_reg_redirect ? _GEN_10 : btb_pc_10; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_203 = fb_reg_redirect ? _GEN_11 : btb_pc_11; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_204 = fb_reg_redirect ? _GEN_12 : btb_pc_12; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_205 = fb_reg_redirect ? _GEN_13 : btb_pc_13; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_206 = fb_reg_redirect ? _GEN_14 : btb_pc_14; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_207 = fb_reg_redirect ? _GEN_15 : btb_pc_15; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_208 = fb_reg_redirect ? _GEN_16 : btb_pc_16; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_209 = fb_reg_redirect ? _GEN_17 : btb_pc_17; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_210 = fb_reg_redirect ? _GEN_18 : btb_pc_18; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_211 = fb_reg_redirect ? _GEN_19 : btb_pc_19; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_212 = fb_reg_redirect ? _GEN_20 : btb_pc_20; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_213 = fb_reg_redirect ? _GEN_21 : btb_pc_21; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_214 = fb_reg_redirect ? _GEN_22 : btb_pc_22; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_215 = fb_reg_redirect ? _GEN_23 : btb_pc_23; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_216 = fb_reg_redirect ? _GEN_24 : btb_pc_24; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_217 = fb_reg_redirect ? _GEN_25 : btb_pc_25; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_218 = fb_reg_redirect ? _GEN_26 : btb_pc_26; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_219 = fb_reg_redirect ? _GEN_27 : btb_pc_27; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_220 = fb_reg_redirect ? _GEN_28 : btb_pc_28; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_221 = fb_reg_redirect ? _GEN_29 : btb_pc_29; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_222 = fb_reg_redirect ? _GEN_30 : btb_pc_30; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_223 = fb_reg_redirect ? _GEN_31 : btb_pc_31; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_224 = fb_reg_redirect ? _GEN_32 : btb_pc_32; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_225 = fb_reg_redirect ? _GEN_33 : btb_pc_33; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_226 = fb_reg_redirect ? _GEN_34 : btb_pc_34; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_227 = fb_reg_redirect ? _GEN_35 : btb_pc_35; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_228 = fb_reg_redirect ? _GEN_36 : btb_pc_36; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_229 = fb_reg_redirect ? _GEN_37 : btb_pc_37; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_230 = fb_reg_redirect ? _GEN_38 : btb_pc_38; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_231 = fb_reg_redirect ? _GEN_39 : btb_pc_39; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_232 = fb_reg_redirect ? _GEN_40 : btb_pc_40; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_233 = fb_reg_redirect ? _GEN_41 : btb_pc_41; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_234 = fb_reg_redirect ? _GEN_42 : btb_pc_42; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_235 = fb_reg_redirect ? _GEN_43 : btb_pc_43; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_236 = fb_reg_redirect ? _GEN_44 : btb_pc_44; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_237 = fb_reg_redirect ? _GEN_45 : btb_pc_45; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_238 = fb_reg_redirect ? _GEN_46 : btb_pc_46; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_239 = fb_reg_redirect ? _GEN_47 : btb_pc_47; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_240 = fb_reg_redirect ? _GEN_48 : btb_pc_48; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_241 = fb_reg_redirect ? _GEN_49 : btb_pc_49; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_242 = fb_reg_redirect ? _GEN_50 : btb_pc_50; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_243 = fb_reg_redirect ? _GEN_51 : btb_pc_51; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_244 = fb_reg_redirect ? _GEN_52 : btb_pc_52; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_245 = fb_reg_redirect ? _GEN_53 : btb_pc_53; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_246 = fb_reg_redirect ? _GEN_54 : btb_pc_54; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_247 = fb_reg_redirect ? _GEN_55 : btb_pc_55; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_248 = fb_reg_redirect ? _GEN_56 : btb_pc_56; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_249 = fb_reg_redirect ? _GEN_57 : btb_pc_57; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_250 = fb_reg_redirect ? _GEN_58 : btb_pc_58; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_251 = fb_reg_redirect ? _GEN_59 : btb_pc_59; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_252 = fb_reg_redirect ? _GEN_60 : btb_pc_60; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_253 = fb_reg_redirect ? _GEN_61 : btb_pc_61; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_254 = fb_reg_redirect ? _GEN_62 : btb_pc_62; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_255 = fb_reg_redirect ? _GEN_63 : btb_pc_63; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_256 = fb_reg_redirect ? _GEN_64 : btb_target_0; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_257 = fb_reg_redirect ? _GEN_65 : btb_target_1; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_258 = fb_reg_redirect ? _GEN_66 : btb_target_2; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_259 = fb_reg_redirect ? _GEN_67 : btb_target_3; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_260 = fb_reg_redirect ? _GEN_68 : btb_target_4; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_261 = fb_reg_redirect ? _GEN_69 : btb_target_5; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_262 = fb_reg_redirect ? _GEN_70 : btb_target_6; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_263 = fb_reg_redirect ? _GEN_71 : btb_target_7; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_264 = fb_reg_redirect ? _GEN_72 : btb_target_8; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_265 = fb_reg_redirect ? _GEN_73 : btb_target_9; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_266 = fb_reg_redirect ? _GEN_74 : btb_target_10; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_267 = fb_reg_redirect ? _GEN_75 : btb_target_11; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_268 = fb_reg_redirect ? _GEN_76 : btb_target_12; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_269 = fb_reg_redirect ? _GEN_77 : btb_target_13; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_270 = fb_reg_redirect ? _GEN_78 : btb_target_14; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_271 = fb_reg_redirect ? _GEN_79 : btb_target_15; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_272 = fb_reg_redirect ? _GEN_80 : btb_target_16; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_273 = fb_reg_redirect ? _GEN_81 : btb_target_17; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_274 = fb_reg_redirect ? _GEN_82 : btb_target_18; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_275 = fb_reg_redirect ? _GEN_83 : btb_target_19; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_276 = fb_reg_redirect ? _GEN_84 : btb_target_20; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_277 = fb_reg_redirect ? _GEN_85 : btb_target_21; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_278 = fb_reg_redirect ? _GEN_86 : btb_target_22; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_279 = fb_reg_redirect ? _GEN_87 : btb_target_23; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_280 = fb_reg_redirect ? _GEN_88 : btb_target_24; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_281 = fb_reg_redirect ? _GEN_89 : btb_target_25; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_282 = fb_reg_redirect ? _GEN_90 : btb_target_26; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_283 = fb_reg_redirect ? _GEN_91 : btb_target_27; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_284 = fb_reg_redirect ? _GEN_92 : btb_target_28; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_285 = fb_reg_redirect ? _GEN_93 : btb_target_29; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_286 = fb_reg_redirect ? _GEN_94 : btb_target_30; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_287 = fb_reg_redirect ? _GEN_95 : btb_target_31; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_288 = fb_reg_redirect ? _GEN_96 : btb_target_32; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_289 = fb_reg_redirect ? _GEN_97 : btb_target_33; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_290 = fb_reg_redirect ? _GEN_98 : btb_target_34; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_291 = fb_reg_redirect ? _GEN_99 : btb_target_35; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_292 = fb_reg_redirect ? _GEN_100 : btb_target_36; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_293 = fb_reg_redirect ? _GEN_101 : btb_target_37; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_294 = fb_reg_redirect ? _GEN_102 : btb_target_38; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_295 = fb_reg_redirect ? _GEN_103 : btb_target_39; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_296 = fb_reg_redirect ? _GEN_104 : btb_target_40; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_297 = fb_reg_redirect ? _GEN_105 : btb_target_41; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_298 = fb_reg_redirect ? _GEN_106 : btb_target_42; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_299 = fb_reg_redirect ? _GEN_107 : btb_target_43; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_300 = fb_reg_redirect ? _GEN_108 : btb_target_44; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_301 = fb_reg_redirect ? _GEN_109 : btb_target_45; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_302 = fb_reg_redirect ? _GEN_110 : btb_target_46; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_303 = fb_reg_redirect ? _GEN_111 : btb_target_47; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_304 = fb_reg_redirect ? _GEN_112 : btb_target_48; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_305 = fb_reg_redirect ? _GEN_113 : btb_target_49; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_306 = fb_reg_redirect ? _GEN_114 : btb_target_50; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_307 = fb_reg_redirect ? _GEN_115 : btb_target_51; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_308 = fb_reg_redirect ? _GEN_116 : btb_target_52; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_309 = fb_reg_redirect ? _GEN_117 : btb_target_53; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_310 = fb_reg_redirect ? _GEN_118 : btb_target_54; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_311 = fb_reg_redirect ? _GEN_119 : btb_target_55; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_312 = fb_reg_redirect ? _GEN_120 : btb_target_56; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_313 = fb_reg_redirect ? _GEN_121 : btb_target_57; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_314 = fb_reg_redirect ? _GEN_122 : btb_target_58; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_315 = fb_reg_redirect ? _GEN_123 : btb_target_59; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_316 = fb_reg_redirect ? _GEN_124 : btb_target_60; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_317 = fb_reg_redirect ? _GEN_125 : btb_target_61; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_318 = fb_reg_redirect ? _GEN_126 : btb_target_62; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_319 = fb_reg_redirect ? _GEN_127 : btb_target_63; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_320 = fb_reg_redirect ? _GEN_128 : btb_btype_0; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_321 = fb_reg_redirect ? _GEN_129 : btb_btype_1; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_322 = fb_reg_redirect ? _GEN_130 : btb_btype_2; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_323 = fb_reg_redirect ? _GEN_131 : btb_btype_3; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_324 = fb_reg_redirect ? _GEN_132 : btb_btype_4; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_325 = fb_reg_redirect ? _GEN_133 : btb_btype_5; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_326 = fb_reg_redirect ? _GEN_134 : btb_btype_6; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_327 = fb_reg_redirect ? _GEN_135 : btb_btype_7; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_328 = fb_reg_redirect ? _GEN_136 : btb_btype_8; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_329 = fb_reg_redirect ? _GEN_137 : btb_btype_9; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_330 = fb_reg_redirect ? _GEN_138 : btb_btype_10; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_331 = fb_reg_redirect ? _GEN_139 : btb_btype_11; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_332 = fb_reg_redirect ? _GEN_140 : btb_btype_12; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_333 = fb_reg_redirect ? _GEN_141 : btb_btype_13; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_334 = fb_reg_redirect ? _GEN_142 : btb_btype_14; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_335 = fb_reg_redirect ? _GEN_143 : btb_btype_15; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_336 = fb_reg_redirect ? _GEN_144 : btb_btype_16; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_337 = fb_reg_redirect ? _GEN_145 : btb_btype_17; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_338 = fb_reg_redirect ? _GEN_146 : btb_btype_18; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_339 = fb_reg_redirect ? _GEN_147 : btb_btype_19; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_340 = fb_reg_redirect ? _GEN_148 : btb_btype_20; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_341 = fb_reg_redirect ? _GEN_149 : btb_btype_21; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_342 = fb_reg_redirect ? _GEN_150 : btb_btype_22; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_343 = fb_reg_redirect ? _GEN_151 : btb_btype_23; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_344 = fb_reg_redirect ? _GEN_152 : btb_btype_24; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_345 = fb_reg_redirect ? _GEN_153 : btb_btype_25; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_346 = fb_reg_redirect ? _GEN_154 : btb_btype_26; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_347 = fb_reg_redirect ? _GEN_155 : btb_btype_27; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_348 = fb_reg_redirect ? _GEN_156 : btb_btype_28; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_349 = fb_reg_redirect ? _GEN_157 : btb_btype_29; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_350 = fb_reg_redirect ? _GEN_158 : btb_btype_30; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_351 = fb_reg_redirect ? _GEN_159 : btb_btype_31; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_352 = fb_reg_redirect ? _GEN_160 : btb_btype_32; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_353 = fb_reg_redirect ? _GEN_161 : btb_btype_33; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_354 = fb_reg_redirect ? _GEN_162 : btb_btype_34; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_355 = fb_reg_redirect ? _GEN_163 : btb_btype_35; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_356 = fb_reg_redirect ? _GEN_164 : btb_btype_36; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_357 = fb_reg_redirect ? _GEN_165 : btb_btype_37; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_358 = fb_reg_redirect ? _GEN_166 : btb_btype_38; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_359 = fb_reg_redirect ? _GEN_167 : btb_btype_39; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_360 = fb_reg_redirect ? _GEN_168 : btb_btype_40; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_361 = fb_reg_redirect ? _GEN_169 : btb_btype_41; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_362 = fb_reg_redirect ? _GEN_170 : btb_btype_42; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_363 = fb_reg_redirect ? _GEN_171 : btb_btype_43; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_364 = fb_reg_redirect ? _GEN_172 : btb_btype_44; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_365 = fb_reg_redirect ? _GEN_173 : btb_btype_45; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_366 = fb_reg_redirect ? _GEN_174 : btb_btype_46; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_367 = fb_reg_redirect ? _GEN_175 : btb_btype_47; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_368 = fb_reg_redirect ? _GEN_176 : btb_btype_48; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_369 = fb_reg_redirect ? _GEN_177 : btb_btype_49; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_370 = fb_reg_redirect ? _GEN_178 : btb_btype_50; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_371 = fb_reg_redirect ? _GEN_179 : btb_btype_51; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_372 = fb_reg_redirect ? _GEN_180 : btb_btype_52; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_373 = fb_reg_redirect ? _GEN_181 : btb_btype_53; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_374 = fb_reg_redirect ? _GEN_182 : btb_btype_54; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_375 = fb_reg_redirect ? _GEN_183 : btb_btype_55; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_376 = fb_reg_redirect ? _GEN_184 : btb_btype_56; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_377 = fb_reg_redirect ? _GEN_185 : btb_btype_57; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_378 = fb_reg_redirect ? _GEN_186 : btb_btype_58; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_379 = fb_reg_redirect ? _GEN_187 : btb_btype_59; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_380 = fb_reg_redirect ? _GEN_188 : btb_btype_60; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_381 = fb_reg_redirect ? _GEN_189 : btb_btype_61; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_382 = fb_reg_redirect ? _GEN_190 : btb_btype_62; // @[BTB.scala 123:28:@2488.6]
  assign _GEN_383 = fb_reg_redirect ? _GEN_191 : btb_btype_63; // @[BTB.scala 123:28:@2488.6]
  assign _T_2858 = fb_reg_btype == 2'h2; // @[BTB.scala 128:24:@2493.6]
  assign _T_2862 = fb_wire_hcount != 2'h0; // @[BTB.scala 51:42:@2498.12]
  assign _T_2863 = fb_wire_hcount[1]; // @[BTB.scala 51:49:@2499.12]
  assign _T_2864 = fb_wire_hcount[0]; // @[BTB.scala 51:58:@2500.12]
  assign _T_2866 = _T_2864 == 1'h0; // @[BTB.scala 51:56:@2501.12]
  assign _T_2867 = _T_2863 | _T_2866; // @[BTB.scala 51:53:@2502.12]
  assign _T_2868 = {_T_2862,_T_2867}; // @[Cat.scala 30:58:@2503.12]
  assign _GEN_384 = 6'h0 == fb_wire_bindex ? _T_2868 : btb_hcount_0; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_385 = 6'h1 == fb_wire_bindex ? _T_2868 : btb_hcount_1; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_386 = 6'h2 == fb_wire_bindex ? _T_2868 : btb_hcount_2; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_387 = 6'h3 == fb_wire_bindex ? _T_2868 : btb_hcount_3; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_388 = 6'h4 == fb_wire_bindex ? _T_2868 : btb_hcount_4; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_389 = 6'h5 == fb_wire_bindex ? _T_2868 : btb_hcount_5; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_390 = 6'h6 == fb_wire_bindex ? _T_2868 : btb_hcount_6; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_391 = 6'h7 == fb_wire_bindex ? _T_2868 : btb_hcount_7; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_392 = 6'h8 == fb_wire_bindex ? _T_2868 : btb_hcount_8; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_393 = 6'h9 == fb_wire_bindex ? _T_2868 : btb_hcount_9; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_394 = 6'ha == fb_wire_bindex ? _T_2868 : btb_hcount_10; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_395 = 6'hb == fb_wire_bindex ? _T_2868 : btb_hcount_11; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_396 = 6'hc == fb_wire_bindex ? _T_2868 : btb_hcount_12; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_397 = 6'hd == fb_wire_bindex ? _T_2868 : btb_hcount_13; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_398 = 6'he == fb_wire_bindex ? _T_2868 : btb_hcount_14; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_399 = 6'hf == fb_wire_bindex ? _T_2868 : btb_hcount_15; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_400 = 6'h10 == fb_wire_bindex ? _T_2868 : btb_hcount_16; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_401 = 6'h11 == fb_wire_bindex ? _T_2868 : btb_hcount_17; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_402 = 6'h12 == fb_wire_bindex ? _T_2868 : btb_hcount_18; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_403 = 6'h13 == fb_wire_bindex ? _T_2868 : btb_hcount_19; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_404 = 6'h14 == fb_wire_bindex ? _T_2868 : btb_hcount_20; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_405 = 6'h15 == fb_wire_bindex ? _T_2868 : btb_hcount_21; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_406 = 6'h16 == fb_wire_bindex ? _T_2868 : btb_hcount_22; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_407 = 6'h17 == fb_wire_bindex ? _T_2868 : btb_hcount_23; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_408 = 6'h18 == fb_wire_bindex ? _T_2868 : btb_hcount_24; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_409 = 6'h19 == fb_wire_bindex ? _T_2868 : btb_hcount_25; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_410 = 6'h1a == fb_wire_bindex ? _T_2868 : btb_hcount_26; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_411 = 6'h1b == fb_wire_bindex ? _T_2868 : btb_hcount_27; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_412 = 6'h1c == fb_wire_bindex ? _T_2868 : btb_hcount_28; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_413 = 6'h1d == fb_wire_bindex ? _T_2868 : btb_hcount_29; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_414 = 6'h1e == fb_wire_bindex ? _T_2868 : btb_hcount_30; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_415 = 6'h1f == fb_wire_bindex ? _T_2868 : btb_hcount_31; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_416 = 6'h20 == fb_wire_bindex ? _T_2868 : btb_hcount_32; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_417 = 6'h21 == fb_wire_bindex ? _T_2868 : btb_hcount_33; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_418 = 6'h22 == fb_wire_bindex ? _T_2868 : btb_hcount_34; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_419 = 6'h23 == fb_wire_bindex ? _T_2868 : btb_hcount_35; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_420 = 6'h24 == fb_wire_bindex ? _T_2868 : btb_hcount_36; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_421 = 6'h25 == fb_wire_bindex ? _T_2868 : btb_hcount_37; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_422 = 6'h26 == fb_wire_bindex ? _T_2868 : btb_hcount_38; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_423 = 6'h27 == fb_wire_bindex ? _T_2868 : btb_hcount_39; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_424 = 6'h28 == fb_wire_bindex ? _T_2868 : btb_hcount_40; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_425 = 6'h29 == fb_wire_bindex ? _T_2868 : btb_hcount_41; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_426 = 6'h2a == fb_wire_bindex ? _T_2868 : btb_hcount_42; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_427 = 6'h2b == fb_wire_bindex ? _T_2868 : btb_hcount_43; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_428 = 6'h2c == fb_wire_bindex ? _T_2868 : btb_hcount_44; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_429 = 6'h2d == fb_wire_bindex ? _T_2868 : btb_hcount_45; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_430 = 6'h2e == fb_wire_bindex ? _T_2868 : btb_hcount_46; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_431 = 6'h2f == fb_wire_bindex ? _T_2868 : btb_hcount_47; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_432 = 6'h30 == fb_wire_bindex ? _T_2868 : btb_hcount_48; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_433 = 6'h31 == fb_wire_bindex ? _T_2868 : btb_hcount_49; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_434 = 6'h32 == fb_wire_bindex ? _T_2868 : btb_hcount_50; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_435 = 6'h33 == fb_wire_bindex ? _T_2868 : btb_hcount_51; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_436 = 6'h34 == fb_wire_bindex ? _T_2868 : btb_hcount_52; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_437 = 6'h35 == fb_wire_bindex ? _T_2868 : btb_hcount_53; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_438 = 6'h36 == fb_wire_bindex ? _T_2868 : btb_hcount_54; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_439 = 6'h37 == fb_wire_bindex ? _T_2868 : btb_hcount_55; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_440 = 6'h38 == fb_wire_bindex ? _T_2868 : btb_hcount_56; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_441 = 6'h39 == fb_wire_bindex ? _T_2868 : btb_hcount_57; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_442 = 6'h3a == fb_wire_bindex ? _T_2868 : btb_hcount_58; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_443 = 6'h3b == fb_wire_bindex ? _T_2868 : btb_hcount_59; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_444 = 6'h3c == fb_wire_bindex ? _T_2868 : btb_hcount_60; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_445 = 6'h3d == fb_wire_bindex ? _T_2868 : btb_hcount_61; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_446 = 6'h3e == fb_wire_bindex ? _T_2868 : btb_hcount_62; // @[BTB.scala 131:38:@2504.12]
  assign _GEN_447 = 6'h3f == fb_wire_bindex ? _T_2868 : btb_hcount_63; // @[BTB.scala 131:38:@2504.12]
  assign _T_2869 = ~ fb_wire_hcount; // @[BTB.scala 52:42:@2507.12]
  assign _T_2871 = _T_2869 == 2'h0; // @[BTB.scala 52:42:@2508.12]
  assign _T_2876 = _T_2863 & _T_2866; // @[BTB.scala 52:53:@2512.12]
  assign _T_2877 = {_T_2871,_T_2876}; // @[Cat.scala 30:58:@2513.12]
  assign _GEN_448 = 6'h0 == fb_wire_bindex ? _T_2877 : btb_hcount_0; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_449 = 6'h1 == fb_wire_bindex ? _T_2877 : btb_hcount_1; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_450 = 6'h2 == fb_wire_bindex ? _T_2877 : btb_hcount_2; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_451 = 6'h3 == fb_wire_bindex ? _T_2877 : btb_hcount_3; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_452 = 6'h4 == fb_wire_bindex ? _T_2877 : btb_hcount_4; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_453 = 6'h5 == fb_wire_bindex ? _T_2877 : btb_hcount_5; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_454 = 6'h6 == fb_wire_bindex ? _T_2877 : btb_hcount_6; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_455 = 6'h7 == fb_wire_bindex ? _T_2877 : btb_hcount_7; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_456 = 6'h8 == fb_wire_bindex ? _T_2877 : btb_hcount_8; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_457 = 6'h9 == fb_wire_bindex ? _T_2877 : btb_hcount_9; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_458 = 6'ha == fb_wire_bindex ? _T_2877 : btb_hcount_10; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_459 = 6'hb == fb_wire_bindex ? _T_2877 : btb_hcount_11; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_460 = 6'hc == fb_wire_bindex ? _T_2877 : btb_hcount_12; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_461 = 6'hd == fb_wire_bindex ? _T_2877 : btb_hcount_13; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_462 = 6'he == fb_wire_bindex ? _T_2877 : btb_hcount_14; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_463 = 6'hf == fb_wire_bindex ? _T_2877 : btb_hcount_15; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_464 = 6'h10 == fb_wire_bindex ? _T_2877 : btb_hcount_16; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_465 = 6'h11 == fb_wire_bindex ? _T_2877 : btb_hcount_17; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_466 = 6'h12 == fb_wire_bindex ? _T_2877 : btb_hcount_18; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_467 = 6'h13 == fb_wire_bindex ? _T_2877 : btb_hcount_19; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_468 = 6'h14 == fb_wire_bindex ? _T_2877 : btb_hcount_20; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_469 = 6'h15 == fb_wire_bindex ? _T_2877 : btb_hcount_21; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_470 = 6'h16 == fb_wire_bindex ? _T_2877 : btb_hcount_22; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_471 = 6'h17 == fb_wire_bindex ? _T_2877 : btb_hcount_23; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_472 = 6'h18 == fb_wire_bindex ? _T_2877 : btb_hcount_24; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_473 = 6'h19 == fb_wire_bindex ? _T_2877 : btb_hcount_25; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_474 = 6'h1a == fb_wire_bindex ? _T_2877 : btb_hcount_26; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_475 = 6'h1b == fb_wire_bindex ? _T_2877 : btb_hcount_27; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_476 = 6'h1c == fb_wire_bindex ? _T_2877 : btb_hcount_28; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_477 = 6'h1d == fb_wire_bindex ? _T_2877 : btb_hcount_29; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_478 = 6'h1e == fb_wire_bindex ? _T_2877 : btb_hcount_30; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_479 = 6'h1f == fb_wire_bindex ? _T_2877 : btb_hcount_31; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_480 = 6'h20 == fb_wire_bindex ? _T_2877 : btb_hcount_32; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_481 = 6'h21 == fb_wire_bindex ? _T_2877 : btb_hcount_33; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_482 = 6'h22 == fb_wire_bindex ? _T_2877 : btb_hcount_34; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_483 = 6'h23 == fb_wire_bindex ? _T_2877 : btb_hcount_35; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_484 = 6'h24 == fb_wire_bindex ? _T_2877 : btb_hcount_36; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_485 = 6'h25 == fb_wire_bindex ? _T_2877 : btb_hcount_37; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_486 = 6'h26 == fb_wire_bindex ? _T_2877 : btb_hcount_38; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_487 = 6'h27 == fb_wire_bindex ? _T_2877 : btb_hcount_39; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_488 = 6'h28 == fb_wire_bindex ? _T_2877 : btb_hcount_40; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_489 = 6'h29 == fb_wire_bindex ? _T_2877 : btb_hcount_41; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_490 = 6'h2a == fb_wire_bindex ? _T_2877 : btb_hcount_42; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_491 = 6'h2b == fb_wire_bindex ? _T_2877 : btb_hcount_43; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_492 = 6'h2c == fb_wire_bindex ? _T_2877 : btb_hcount_44; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_493 = 6'h2d == fb_wire_bindex ? _T_2877 : btb_hcount_45; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_494 = 6'h2e == fb_wire_bindex ? _T_2877 : btb_hcount_46; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_495 = 6'h2f == fb_wire_bindex ? _T_2877 : btb_hcount_47; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_496 = 6'h30 == fb_wire_bindex ? _T_2877 : btb_hcount_48; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_497 = 6'h31 == fb_wire_bindex ? _T_2877 : btb_hcount_49; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_498 = 6'h32 == fb_wire_bindex ? _T_2877 : btb_hcount_50; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_499 = 6'h33 == fb_wire_bindex ? _T_2877 : btb_hcount_51; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_500 = 6'h34 == fb_wire_bindex ? _T_2877 : btb_hcount_52; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_501 = 6'h35 == fb_wire_bindex ? _T_2877 : btb_hcount_53; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_502 = 6'h36 == fb_wire_bindex ? _T_2877 : btb_hcount_54; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_503 = 6'h37 == fb_wire_bindex ? _T_2877 : btb_hcount_55; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_504 = 6'h38 == fb_wire_bindex ? _T_2877 : btb_hcount_56; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_505 = 6'h39 == fb_wire_bindex ? _T_2877 : btb_hcount_57; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_506 = 6'h3a == fb_wire_bindex ? _T_2877 : btb_hcount_58; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_507 = 6'h3b == fb_wire_bindex ? _T_2877 : btb_hcount_59; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_508 = 6'h3c == fb_wire_bindex ? _T_2877 : btb_hcount_60; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_509 = 6'h3d == fb_wire_bindex ? _T_2877 : btb_hcount_61; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_510 = 6'h3e == fb_wire_bindex ? _T_2877 : btb_hcount_62; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_511 = 6'h3f == fb_wire_bindex ? _T_2877 : btb_hcount_63; // @[BTB.scala 133:38:@2514.12]
  assign _GEN_512 = fb_reg_redirect ? _GEN_384 : _GEN_448; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_513 = fb_reg_redirect ? _GEN_385 : _GEN_449; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_514 = fb_reg_redirect ? _GEN_386 : _GEN_450; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_515 = fb_reg_redirect ? _GEN_387 : _GEN_451; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_516 = fb_reg_redirect ? _GEN_388 : _GEN_452; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_517 = fb_reg_redirect ? _GEN_389 : _GEN_453; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_518 = fb_reg_redirect ? _GEN_390 : _GEN_454; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_519 = fb_reg_redirect ? _GEN_391 : _GEN_455; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_520 = fb_reg_redirect ? _GEN_392 : _GEN_456; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_521 = fb_reg_redirect ? _GEN_393 : _GEN_457; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_522 = fb_reg_redirect ? _GEN_394 : _GEN_458; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_523 = fb_reg_redirect ? _GEN_395 : _GEN_459; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_524 = fb_reg_redirect ? _GEN_396 : _GEN_460; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_525 = fb_reg_redirect ? _GEN_397 : _GEN_461; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_526 = fb_reg_redirect ? _GEN_398 : _GEN_462; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_527 = fb_reg_redirect ? _GEN_399 : _GEN_463; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_528 = fb_reg_redirect ? _GEN_400 : _GEN_464; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_529 = fb_reg_redirect ? _GEN_401 : _GEN_465; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_530 = fb_reg_redirect ? _GEN_402 : _GEN_466; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_531 = fb_reg_redirect ? _GEN_403 : _GEN_467; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_532 = fb_reg_redirect ? _GEN_404 : _GEN_468; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_533 = fb_reg_redirect ? _GEN_405 : _GEN_469; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_534 = fb_reg_redirect ? _GEN_406 : _GEN_470; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_535 = fb_reg_redirect ? _GEN_407 : _GEN_471; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_536 = fb_reg_redirect ? _GEN_408 : _GEN_472; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_537 = fb_reg_redirect ? _GEN_409 : _GEN_473; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_538 = fb_reg_redirect ? _GEN_410 : _GEN_474; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_539 = fb_reg_redirect ? _GEN_411 : _GEN_475; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_540 = fb_reg_redirect ? _GEN_412 : _GEN_476; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_541 = fb_reg_redirect ? _GEN_413 : _GEN_477; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_542 = fb_reg_redirect ? _GEN_414 : _GEN_478; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_543 = fb_reg_redirect ? _GEN_415 : _GEN_479; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_544 = fb_reg_redirect ? _GEN_416 : _GEN_480; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_545 = fb_reg_redirect ? _GEN_417 : _GEN_481; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_546 = fb_reg_redirect ? _GEN_418 : _GEN_482; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_547 = fb_reg_redirect ? _GEN_419 : _GEN_483; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_548 = fb_reg_redirect ? _GEN_420 : _GEN_484; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_549 = fb_reg_redirect ? _GEN_421 : _GEN_485; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_550 = fb_reg_redirect ? _GEN_422 : _GEN_486; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_551 = fb_reg_redirect ? _GEN_423 : _GEN_487; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_552 = fb_reg_redirect ? _GEN_424 : _GEN_488; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_553 = fb_reg_redirect ? _GEN_425 : _GEN_489; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_554 = fb_reg_redirect ? _GEN_426 : _GEN_490; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_555 = fb_reg_redirect ? _GEN_427 : _GEN_491; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_556 = fb_reg_redirect ? _GEN_428 : _GEN_492; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_557 = fb_reg_redirect ? _GEN_429 : _GEN_493; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_558 = fb_reg_redirect ? _GEN_430 : _GEN_494; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_559 = fb_reg_redirect ? _GEN_431 : _GEN_495; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_560 = fb_reg_redirect ? _GEN_432 : _GEN_496; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_561 = fb_reg_redirect ? _GEN_433 : _GEN_497; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_562 = fb_reg_redirect ? _GEN_434 : _GEN_498; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_563 = fb_reg_redirect ? _GEN_435 : _GEN_499; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_564 = fb_reg_redirect ? _GEN_436 : _GEN_500; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_565 = fb_reg_redirect ? _GEN_437 : _GEN_501; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_566 = fb_reg_redirect ? _GEN_438 : _GEN_502; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_567 = fb_reg_redirect ? _GEN_439 : _GEN_503; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_568 = fb_reg_redirect ? _GEN_440 : _GEN_504; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_569 = fb_reg_redirect ? _GEN_441 : _GEN_505; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_570 = fb_reg_redirect ? _GEN_442 : _GEN_506; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_571 = fb_reg_redirect ? _GEN_443 : _GEN_507; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_572 = fb_reg_redirect ? _GEN_444 : _GEN_508; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_573 = fb_reg_redirect ? _GEN_445 : _GEN_509; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_574 = fb_reg_redirect ? _GEN_446 : _GEN_510; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_575 = fb_reg_redirect ? _GEN_447 : _GEN_511; // @[BTB.scala 130:32:@2497.10]
  assign _GEN_576 = 6'h0 == fb_wire_bindex ? 2'h2 : btb_hcount_0; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_577 = 6'h1 == fb_wire_bindex ? 2'h2 : btb_hcount_1; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_578 = 6'h2 == fb_wire_bindex ? 2'h2 : btb_hcount_2; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_579 = 6'h3 == fb_wire_bindex ? 2'h2 : btb_hcount_3; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_580 = 6'h4 == fb_wire_bindex ? 2'h2 : btb_hcount_4; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_581 = 6'h5 == fb_wire_bindex ? 2'h2 : btb_hcount_5; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_582 = 6'h6 == fb_wire_bindex ? 2'h2 : btb_hcount_6; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_583 = 6'h7 == fb_wire_bindex ? 2'h2 : btb_hcount_7; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_584 = 6'h8 == fb_wire_bindex ? 2'h2 : btb_hcount_8; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_585 = 6'h9 == fb_wire_bindex ? 2'h2 : btb_hcount_9; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_586 = 6'ha == fb_wire_bindex ? 2'h2 : btb_hcount_10; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_587 = 6'hb == fb_wire_bindex ? 2'h2 : btb_hcount_11; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_588 = 6'hc == fb_wire_bindex ? 2'h2 : btb_hcount_12; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_589 = 6'hd == fb_wire_bindex ? 2'h2 : btb_hcount_13; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_590 = 6'he == fb_wire_bindex ? 2'h2 : btb_hcount_14; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_591 = 6'hf == fb_wire_bindex ? 2'h2 : btb_hcount_15; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_592 = 6'h10 == fb_wire_bindex ? 2'h2 : btb_hcount_16; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_593 = 6'h11 == fb_wire_bindex ? 2'h2 : btb_hcount_17; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_594 = 6'h12 == fb_wire_bindex ? 2'h2 : btb_hcount_18; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_595 = 6'h13 == fb_wire_bindex ? 2'h2 : btb_hcount_19; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_596 = 6'h14 == fb_wire_bindex ? 2'h2 : btb_hcount_20; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_597 = 6'h15 == fb_wire_bindex ? 2'h2 : btb_hcount_21; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_598 = 6'h16 == fb_wire_bindex ? 2'h2 : btb_hcount_22; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_599 = 6'h17 == fb_wire_bindex ? 2'h2 : btb_hcount_23; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_600 = 6'h18 == fb_wire_bindex ? 2'h2 : btb_hcount_24; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_601 = 6'h19 == fb_wire_bindex ? 2'h2 : btb_hcount_25; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_602 = 6'h1a == fb_wire_bindex ? 2'h2 : btb_hcount_26; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_603 = 6'h1b == fb_wire_bindex ? 2'h2 : btb_hcount_27; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_604 = 6'h1c == fb_wire_bindex ? 2'h2 : btb_hcount_28; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_605 = 6'h1d == fb_wire_bindex ? 2'h2 : btb_hcount_29; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_606 = 6'h1e == fb_wire_bindex ? 2'h2 : btb_hcount_30; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_607 = 6'h1f == fb_wire_bindex ? 2'h2 : btb_hcount_31; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_608 = 6'h20 == fb_wire_bindex ? 2'h2 : btb_hcount_32; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_609 = 6'h21 == fb_wire_bindex ? 2'h2 : btb_hcount_33; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_610 = 6'h22 == fb_wire_bindex ? 2'h2 : btb_hcount_34; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_611 = 6'h23 == fb_wire_bindex ? 2'h2 : btb_hcount_35; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_612 = 6'h24 == fb_wire_bindex ? 2'h2 : btb_hcount_36; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_613 = 6'h25 == fb_wire_bindex ? 2'h2 : btb_hcount_37; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_614 = 6'h26 == fb_wire_bindex ? 2'h2 : btb_hcount_38; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_615 = 6'h27 == fb_wire_bindex ? 2'h2 : btb_hcount_39; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_616 = 6'h28 == fb_wire_bindex ? 2'h2 : btb_hcount_40; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_617 = 6'h29 == fb_wire_bindex ? 2'h2 : btb_hcount_41; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_618 = 6'h2a == fb_wire_bindex ? 2'h2 : btb_hcount_42; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_619 = 6'h2b == fb_wire_bindex ? 2'h2 : btb_hcount_43; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_620 = 6'h2c == fb_wire_bindex ? 2'h2 : btb_hcount_44; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_621 = 6'h2d == fb_wire_bindex ? 2'h2 : btb_hcount_45; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_622 = 6'h2e == fb_wire_bindex ? 2'h2 : btb_hcount_46; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_623 = 6'h2f == fb_wire_bindex ? 2'h2 : btb_hcount_47; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_624 = 6'h30 == fb_wire_bindex ? 2'h2 : btb_hcount_48; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_625 = 6'h31 == fb_wire_bindex ? 2'h2 : btb_hcount_49; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_626 = 6'h32 == fb_wire_bindex ? 2'h2 : btb_hcount_50; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_627 = 6'h33 == fb_wire_bindex ? 2'h2 : btb_hcount_51; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_628 = 6'h34 == fb_wire_bindex ? 2'h2 : btb_hcount_52; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_629 = 6'h35 == fb_wire_bindex ? 2'h2 : btb_hcount_53; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_630 = 6'h36 == fb_wire_bindex ? 2'h2 : btb_hcount_54; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_631 = 6'h37 == fb_wire_bindex ? 2'h2 : btb_hcount_55; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_632 = 6'h38 == fb_wire_bindex ? 2'h2 : btb_hcount_56; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_633 = 6'h39 == fb_wire_bindex ? 2'h2 : btb_hcount_57; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_634 = 6'h3a == fb_wire_bindex ? 2'h2 : btb_hcount_58; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_635 = 6'h3b == fb_wire_bindex ? 2'h2 : btb_hcount_59; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_636 = 6'h3c == fb_wire_bindex ? 2'h2 : btb_hcount_60; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_637 = 6'h3d == fb_wire_bindex ? 2'h2 : btb_hcount_61; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_638 = 6'h3e == fb_wire_bindex ? 2'h2 : btb_hcount_62; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_639 = 6'h3f == fb_wire_bindex ? 2'h2 : btb_hcount_63; // @[BTB.scala 136:36:@2519.12]
  assign _GEN_640 = fb_reg_redirect ? _GEN_576 : btb_hcount_0; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_641 = fb_reg_redirect ? _GEN_577 : btb_hcount_1; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_642 = fb_reg_redirect ? _GEN_578 : btb_hcount_2; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_643 = fb_reg_redirect ? _GEN_579 : btb_hcount_3; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_644 = fb_reg_redirect ? _GEN_580 : btb_hcount_4; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_645 = fb_reg_redirect ? _GEN_581 : btb_hcount_5; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_646 = fb_reg_redirect ? _GEN_582 : btb_hcount_6; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_647 = fb_reg_redirect ? _GEN_583 : btb_hcount_7; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_648 = fb_reg_redirect ? _GEN_584 : btb_hcount_8; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_649 = fb_reg_redirect ? _GEN_585 : btb_hcount_9; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_650 = fb_reg_redirect ? _GEN_586 : btb_hcount_10; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_651 = fb_reg_redirect ? _GEN_587 : btb_hcount_11; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_652 = fb_reg_redirect ? _GEN_588 : btb_hcount_12; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_653 = fb_reg_redirect ? _GEN_589 : btb_hcount_13; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_654 = fb_reg_redirect ? _GEN_590 : btb_hcount_14; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_655 = fb_reg_redirect ? _GEN_591 : btb_hcount_15; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_656 = fb_reg_redirect ? _GEN_592 : btb_hcount_16; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_657 = fb_reg_redirect ? _GEN_593 : btb_hcount_17; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_658 = fb_reg_redirect ? _GEN_594 : btb_hcount_18; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_659 = fb_reg_redirect ? _GEN_595 : btb_hcount_19; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_660 = fb_reg_redirect ? _GEN_596 : btb_hcount_20; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_661 = fb_reg_redirect ? _GEN_597 : btb_hcount_21; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_662 = fb_reg_redirect ? _GEN_598 : btb_hcount_22; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_663 = fb_reg_redirect ? _GEN_599 : btb_hcount_23; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_664 = fb_reg_redirect ? _GEN_600 : btb_hcount_24; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_665 = fb_reg_redirect ? _GEN_601 : btb_hcount_25; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_666 = fb_reg_redirect ? _GEN_602 : btb_hcount_26; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_667 = fb_reg_redirect ? _GEN_603 : btb_hcount_27; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_668 = fb_reg_redirect ? _GEN_604 : btb_hcount_28; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_669 = fb_reg_redirect ? _GEN_605 : btb_hcount_29; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_670 = fb_reg_redirect ? _GEN_606 : btb_hcount_30; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_671 = fb_reg_redirect ? _GEN_607 : btb_hcount_31; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_672 = fb_reg_redirect ? _GEN_608 : btb_hcount_32; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_673 = fb_reg_redirect ? _GEN_609 : btb_hcount_33; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_674 = fb_reg_redirect ? _GEN_610 : btb_hcount_34; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_675 = fb_reg_redirect ? _GEN_611 : btb_hcount_35; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_676 = fb_reg_redirect ? _GEN_612 : btb_hcount_36; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_677 = fb_reg_redirect ? _GEN_613 : btb_hcount_37; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_678 = fb_reg_redirect ? _GEN_614 : btb_hcount_38; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_679 = fb_reg_redirect ? _GEN_615 : btb_hcount_39; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_680 = fb_reg_redirect ? _GEN_616 : btb_hcount_40; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_681 = fb_reg_redirect ? _GEN_617 : btb_hcount_41; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_682 = fb_reg_redirect ? _GEN_618 : btb_hcount_42; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_683 = fb_reg_redirect ? _GEN_619 : btb_hcount_43; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_684 = fb_reg_redirect ? _GEN_620 : btb_hcount_44; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_685 = fb_reg_redirect ? _GEN_621 : btb_hcount_45; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_686 = fb_reg_redirect ? _GEN_622 : btb_hcount_46; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_687 = fb_reg_redirect ? _GEN_623 : btb_hcount_47; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_688 = fb_reg_redirect ? _GEN_624 : btb_hcount_48; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_689 = fb_reg_redirect ? _GEN_625 : btb_hcount_49; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_690 = fb_reg_redirect ? _GEN_626 : btb_hcount_50; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_691 = fb_reg_redirect ? _GEN_627 : btb_hcount_51; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_692 = fb_reg_redirect ? _GEN_628 : btb_hcount_52; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_693 = fb_reg_redirect ? _GEN_629 : btb_hcount_53; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_694 = fb_reg_redirect ? _GEN_630 : btb_hcount_54; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_695 = fb_reg_redirect ? _GEN_631 : btb_hcount_55; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_696 = fb_reg_redirect ? _GEN_632 : btb_hcount_56; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_697 = fb_reg_redirect ? _GEN_633 : btb_hcount_57; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_698 = fb_reg_redirect ? _GEN_634 : btb_hcount_58; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_699 = fb_reg_redirect ? _GEN_635 : btb_hcount_59; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_700 = fb_reg_redirect ? _GEN_636 : btb_hcount_60; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_701 = fb_reg_redirect ? _GEN_637 : btb_hcount_61; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_702 = fb_reg_redirect ? _GEN_638 : btb_hcount_62; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_703 = fb_reg_redirect ? _GEN_639 : btb_hcount_63; // @[BTB.scala 135:35:@2518.10]
  assign _GEN_704 = _T_2106 ? _GEN_512 : _GEN_640; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_705 = _T_2106 ? _GEN_513 : _GEN_641; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_706 = _T_2106 ? _GEN_514 : _GEN_642; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_707 = _T_2106 ? _GEN_515 : _GEN_643; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_708 = _T_2106 ? _GEN_516 : _GEN_644; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_709 = _T_2106 ? _GEN_517 : _GEN_645; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_710 = _T_2106 ? _GEN_518 : _GEN_646; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_711 = _T_2106 ? _GEN_519 : _GEN_647; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_712 = _T_2106 ? _GEN_520 : _GEN_648; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_713 = _T_2106 ? _GEN_521 : _GEN_649; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_714 = _T_2106 ? _GEN_522 : _GEN_650; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_715 = _T_2106 ? _GEN_523 : _GEN_651; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_716 = _T_2106 ? _GEN_524 : _GEN_652; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_717 = _T_2106 ? _GEN_525 : _GEN_653; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_718 = _T_2106 ? _GEN_526 : _GEN_654; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_719 = _T_2106 ? _GEN_527 : _GEN_655; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_720 = _T_2106 ? _GEN_528 : _GEN_656; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_721 = _T_2106 ? _GEN_529 : _GEN_657; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_722 = _T_2106 ? _GEN_530 : _GEN_658; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_723 = _T_2106 ? _GEN_531 : _GEN_659; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_724 = _T_2106 ? _GEN_532 : _GEN_660; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_725 = _T_2106 ? _GEN_533 : _GEN_661; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_726 = _T_2106 ? _GEN_534 : _GEN_662; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_727 = _T_2106 ? _GEN_535 : _GEN_663; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_728 = _T_2106 ? _GEN_536 : _GEN_664; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_729 = _T_2106 ? _GEN_537 : _GEN_665; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_730 = _T_2106 ? _GEN_538 : _GEN_666; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_731 = _T_2106 ? _GEN_539 : _GEN_667; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_732 = _T_2106 ? _GEN_540 : _GEN_668; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_733 = _T_2106 ? _GEN_541 : _GEN_669; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_734 = _T_2106 ? _GEN_542 : _GEN_670; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_735 = _T_2106 ? _GEN_543 : _GEN_671; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_736 = _T_2106 ? _GEN_544 : _GEN_672; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_737 = _T_2106 ? _GEN_545 : _GEN_673; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_738 = _T_2106 ? _GEN_546 : _GEN_674; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_739 = _T_2106 ? _GEN_547 : _GEN_675; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_740 = _T_2106 ? _GEN_548 : _GEN_676; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_741 = _T_2106 ? _GEN_549 : _GEN_677; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_742 = _T_2106 ? _GEN_550 : _GEN_678; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_743 = _T_2106 ? _GEN_551 : _GEN_679; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_744 = _T_2106 ? _GEN_552 : _GEN_680; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_745 = _T_2106 ? _GEN_553 : _GEN_681; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_746 = _T_2106 ? _GEN_554 : _GEN_682; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_747 = _T_2106 ? _GEN_555 : _GEN_683; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_748 = _T_2106 ? _GEN_556 : _GEN_684; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_749 = _T_2106 ? _GEN_557 : _GEN_685; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_750 = _T_2106 ? _GEN_558 : _GEN_686; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_751 = _T_2106 ? _GEN_559 : _GEN_687; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_752 = _T_2106 ? _GEN_560 : _GEN_688; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_753 = _T_2106 ? _GEN_561 : _GEN_689; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_754 = _T_2106 ? _GEN_562 : _GEN_690; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_755 = _T_2106 ? _GEN_563 : _GEN_691; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_756 = _T_2106 ? _GEN_564 : _GEN_692; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_757 = _T_2106 ? _GEN_565 : _GEN_693; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_758 = _T_2106 ? _GEN_566 : _GEN_694; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_759 = _T_2106 ? _GEN_567 : _GEN_695; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_760 = _T_2106 ? _GEN_568 : _GEN_696; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_761 = _T_2106 ? _GEN_569 : _GEN_697; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_762 = _T_2106 ? _GEN_570 : _GEN_698; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_763 = _T_2106 ? _GEN_571 : _GEN_699; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_764 = _T_2106 ? _GEN_572 : _GEN_700; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_765 = _T_2106 ? _GEN_573 : _GEN_701; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_766 = _T_2106 ? _GEN_574 : _GEN_702; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_767 = _T_2106 ? _GEN_575 : _GEN_703; // @[BTB.scala 129:28:@2496.8]
  assign _GEN_768 = _T_2858 ? _GEN_704 : btb_hcount_0; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_769 = _T_2858 ? _GEN_705 : btb_hcount_1; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_770 = _T_2858 ? _GEN_706 : btb_hcount_2; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_771 = _T_2858 ? _GEN_707 : btb_hcount_3; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_772 = _T_2858 ? _GEN_708 : btb_hcount_4; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_773 = _T_2858 ? _GEN_709 : btb_hcount_5; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_774 = _T_2858 ? _GEN_710 : btb_hcount_6; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_775 = _T_2858 ? _GEN_711 : btb_hcount_7; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_776 = _T_2858 ? _GEN_712 : btb_hcount_8; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_777 = _T_2858 ? _GEN_713 : btb_hcount_9; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_778 = _T_2858 ? _GEN_714 : btb_hcount_10; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_779 = _T_2858 ? _GEN_715 : btb_hcount_11; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_780 = _T_2858 ? _GEN_716 : btb_hcount_12; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_781 = _T_2858 ? _GEN_717 : btb_hcount_13; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_782 = _T_2858 ? _GEN_718 : btb_hcount_14; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_783 = _T_2858 ? _GEN_719 : btb_hcount_15; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_784 = _T_2858 ? _GEN_720 : btb_hcount_16; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_785 = _T_2858 ? _GEN_721 : btb_hcount_17; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_786 = _T_2858 ? _GEN_722 : btb_hcount_18; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_787 = _T_2858 ? _GEN_723 : btb_hcount_19; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_788 = _T_2858 ? _GEN_724 : btb_hcount_20; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_789 = _T_2858 ? _GEN_725 : btb_hcount_21; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_790 = _T_2858 ? _GEN_726 : btb_hcount_22; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_791 = _T_2858 ? _GEN_727 : btb_hcount_23; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_792 = _T_2858 ? _GEN_728 : btb_hcount_24; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_793 = _T_2858 ? _GEN_729 : btb_hcount_25; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_794 = _T_2858 ? _GEN_730 : btb_hcount_26; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_795 = _T_2858 ? _GEN_731 : btb_hcount_27; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_796 = _T_2858 ? _GEN_732 : btb_hcount_28; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_797 = _T_2858 ? _GEN_733 : btb_hcount_29; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_798 = _T_2858 ? _GEN_734 : btb_hcount_30; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_799 = _T_2858 ? _GEN_735 : btb_hcount_31; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_800 = _T_2858 ? _GEN_736 : btb_hcount_32; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_801 = _T_2858 ? _GEN_737 : btb_hcount_33; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_802 = _T_2858 ? _GEN_738 : btb_hcount_34; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_803 = _T_2858 ? _GEN_739 : btb_hcount_35; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_804 = _T_2858 ? _GEN_740 : btb_hcount_36; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_805 = _T_2858 ? _GEN_741 : btb_hcount_37; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_806 = _T_2858 ? _GEN_742 : btb_hcount_38; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_807 = _T_2858 ? _GEN_743 : btb_hcount_39; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_808 = _T_2858 ? _GEN_744 : btb_hcount_40; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_809 = _T_2858 ? _GEN_745 : btb_hcount_41; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_810 = _T_2858 ? _GEN_746 : btb_hcount_42; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_811 = _T_2858 ? _GEN_747 : btb_hcount_43; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_812 = _T_2858 ? _GEN_748 : btb_hcount_44; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_813 = _T_2858 ? _GEN_749 : btb_hcount_45; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_814 = _T_2858 ? _GEN_750 : btb_hcount_46; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_815 = _T_2858 ? _GEN_751 : btb_hcount_47; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_816 = _T_2858 ? _GEN_752 : btb_hcount_48; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_817 = _T_2858 ? _GEN_753 : btb_hcount_49; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_818 = _T_2858 ? _GEN_754 : btb_hcount_50; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_819 = _T_2858 ? _GEN_755 : btb_hcount_51; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_820 = _T_2858 ? _GEN_756 : btb_hcount_52; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_821 = _T_2858 ? _GEN_757 : btb_hcount_53; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_822 = _T_2858 ? _GEN_758 : btb_hcount_54; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_823 = _T_2858 ? _GEN_759 : btb_hcount_55; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_824 = _T_2858 ? _GEN_760 : btb_hcount_56; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_825 = _T_2858 ? _GEN_761 : btb_hcount_57; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_826 = _T_2858 ? _GEN_762 : btb_hcount_58; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_827 = _T_2858 ? _GEN_763 : btb_hcount_59; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_828 = _T_2858 ? _GEN_764 : btb_hcount_60; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_829 = _T_2858 ? _GEN_765 : btb_hcount_61; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_830 = _T_2858 ? _GEN_766 : btb_hcount_62; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_831 = _T_2858 ? _GEN_767 : btb_hcount_63; // @[BTB.scala 128:46:@2494.6]
  assign _GEN_832 = fb_reg_valid ? _GEN_192 : btb_pc_0; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_833 = fb_reg_valid ? _GEN_193 : btb_pc_1; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_834 = fb_reg_valid ? _GEN_194 : btb_pc_2; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_835 = fb_reg_valid ? _GEN_195 : btb_pc_3; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_836 = fb_reg_valid ? _GEN_196 : btb_pc_4; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_837 = fb_reg_valid ? _GEN_197 : btb_pc_5; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_838 = fb_reg_valid ? _GEN_198 : btb_pc_6; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_839 = fb_reg_valid ? _GEN_199 : btb_pc_7; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_840 = fb_reg_valid ? _GEN_200 : btb_pc_8; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_841 = fb_reg_valid ? _GEN_201 : btb_pc_9; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_842 = fb_reg_valid ? _GEN_202 : btb_pc_10; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_843 = fb_reg_valid ? _GEN_203 : btb_pc_11; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_844 = fb_reg_valid ? _GEN_204 : btb_pc_12; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_845 = fb_reg_valid ? _GEN_205 : btb_pc_13; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_846 = fb_reg_valid ? _GEN_206 : btb_pc_14; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_847 = fb_reg_valid ? _GEN_207 : btb_pc_15; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_848 = fb_reg_valid ? _GEN_208 : btb_pc_16; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_849 = fb_reg_valid ? _GEN_209 : btb_pc_17; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_850 = fb_reg_valid ? _GEN_210 : btb_pc_18; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_851 = fb_reg_valid ? _GEN_211 : btb_pc_19; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_852 = fb_reg_valid ? _GEN_212 : btb_pc_20; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_853 = fb_reg_valid ? _GEN_213 : btb_pc_21; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_854 = fb_reg_valid ? _GEN_214 : btb_pc_22; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_855 = fb_reg_valid ? _GEN_215 : btb_pc_23; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_856 = fb_reg_valid ? _GEN_216 : btb_pc_24; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_857 = fb_reg_valid ? _GEN_217 : btb_pc_25; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_858 = fb_reg_valid ? _GEN_218 : btb_pc_26; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_859 = fb_reg_valid ? _GEN_219 : btb_pc_27; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_860 = fb_reg_valid ? _GEN_220 : btb_pc_28; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_861 = fb_reg_valid ? _GEN_221 : btb_pc_29; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_862 = fb_reg_valid ? _GEN_222 : btb_pc_30; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_863 = fb_reg_valid ? _GEN_223 : btb_pc_31; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_864 = fb_reg_valid ? _GEN_224 : btb_pc_32; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_865 = fb_reg_valid ? _GEN_225 : btb_pc_33; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_866 = fb_reg_valid ? _GEN_226 : btb_pc_34; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_867 = fb_reg_valid ? _GEN_227 : btb_pc_35; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_868 = fb_reg_valid ? _GEN_228 : btb_pc_36; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_869 = fb_reg_valid ? _GEN_229 : btb_pc_37; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_870 = fb_reg_valid ? _GEN_230 : btb_pc_38; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_871 = fb_reg_valid ? _GEN_231 : btb_pc_39; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_872 = fb_reg_valid ? _GEN_232 : btb_pc_40; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_873 = fb_reg_valid ? _GEN_233 : btb_pc_41; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_874 = fb_reg_valid ? _GEN_234 : btb_pc_42; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_875 = fb_reg_valid ? _GEN_235 : btb_pc_43; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_876 = fb_reg_valid ? _GEN_236 : btb_pc_44; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_877 = fb_reg_valid ? _GEN_237 : btb_pc_45; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_878 = fb_reg_valid ? _GEN_238 : btb_pc_46; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_879 = fb_reg_valid ? _GEN_239 : btb_pc_47; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_880 = fb_reg_valid ? _GEN_240 : btb_pc_48; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_881 = fb_reg_valid ? _GEN_241 : btb_pc_49; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_882 = fb_reg_valid ? _GEN_242 : btb_pc_50; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_883 = fb_reg_valid ? _GEN_243 : btb_pc_51; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_884 = fb_reg_valid ? _GEN_244 : btb_pc_52; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_885 = fb_reg_valid ? _GEN_245 : btb_pc_53; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_886 = fb_reg_valid ? _GEN_246 : btb_pc_54; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_887 = fb_reg_valid ? _GEN_247 : btb_pc_55; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_888 = fb_reg_valid ? _GEN_248 : btb_pc_56; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_889 = fb_reg_valid ? _GEN_249 : btb_pc_57; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_890 = fb_reg_valid ? _GEN_250 : btb_pc_58; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_891 = fb_reg_valid ? _GEN_251 : btb_pc_59; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_892 = fb_reg_valid ? _GEN_252 : btb_pc_60; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_893 = fb_reg_valid ? _GEN_253 : btb_pc_61; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_894 = fb_reg_valid ? _GEN_254 : btb_pc_62; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_895 = fb_reg_valid ? _GEN_255 : btb_pc_63; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_896 = fb_reg_valid ? _GEN_256 : btb_target_0; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_897 = fb_reg_valid ? _GEN_257 : btb_target_1; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_898 = fb_reg_valid ? _GEN_258 : btb_target_2; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_899 = fb_reg_valid ? _GEN_259 : btb_target_3; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_900 = fb_reg_valid ? _GEN_260 : btb_target_4; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_901 = fb_reg_valid ? _GEN_261 : btb_target_5; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_902 = fb_reg_valid ? _GEN_262 : btb_target_6; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_903 = fb_reg_valid ? _GEN_263 : btb_target_7; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_904 = fb_reg_valid ? _GEN_264 : btb_target_8; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_905 = fb_reg_valid ? _GEN_265 : btb_target_9; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_906 = fb_reg_valid ? _GEN_266 : btb_target_10; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_907 = fb_reg_valid ? _GEN_267 : btb_target_11; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_908 = fb_reg_valid ? _GEN_268 : btb_target_12; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_909 = fb_reg_valid ? _GEN_269 : btb_target_13; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_910 = fb_reg_valid ? _GEN_270 : btb_target_14; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_911 = fb_reg_valid ? _GEN_271 : btb_target_15; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_912 = fb_reg_valid ? _GEN_272 : btb_target_16; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_913 = fb_reg_valid ? _GEN_273 : btb_target_17; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_914 = fb_reg_valid ? _GEN_274 : btb_target_18; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_915 = fb_reg_valid ? _GEN_275 : btb_target_19; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_916 = fb_reg_valid ? _GEN_276 : btb_target_20; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_917 = fb_reg_valid ? _GEN_277 : btb_target_21; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_918 = fb_reg_valid ? _GEN_278 : btb_target_22; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_919 = fb_reg_valid ? _GEN_279 : btb_target_23; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_920 = fb_reg_valid ? _GEN_280 : btb_target_24; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_921 = fb_reg_valid ? _GEN_281 : btb_target_25; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_922 = fb_reg_valid ? _GEN_282 : btb_target_26; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_923 = fb_reg_valid ? _GEN_283 : btb_target_27; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_924 = fb_reg_valid ? _GEN_284 : btb_target_28; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_925 = fb_reg_valid ? _GEN_285 : btb_target_29; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_926 = fb_reg_valid ? _GEN_286 : btb_target_30; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_927 = fb_reg_valid ? _GEN_287 : btb_target_31; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_928 = fb_reg_valid ? _GEN_288 : btb_target_32; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_929 = fb_reg_valid ? _GEN_289 : btb_target_33; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_930 = fb_reg_valid ? _GEN_290 : btb_target_34; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_931 = fb_reg_valid ? _GEN_291 : btb_target_35; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_932 = fb_reg_valid ? _GEN_292 : btb_target_36; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_933 = fb_reg_valid ? _GEN_293 : btb_target_37; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_934 = fb_reg_valid ? _GEN_294 : btb_target_38; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_935 = fb_reg_valid ? _GEN_295 : btb_target_39; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_936 = fb_reg_valid ? _GEN_296 : btb_target_40; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_937 = fb_reg_valid ? _GEN_297 : btb_target_41; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_938 = fb_reg_valid ? _GEN_298 : btb_target_42; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_939 = fb_reg_valid ? _GEN_299 : btb_target_43; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_940 = fb_reg_valid ? _GEN_300 : btb_target_44; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_941 = fb_reg_valid ? _GEN_301 : btb_target_45; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_942 = fb_reg_valid ? _GEN_302 : btb_target_46; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_943 = fb_reg_valid ? _GEN_303 : btb_target_47; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_944 = fb_reg_valid ? _GEN_304 : btb_target_48; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_945 = fb_reg_valid ? _GEN_305 : btb_target_49; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_946 = fb_reg_valid ? _GEN_306 : btb_target_50; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_947 = fb_reg_valid ? _GEN_307 : btb_target_51; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_948 = fb_reg_valid ? _GEN_308 : btb_target_52; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_949 = fb_reg_valid ? _GEN_309 : btb_target_53; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_950 = fb_reg_valid ? _GEN_310 : btb_target_54; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_951 = fb_reg_valid ? _GEN_311 : btb_target_55; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_952 = fb_reg_valid ? _GEN_312 : btb_target_56; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_953 = fb_reg_valid ? _GEN_313 : btb_target_57; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_954 = fb_reg_valid ? _GEN_314 : btb_target_58; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_955 = fb_reg_valid ? _GEN_315 : btb_target_59; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_956 = fb_reg_valid ? _GEN_316 : btb_target_60; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_957 = fb_reg_valid ? _GEN_317 : btb_target_61; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_958 = fb_reg_valid ? _GEN_318 : btb_target_62; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_959 = fb_reg_valid ? _GEN_319 : btb_target_63; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_960 = fb_reg_valid ? _GEN_320 : btb_btype_0; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_961 = fb_reg_valid ? _GEN_321 : btb_btype_1; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_962 = fb_reg_valid ? _GEN_322 : btb_btype_2; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_963 = fb_reg_valid ? _GEN_323 : btb_btype_3; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_964 = fb_reg_valid ? _GEN_324 : btb_btype_4; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_965 = fb_reg_valid ? _GEN_325 : btb_btype_5; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_966 = fb_reg_valid ? _GEN_326 : btb_btype_6; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_967 = fb_reg_valid ? _GEN_327 : btb_btype_7; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_968 = fb_reg_valid ? _GEN_328 : btb_btype_8; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_969 = fb_reg_valid ? _GEN_329 : btb_btype_9; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_970 = fb_reg_valid ? _GEN_330 : btb_btype_10; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_971 = fb_reg_valid ? _GEN_331 : btb_btype_11; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_972 = fb_reg_valid ? _GEN_332 : btb_btype_12; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_973 = fb_reg_valid ? _GEN_333 : btb_btype_13; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_974 = fb_reg_valid ? _GEN_334 : btb_btype_14; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_975 = fb_reg_valid ? _GEN_335 : btb_btype_15; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_976 = fb_reg_valid ? _GEN_336 : btb_btype_16; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_977 = fb_reg_valid ? _GEN_337 : btb_btype_17; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_978 = fb_reg_valid ? _GEN_338 : btb_btype_18; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_979 = fb_reg_valid ? _GEN_339 : btb_btype_19; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_980 = fb_reg_valid ? _GEN_340 : btb_btype_20; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_981 = fb_reg_valid ? _GEN_341 : btb_btype_21; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_982 = fb_reg_valid ? _GEN_342 : btb_btype_22; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_983 = fb_reg_valid ? _GEN_343 : btb_btype_23; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_984 = fb_reg_valid ? _GEN_344 : btb_btype_24; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_985 = fb_reg_valid ? _GEN_345 : btb_btype_25; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_986 = fb_reg_valid ? _GEN_346 : btb_btype_26; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_987 = fb_reg_valid ? _GEN_347 : btb_btype_27; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_988 = fb_reg_valid ? _GEN_348 : btb_btype_28; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_989 = fb_reg_valid ? _GEN_349 : btb_btype_29; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_990 = fb_reg_valid ? _GEN_350 : btb_btype_30; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_991 = fb_reg_valid ? _GEN_351 : btb_btype_31; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_992 = fb_reg_valid ? _GEN_352 : btb_btype_32; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_993 = fb_reg_valid ? _GEN_353 : btb_btype_33; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_994 = fb_reg_valid ? _GEN_354 : btb_btype_34; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_995 = fb_reg_valid ? _GEN_355 : btb_btype_35; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_996 = fb_reg_valid ? _GEN_356 : btb_btype_36; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_997 = fb_reg_valid ? _GEN_357 : btb_btype_37; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_998 = fb_reg_valid ? _GEN_358 : btb_btype_38; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_999 = fb_reg_valid ? _GEN_359 : btb_btype_39; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1000 = fb_reg_valid ? _GEN_360 : btb_btype_40; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1001 = fb_reg_valid ? _GEN_361 : btb_btype_41; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1002 = fb_reg_valid ? _GEN_362 : btb_btype_42; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1003 = fb_reg_valid ? _GEN_363 : btb_btype_43; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1004 = fb_reg_valid ? _GEN_364 : btb_btype_44; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1005 = fb_reg_valid ? _GEN_365 : btb_btype_45; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1006 = fb_reg_valid ? _GEN_366 : btb_btype_46; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1007 = fb_reg_valid ? _GEN_367 : btb_btype_47; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1008 = fb_reg_valid ? _GEN_368 : btb_btype_48; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1009 = fb_reg_valid ? _GEN_369 : btb_btype_49; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1010 = fb_reg_valid ? _GEN_370 : btb_btype_50; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1011 = fb_reg_valid ? _GEN_371 : btb_btype_51; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1012 = fb_reg_valid ? _GEN_372 : btb_btype_52; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1013 = fb_reg_valid ? _GEN_373 : btb_btype_53; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1014 = fb_reg_valid ? _GEN_374 : btb_btype_54; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1015 = fb_reg_valid ? _GEN_375 : btb_btype_55; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1016 = fb_reg_valid ? _GEN_376 : btb_btype_56; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1017 = fb_reg_valid ? _GEN_377 : btb_btype_57; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1018 = fb_reg_valid ? _GEN_378 : btb_btype_58; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1019 = fb_reg_valid ? _GEN_379 : btb_btype_59; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1020 = fb_reg_valid ? _GEN_380 : btb_btype_60; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1021 = fb_reg_valid ? _GEN_381 : btb_btype_61; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1022 = fb_reg_valid ? _GEN_382 : btb_btype_62; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1023 = fb_reg_valid ? _GEN_383 : btb_btype_63; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1024 = fb_reg_valid ? _GEN_768 : btb_hcount_0; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1025 = fb_reg_valid ? _GEN_769 : btb_hcount_1; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1026 = fb_reg_valid ? _GEN_770 : btb_hcount_2; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1027 = fb_reg_valid ? _GEN_771 : btb_hcount_3; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1028 = fb_reg_valid ? _GEN_772 : btb_hcount_4; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1029 = fb_reg_valid ? _GEN_773 : btb_hcount_5; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1030 = fb_reg_valid ? _GEN_774 : btb_hcount_6; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1031 = fb_reg_valid ? _GEN_775 : btb_hcount_7; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1032 = fb_reg_valid ? _GEN_776 : btb_hcount_8; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1033 = fb_reg_valid ? _GEN_777 : btb_hcount_9; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1034 = fb_reg_valid ? _GEN_778 : btb_hcount_10; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1035 = fb_reg_valid ? _GEN_779 : btb_hcount_11; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1036 = fb_reg_valid ? _GEN_780 : btb_hcount_12; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1037 = fb_reg_valid ? _GEN_781 : btb_hcount_13; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1038 = fb_reg_valid ? _GEN_782 : btb_hcount_14; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1039 = fb_reg_valid ? _GEN_783 : btb_hcount_15; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1040 = fb_reg_valid ? _GEN_784 : btb_hcount_16; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1041 = fb_reg_valid ? _GEN_785 : btb_hcount_17; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1042 = fb_reg_valid ? _GEN_786 : btb_hcount_18; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1043 = fb_reg_valid ? _GEN_787 : btb_hcount_19; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1044 = fb_reg_valid ? _GEN_788 : btb_hcount_20; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1045 = fb_reg_valid ? _GEN_789 : btb_hcount_21; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1046 = fb_reg_valid ? _GEN_790 : btb_hcount_22; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1047 = fb_reg_valid ? _GEN_791 : btb_hcount_23; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1048 = fb_reg_valid ? _GEN_792 : btb_hcount_24; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1049 = fb_reg_valid ? _GEN_793 : btb_hcount_25; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1050 = fb_reg_valid ? _GEN_794 : btb_hcount_26; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1051 = fb_reg_valid ? _GEN_795 : btb_hcount_27; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1052 = fb_reg_valid ? _GEN_796 : btb_hcount_28; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1053 = fb_reg_valid ? _GEN_797 : btb_hcount_29; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1054 = fb_reg_valid ? _GEN_798 : btb_hcount_30; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1055 = fb_reg_valid ? _GEN_799 : btb_hcount_31; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1056 = fb_reg_valid ? _GEN_800 : btb_hcount_32; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1057 = fb_reg_valid ? _GEN_801 : btb_hcount_33; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1058 = fb_reg_valid ? _GEN_802 : btb_hcount_34; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1059 = fb_reg_valid ? _GEN_803 : btb_hcount_35; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1060 = fb_reg_valid ? _GEN_804 : btb_hcount_36; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1061 = fb_reg_valid ? _GEN_805 : btb_hcount_37; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1062 = fb_reg_valid ? _GEN_806 : btb_hcount_38; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1063 = fb_reg_valid ? _GEN_807 : btb_hcount_39; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1064 = fb_reg_valid ? _GEN_808 : btb_hcount_40; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1065 = fb_reg_valid ? _GEN_809 : btb_hcount_41; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1066 = fb_reg_valid ? _GEN_810 : btb_hcount_42; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1067 = fb_reg_valid ? _GEN_811 : btb_hcount_43; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1068 = fb_reg_valid ? _GEN_812 : btb_hcount_44; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1069 = fb_reg_valid ? _GEN_813 : btb_hcount_45; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1070 = fb_reg_valid ? _GEN_814 : btb_hcount_46; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1071 = fb_reg_valid ? _GEN_815 : btb_hcount_47; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1072 = fb_reg_valid ? _GEN_816 : btb_hcount_48; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1073 = fb_reg_valid ? _GEN_817 : btb_hcount_49; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1074 = fb_reg_valid ? _GEN_818 : btb_hcount_50; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1075 = fb_reg_valid ? _GEN_819 : btb_hcount_51; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1076 = fb_reg_valid ? _GEN_820 : btb_hcount_52; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1077 = fb_reg_valid ? _GEN_821 : btb_hcount_53; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1078 = fb_reg_valid ? _GEN_822 : btb_hcount_54; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1079 = fb_reg_valid ? _GEN_823 : btb_hcount_55; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1080 = fb_reg_valid ? _GEN_824 : btb_hcount_56; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1081 = fb_reg_valid ? _GEN_825 : btb_hcount_57; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1082 = fb_reg_valid ? _GEN_826 : btb_hcount_58; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1083 = fb_reg_valid ? _GEN_827 : btb_hcount_59; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1084 = fb_reg_valid ? _GEN_828 : btb_hcount_60; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1085 = fb_reg_valid ? _GEN_829 : btb_hcount_61; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1086 = fb_reg_valid ? _GEN_830 : btb_hcount_62; // @[BTB.scala 122:23:@2487.4]
  assign _GEN_1087 = fb_reg_valid ? _GEN_831 : btb_hcount_63; // @[BTB.scala 122:23:@2487.4]
  assign io_pred_pc = _T_1362 ? io_ras_peek : _T_1374; // @[BTB.scala 76:14:@1342.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  btb_pc_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  btb_pc_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  btb_pc_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  btb_pc_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  btb_pc_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  btb_pc_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  btb_pc_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  btb_pc_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  btb_pc_8 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  btb_pc_9 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  btb_pc_10 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  btb_pc_11 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  btb_pc_12 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  btb_pc_13 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  btb_pc_14 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  btb_pc_15 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  btb_pc_16 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  btb_pc_17 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  btb_pc_18 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  btb_pc_19 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  btb_pc_20 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  btb_pc_21 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  btb_pc_22 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  btb_pc_23 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  btb_pc_24 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  btb_pc_25 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  btb_pc_26 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  btb_pc_27 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  btb_pc_28 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  btb_pc_29 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  btb_pc_30 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  btb_pc_31 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  btb_pc_32 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  btb_pc_33 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  btb_pc_34 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  btb_pc_35 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  btb_pc_36 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  btb_pc_37 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  btb_pc_38 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  btb_pc_39 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  btb_pc_40 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  btb_pc_41 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{`RANDOM}};
  btb_pc_42 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{`RANDOM}};
  btb_pc_43 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{`RANDOM}};
  btb_pc_44 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{`RANDOM}};
  btb_pc_45 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{`RANDOM}};
  btb_pc_46 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{`RANDOM}};
  btb_pc_47 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  btb_pc_48 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{`RANDOM}};
  btb_pc_49 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{`RANDOM}};
  btb_pc_50 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{`RANDOM}};
  btb_pc_51 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{`RANDOM}};
  btb_pc_52 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{`RANDOM}};
  btb_pc_53 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{`RANDOM}};
  btb_pc_54 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{`RANDOM}};
  btb_pc_55 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{`RANDOM}};
  btb_pc_56 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{`RANDOM}};
  btb_pc_57 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{`RANDOM}};
  btb_pc_58 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{`RANDOM}};
  btb_pc_59 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{`RANDOM}};
  btb_pc_60 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{`RANDOM}};
  btb_pc_61 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{`RANDOM}};
  btb_pc_62 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{`RANDOM}};
  btb_pc_63 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{`RANDOM}};
  btb_target_0 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{`RANDOM}};
  btb_target_1 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{`RANDOM}};
  btb_target_2 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{`RANDOM}};
  btb_target_3 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{`RANDOM}};
  btb_target_4 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{`RANDOM}};
  btb_target_5 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{`RANDOM}};
  btb_target_6 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{`RANDOM}};
  btb_target_7 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{`RANDOM}};
  btb_target_8 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{`RANDOM}};
  btb_target_9 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{`RANDOM}};
  btb_target_10 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{`RANDOM}};
  btb_target_11 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{`RANDOM}};
  btb_target_12 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{`RANDOM}};
  btb_target_13 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{`RANDOM}};
  btb_target_14 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{`RANDOM}};
  btb_target_15 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{`RANDOM}};
  btb_target_16 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{`RANDOM}};
  btb_target_17 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{`RANDOM}};
  btb_target_18 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{`RANDOM}};
  btb_target_19 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{`RANDOM}};
  btb_target_20 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{`RANDOM}};
  btb_target_21 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{`RANDOM}};
  btb_target_22 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{`RANDOM}};
  btb_target_23 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{`RANDOM}};
  btb_target_24 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{`RANDOM}};
  btb_target_25 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{`RANDOM}};
  btb_target_26 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{`RANDOM}};
  btb_target_27 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{`RANDOM}};
  btb_target_28 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{`RANDOM}};
  btb_target_29 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{`RANDOM}};
  btb_target_30 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{`RANDOM}};
  btb_target_31 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{`RANDOM}};
  btb_target_32 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{`RANDOM}};
  btb_target_33 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{`RANDOM}};
  btb_target_34 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{`RANDOM}};
  btb_target_35 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{`RANDOM}};
  btb_target_36 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{`RANDOM}};
  btb_target_37 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{`RANDOM}};
  btb_target_38 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{`RANDOM}};
  btb_target_39 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{`RANDOM}};
  btb_target_40 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{`RANDOM}};
  btb_target_41 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{`RANDOM}};
  btb_target_42 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{`RANDOM}};
  btb_target_43 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{`RANDOM}};
  btb_target_44 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{`RANDOM}};
  btb_target_45 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{`RANDOM}};
  btb_target_46 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{`RANDOM}};
  btb_target_47 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{`RANDOM}};
  btb_target_48 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{`RANDOM}};
  btb_target_49 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{`RANDOM}};
  btb_target_50 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{`RANDOM}};
  btb_target_51 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{`RANDOM}};
  btb_target_52 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{`RANDOM}};
  btb_target_53 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{`RANDOM}};
  btb_target_54 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{`RANDOM}};
  btb_target_55 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{`RANDOM}};
  btb_target_56 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{`RANDOM}};
  btb_target_57 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{`RANDOM}};
  btb_target_58 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{`RANDOM}};
  btb_target_59 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{`RANDOM}};
  btb_target_60 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{`RANDOM}};
  btb_target_61 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{`RANDOM}};
  btb_target_62 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{`RANDOM}};
  btb_target_63 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{`RANDOM}};
  btb_hcount_0 = _RAND_128[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{`RANDOM}};
  btb_hcount_1 = _RAND_129[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{`RANDOM}};
  btb_hcount_2 = _RAND_130[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{`RANDOM}};
  btb_hcount_3 = _RAND_131[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{`RANDOM}};
  btb_hcount_4 = _RAND_132[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{`RANDOM}};
  btb_hcount_5 = _RAND_133[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{`RANDOM}};
  btb_hcount_6 = _RAND_134[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{`RANDOM}};
  btb_hcount_7 = _RAND_135[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{`RANDOM}};
  btb_hcount_8 = _RAND_136[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{`RANDOM}};
  btb_hcount_9 = _RAND_137[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{`RANDOM}};
  btb_hcount_10 = _RAND_138[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{`RANDOM}};
  btb_hcount_11 = _RAND_139[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{`RANDOM}};
  btb_hcount_12 = _RAND_140[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{`RANDOM}};
  btb_hcount_13 = _RAND_141[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{`RANDOM}};
  btb_hcount_14 = _RAND_142[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{`RANDOM}};
  btb_hcount_15 = _RAND_143[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{`RANDOM}};
  btb_hcount_16 = _RAND_144[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{`RANDOM}};
  btb_hcount_17 = _RAND_145[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{`RANDOM}};
  btb_hcount_18 = _RAND_146[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{`RANDOM}};
  btb_hcount_19 = _RAND_147[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{`RANDOM}};
  btb_hcount_20 = _RAND_148[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{`RANDOM}};
  btb_hcount_21 = _RAND_149[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{`RANDOM}};
  btb_hcount_22 = _RAND_150[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{`RANDOM}};
  btb_hcount_23 = _RAND_151[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{`RANDOM}};
  btb_hcount_24 = _RAND_152[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{`RANDOM}};
  btb_hcount_25 = _RAND_153[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{`RANDOM}};
  btb_hcount_26 = _RAND_154[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{`RANDOM}};
  btb_hcount_27 = _RAND_155[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{`RANDOM}};
  btb_hcount_28 = _RAND_156[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{`RANDOM}};
  btb_hcount_29 = _RAND_157[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{`RANDOM}};
  btb_hcount_30 = _RAND_158[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{`RANDOM}};
  btb_hcount_31 = _RAND_159[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{`RANDOM}};
  btb_hcount_32 = _RAND_160[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{`RANDOM}};
  btb_hcount_33 = _RAND_161[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{`RANDOM}};
  btb_hcount_34 = _RAND_162[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{`RANDOM}};
  btb_hcount_35 = _RAND_163[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{`RANDOM}};
  btb_hcount_36 = _RAND_164[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{`RANDOM}};
  btb_hcount_37 = _RAND_165[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{`RANDOM}};
  btb_hcount_38 = _RAND_166[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{`RANDOM}};
  btb_hcount_39 = _RAND_167[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{`RANDOM}};
  btb_hcount_40 = _RAND_168[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{`RANDOM}};
  btb_hcount_41 = _RAND_169[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{`RANDOM}};
  btb_hcount_42 = _RAND_170[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{`RANDOM}};
  btb_hcount_43 = _RAND_171[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{`RANDOM}};
  btb_hcount_44 = _RAND_172[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{`RANDOM}};
  btb_hcount_45 = _RAND_173[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{`RANDOM}};
  btb_hcount_46 = _RAND_174[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{`RANDOM}};
  btb_hcount_47 = _RAND_175[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{`RANDOM}};
  btb_hcount_48 = _RAND_176[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{`RANDOM}};
  btb_hcount_49 = _RAND_177[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{`RANDOM}};
  btb_hcount_50 = _RAND_178[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{`RANDOM}};
  btb_hcount_51 = _RAND_179[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{`RANDOM}};
  btb_hcount_52 = _RAND_180[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{`RANDOM}};
  btb_hcount_53 = _RAND_181[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{`RANDOM}};
  btb_hcount_54 = _RAND_182[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{`RANDOM}};
  btb_hcount_55 = _RAND_183[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{`RANDOM}};
  btb_hcount_56 = _RAND_184[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{`RANDOM}};
  btb_hcount_57 = _RAND_185[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{`RANDOM}};
  btb_hcount_58 = _RAND_186[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{`RANDOM}};
  btb_hcount_59 = _RAND_187[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{`RANDOM}};
  btb_hcount_60 = _RAND_188[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{`RANDOM}};
  btb_hcount_61 = _RAND_189[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{`RANDOM}};
  btb_hcount_62 = _RAND_190[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{`RANDOM}};
  btb_hcount_63 = _RAND_191[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{`RANDOM}};
  btb_btype_0 = _RAND_192[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{`RANDOM}};
  btb_btype_1 = _RAND_193[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{`RANDOM}};
  btb_btype_2 = _RAND_194[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{`RANDOM}};
  btb_btype_3 = _RAND_195[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{`RANDOM}};
  btb_btype_4 = _RAND_196[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{`RANDOM}};
  btb_btype_5 = _RAND_197[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{`RANDOM}};
  btb_btype_6 = _RAND_198[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{`RANDOM}};
  btb_btype_7 = _RAND_199[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{`RANDOM}};
  btb_btype_8 = _RAND_200[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{`RANDOM}};
  btb_btype_9 = _RAND_201[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{`RANDOM}};
  btb_btype_10 = _RAND_202[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{`RANDOM}};
  btb_btype_11 = _RAND_203[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{`RANDOM}};
  btb_btype_12 = _RAND_204[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{`RANDOM}};
  btb_btype_13 = _RAND_205[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{`RANDOM}};
  btb_btype_14 = _RAND_206[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{`RANDOM}};
  btb_btype_15 = _RAND_207[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{`RANDOM}};
  btb_btype_16 = _RAND_208[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{`RANDOM}};
  btb_btype_17 = _RAND_209[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{`RANDOM}};
  btb_btype_18 = _RAND_210[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{`RANDOM}};
  btb_btype_19 = _RAND_211[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{`RANDOM}};
  btb_btype_20 = _RAND_212[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{`RANDOM}};
  btb_btype_21 = _RAND_213[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{`RANDOM}};
  btb_btype_22 = _RAND_214[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{`RANDOM}};
  btb_btype_23 = _RAND_215[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{`RANDOM}};
  btb_btype_24 = _RAND_216[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{`RANDOM}};
  btb_btype_25 = _RAND_217[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{`RANDOM}};
  btb_btype_26 = _RAND_218[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{`RANDOM}};
  btb_btype_27 = _RAND_219[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{`RANDOM}};
  btb_btype_28 = _RAND_220[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{`RANDOM}};
  btb_btype_29 = _RAND_221[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{`RANDOM}};
  btb_btype_30 = _RAND_222[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{`RANDOM}};
  btb_btype_31 = _RAND_223[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{`RANDOM}};
  btb_btype_32 = _RAND_224[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{`RANDOM}};
  btb_btype_33 = _RAND_225[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{`RANDOM}};
  btb_btype_34 = _RAND_226[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{`RANDOM}};
  btb_btype_35 = _RAND_227[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{`RANDOM}};
  btb_btype_36 = _RAND_228[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{`RANDOM}};
  btb_btype_37 = _RAND_229[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{`RANDOM}};
  btb_btype_38 = _RAND_230[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{`RANDOM}};
  btb_btype_39 = _RAND_231[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{`RANDOM}};
  btb_btype_40 = _RAND_232[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_233 = {1{`RANDOM}};
  btb_btype_41 = _RAND_233[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_234 = {1{`RANDOM}};
  btb_btype_42 = _RAND_234[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_235 = {1{`RANDOM}};
  btb_btype_43 = _RAND_235[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_236 = {1{`RANDOM}};
  btb_btype_44 = _RAND_236[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_237 = {1{`RANDOM}};
  btb_btype_45 = _RAND_237[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_238 = {1{`RANDOM}};
  btb_btype_46 = _RAND_238[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_239 = {1{`RANDOM}};
  btb_btype_47 = _RAND_239[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_240 = {1{`RANDOM}};
  btb_btype_48 = _RAND_240[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_241 = {1{`RANDOM}};
  btb_btype_49 = _RAND_241[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_242 = {1{`RANDOM}};
  btb_btype_50 = _RAND_242[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_243 = {1{`RANDOM}};
  btb_btype_51 = _RAND_243[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_244 = {1{`RANDOM}};
  btb_btype_52 = _RAND_244[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_245 = {1{`RANDOM}};
  btb_btype_53 = _RAND_245[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_246 = {1{`RANDOM}};
  btb_btype_54 = _RAND_246[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_247 = {1{`RANDOM}};
  btb_btype_55 = _RAND_247[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_248 = {1{`RANDOM}};
  btb_btype_56 = _RAND_248[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_249 = {1{`RANDOM}};
  btb_btype_57 = _RAND_249[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_250 = {1{`RANDOM}};
  btb_btype_58 = _RAND_250[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_251 = {1{`RANDOM}};
  btb_btype_59 = _RAND_251[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_252 = {1{`RANDOM}};
  btb_btype_60 = _RAND_252[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_253 = {1{`RANDOM}};
  btb_btype_61 = _RAND_253[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_254 = {1{`RANDOM}};
  btb_btype_62 = _RAND_254[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_255 = {1{`RANDOM}};
  btb_btype_63 = _RAND_255[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_256 = {1{`RANDOM}};
  fb_reg_valid = _RAND_256[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_257 = {1{`RANDOM}};
  fb_reg_redirect = _RAND_257[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_258 = {1{`RANDOM}};
  fb_reg_lfsr = _RAND_258[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_259 = {1{`RANDOM}};
  fb_reg_pc = _RAND_259[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_260 = {1{`RANDOM}};
  fb_reg_target = _RAND_260[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_261 = {1{`RANDOM}};
  fb_reg_btype = _RAND_261[1:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      btb_pc_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_pc_0 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_pc_1 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_pc_2 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_pc_3 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_pc_4 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_pc_5 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_pc_6 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_pc_7 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_pc_8 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_pc_9 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_pc_10 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_pc_11 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_pc_12 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_pc_13 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_pc_14 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_pc_15 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_pc_16 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_pc_17 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_pc_18 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_pc_19 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_pc_20 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_pc_21 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_pc_22 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_pc_23 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_pc_24 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_pc_25 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_pc_26 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_pc_27 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_pc_28 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_pc_29 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_pc_30 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_pc_31 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_pc_32 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_pc_33 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_pc_34 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_pc_35 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_pc_36 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_pc_37 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_pc_38 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_pc_39 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_pc_40 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_pc_41 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_pc_42 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_pc_43 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_pc_44 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_pc_45 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_pc_46 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_pc_47 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_pc_48 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_pc_49 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_pc_50 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_pc_51 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_pc_52 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_pc_53 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_pc_54 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_pc_55 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_pc_56 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_pc_57 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_pc_58 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_pc_59 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_pc_60 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_pc_61 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_pc_62 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_pc_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_pc_63 <= fb_reg_pc;
          end
        end
      end
    end
    if (reset) begin
      btb_target_0 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_target_0 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_1 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_target_1 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_2 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_target_2 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_3 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_target_3 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_4 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_target_4 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_5 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_target_5 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_6 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_target_6 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_7 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_target_7 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_8 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_target_8 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_9 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_target_9 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_10 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_target_10 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_11 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_target_11 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_12 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_target_12 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_13 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_target_13 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_14 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_target_14 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_15 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_target_15 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_16 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_target_16 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_17 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_target_17 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_18 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_target_18 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_19 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_target_19 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_20 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_target_20 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_21 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_target_21 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_22 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_target_22 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_23 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_target_23 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_24 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_target_24 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_25 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_target_25 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_26 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_target_26 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_27 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_target_27 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_28 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_target_28 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_29 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_target_29 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_30 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_target_30 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_31 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_target_31 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_32 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_target_32 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_33 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_target_33 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_34 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_target_34 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_35 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_target_35 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_36 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_target_36 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_37 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_target_37 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_38 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_target_38 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_39 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_target_39 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_40 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_target_40 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_41 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_target_41 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_42 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_target_42 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_43 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_target_43 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_44 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_target_44 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_45 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_target_45 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_46 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_target_46 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_47 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_target_47 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_48 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_target_48 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_49 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_target_49 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_50 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_target_50 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_51 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_target_51 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_52 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_target_52 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_53 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_target_53 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_54 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_target_54 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_55 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_target_55 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_56 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_target_56 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_57 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_target_57 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_58 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_target_58 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_59 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_target_59 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_60 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_target_60 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_61 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_target_61 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_62 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_target_62 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_target_63 <= 32'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_target_63 <= fb_reg_target;
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= _T_2868;
              end
            end else begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h0 == fb_wire_bindex) begin
                btb_hcount_0 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= _T_2868;
              end
            end else begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1 == fb_wire_bindex) begin
                btb_hcount_1 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= _T_2868;
              end
            end else begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2 == fb_wire_bindex) begin
                btb_hcount_2 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= _T_2868;
              end
            end else begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3 == fb_wire_bindex) begin
                btb_hcount_3 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= _T_2868;
              end
            end else begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h4 == fb_wire_bindex) begin
                btb_hcount_4 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= _T_2868;
              end
            end else begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h5 == fb_wire_bindex) begin
                btb_hcount_5 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= _T_2868;
              end
            end else begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h6 == fb_wire_bindex) begin
                btb_hcount_6 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= _T_2868;
              end
            end else begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h7 == fb_wire_bindex) begin
                btb_hcount_7 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= _T_2868;
              end
            end else begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h8 == fb_wire_bindex) begin
                btb_hcount_8 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= _T_2868;
              end
            end else begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h9 == fb_wire_bindex) begin
                btb_hcount_9 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= _T_2868;
              end
            end else begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'ha == fb_wire_bindex) begin
                btb_hcount_10 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= _T_2868;
              end
            end else begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hb == fb_wire_bindex) begin
                btb_hcount_11 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= _T_2868;
              end
            end else begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hc == fb_wire_bindex) begin
                btb_hcount_12 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= _T_2868;
              end
            end else begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hd == fb_wire_bindex) begin
                btb_hcount_13 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= _T_2868;
              end
            end else begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'he == fb_wire_bindex) begin
                btb_hcount_14 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= _T_2868;
              end
            end else begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'hf == fb_wire_bindex) begin
                btb_hcount_15 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= _T_2868;
              end
            end else begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h10 == fb_wire_bindex) begin
                btb_hcount_16 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= _T_2868;
              end
            end else begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h11 == fb_wire_bindex) begin
                btb_hcount_17 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= _T_2868;
              end
            end else begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h12 == fb_wire_bindex) begin
                btb_hcount_18 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= _T_2868;
              end
            end else begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h13 == fb_wire_bindex) begin
                btb_hcount_19 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= _T_2868;
              end
            end else begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h14 == fb_wire_bindex) begin
                btb_hcount_20 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= _T_2868;
              end
            end else begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h15 == fb_wire_bindex) begin
                btb_hcount_21 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= _T_2868;
              end
            end else begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h16 == fb_wire_bindex) begin
                btb_hcount_22 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= _T_2868;
              end
            end else begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h17 == fb_wire_bindex) begin
                btb_hcount_23 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= _T_2868;
              end
            end else begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h18 == fb_wire_bindex) begin
                btb_hcount_24 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= _T_2868;
              end
            end else begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h19 == fb_wire_bindex) begin
                btb_hcount_25 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= _T_2868;
              end
            end else begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1a == fb_wire_bindex) begin
                btb_hcount_26 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= _T_2868;
              end
            end else begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1b == fb_wire_bindex) begin
                btb_hcount_27 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= _T_2868;
              end
            end else begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1c == fb_wire_bindex) begin
                btb_hcount_28 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= _T_2868;
              end
            end else begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1d == fb_wire_bindex) begin
                btb_hcount_29 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= _T_2868;
              end
            end else begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1e == fb_wire_bindex) begin
                btb_hcount_30 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= _T_2868;
              end
            end else begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h1f == fb_wire_bindex) begin
                btb_hcount_31 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= _T_2868;
              end
            end else begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h20 == fb_wire_bindex) begin
                btb_hcount_32 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= _T_2868;
              end
            end else begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h21 == fb_wire_bindex) begin
                btb_hcount_33 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= _T_2868;
              end
            end else begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h22 == fb_wire_bindex) begin
                btb_hcount_34 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= _T_2868;
              end
            end else begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h23 == fb_wire_bindex) begin
                btb_hcount_35 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= _T_2868;
              end
            end else begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h24 == fb_wire_bindex) begin
                btb_hcount_36 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= _T_2868;
              end
            end else begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h25 == fb_wire_bindex) begin
                btb_hcount_37 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= _T_2868;
              end
            end else begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h26 == fb_wire_bindex) begin
                btb_hcount_38 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= _T_2868;
              end
            end else begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h27 == fb_wire_bindex) begin
                btb_hcount_39 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= _T_2868;
              end
            end else begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h28 == fb_wire_bindex) begin
                btb_hcount_40 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= _T_2868;
              end
            end else begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h29 == fb_wire_bindex) begin
                btb_hcount_41 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= _T_2868;
              end
            end else begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2a == fb_wire_bindex) begin
                btb_hcount_42 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= _T_2868;
              end
            end else begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2b == fb_wire_bindex) begin
                btb_hcount_43 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= _T_2868;
              end
            end else begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2c == fb_wire_bindex) begin
                btb_hcount_44 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= _T_2868;
              end
            end else begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2d == fb_wire_bindex) begin
                btb_hcount_45 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= _T_2868;
              end
            end else begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2e == fb_wire_bindex) begin
                btb_hcount_46 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= _T_2868;
              end
            end else begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h2f == fb_wire_bindex) begin
                btb_hcount_47 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= _T_2868;
              end
            end else begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h30 == fb_wire_bindex) begin
                btb_hcount_48 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= _T_2868;
              end
            end else begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h31 == fb_wire_bindex) begin
                btb_hcount_49 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= _T_2868;
              end
            end else begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h32 == fb_wire_bindex) begin
                btb_hcount_50 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= _T_2868;
              end
            end else begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h33 == fb_wire_bindex) begin
                btb_hcount_51 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= _T_2868;
              end
            end else begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h34 == fb_wire_bindex) begin
                btb_hcount_52 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= _T_2868;
              end
            end else begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h35 == fb_wire_bindex) begin
                btb_hcount_53 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= _T_2868;
              end
            end else begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h36 == fb_wire_bindex) begin
                btb_hcount_54 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= _T_2868;
              end
            end else begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h37 == fb_wire_bindex) begin
                btb_hcount_55 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= _T_2868;
              end
            end else begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h38 == fb_wire_bindex) begin
                btb_hcount_56 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= _T_2868;
              end
            end else begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h39 == fb_wire_bindex) begin
                btb_hcount_57 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= _T_2868;
              end
            end else begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3a == fb_wire_bindex) begin
                btb_hcount_58 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= _T_2868;
              end
            end else begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3b == fb_wire_bindex) begin
                btb_hcount_59 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= _T_2868;
              end
            end else begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3c == fb_wire_bindex) begin
                btb_hcount_60 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= _T_2868;
              end
            end else begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3d == fb_wire_bindex) begin
                btb_hcount_61 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= _T_2868;
              end
            end else begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3e == fb_wire_bindex) begin
                btb_hcount_62 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_hcount_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (_T_2858) begin
          if (_T_2106) begin
            if (fb_reg_redirect) begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= _T_2868;
              end
            end else begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= _T_2877;
              end
            end
          end else begin
            if (fb_reg_redirect) begin
              if (6'h3f == fb_wire_bindex) begin
                btb_hcount_63 <= 2'h2;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      btb_btype_0 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h0 == fb_wire_bindex) begin
            btb_btype_0 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_1 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1 == fb_wire_bindex) begin
            btb_btype_1 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_2 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2 == fb_wire_bindex) begin
            btb_btype_2 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_3 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3 == fb_wire_bindex) begin
            btb_btype_3 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_4 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h4 == fb_wire_bindex) begin
            btb_btype_4 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_5 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h5 == fb_wire_bindex) begin
            btb_btype_5 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_6 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h6 == fb_wire_bindex) begin
            btb_btype_6 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_7 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h7 == fb_wire_bindex) begin
            btb_btype_7 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_8 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h8 == fb_wire_bindex) begin
            btb_btype_8 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_9 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h9 == fb_wire_bindex) begin
            btb_btype_9 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_10 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'ha == fb_wire_bindex) begin
            btb_btype_10 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_11 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hb == fb_wire_bindex) begin
            btb_btype_11 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_12 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hc == fb_wire_bindex) begin
            btb_btype_12 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_13 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hd == fb_wire_bindex) begin
            btb_btype_13 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_14 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'he == fb_wire_bindex) begin
            btb_btype_14 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_15 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'hf == fb_wire_bindex) begin
            btb_btype_15 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_16 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h10 == fb_wire_bindex) begin
            btb_btype_16 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_17 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h11 == fb_wire_bindex) begin
            btb_btype_17 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_18 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h12 == fb_wire_bindex) begin
            btb_btype_18 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_19 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h13 == fb_wire_bindex) begin
            btb_btype_19 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_20 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h14 == fb_wire_bindex) begin
            btb_btype_20 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_21 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h15 == fb_wire_bindex) begin
            btb_btype_21 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_22 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h16 == fb_wire_bindex) begin
            btb_btype_22 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_23 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h17 == fb_wire_bindex) begin
            btb_btype_23 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_24 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h18 == fb_wire_bindex) begin
            btb_btype_24 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_25 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h19 == fb_wire_bindex) begin
            btb_btype_25 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_26 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1a == fb_wire_bindex) begin
            btb_btype_26 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_27 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1b == fb_wire_bindex) begin
            btb_btype_27 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_28 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1c == fb_wire_bindex) begin
            btb_btype_28 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_29 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1d == fb_wire_bindex) begin
            btb_btype_29 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_30 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1e == fb_wire_bindex) begin
            btb_btype_30 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_31 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h1f == fb_wire_bindex) begin
            btb_btype_31 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_32 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h20 == fb_wire_bindex) begin
            btb_btype_32 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_33 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h21 == fb_wire_bindex) begin
            btb_btype_33 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_34 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h22 == fb_wire_bindex) begin
            btb_btype_34 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_35 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h23 == fb_wire_bindex) begin
            btb_btype_35 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_36 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h24 == fb_wire_bindex) begin
            btb_btype_36 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_37 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h25 == fb_wire_bindex) begin
            btb_btype_37 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_38 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h26 == fb_wire_bindex) begin
            btb_btype_38 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_39 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h27 == fb_wire_bindex) begin
            btb_btype_39 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_40 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h28 == fb_wire_bindex) begin
            btb_btype_40 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_41 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h29 == fb_wire_bindex) begin
            btb_btype_41 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_42 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2a == fb_wire_bindex) begin
            btb_btype_42 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_43 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2b == fb_wire_bindex) begin
            btb_btype_43 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_44 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2c == fb_wire_bindex) begin
            btb_btype_44 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_45 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2d == fb_wire_bindex) begin
            btb_btype_45 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_46 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2e == fb_wire_bindex) begin
            btb_btype_46 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_47 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h2f == fb_wire_bindex) begin
            btb_btype_47 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_48 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h30 == fb_wire_bindex) begin
            btb_btype_48 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_49 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h31 == fb_wire_bindex) begin
            btb_btype_49 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_50 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h32 == fb_wire_bindex) begin
            btb_btype_50 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_51 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h33 == fb_wire_bindex) begin
            btb_btype_51 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_52 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h34 == fb_wire_bindex) begin
            btb_btype_52 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_53 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h35 == fb_wire_bindex) begin
            btb_btype_53 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_54 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h36 == fb_wire_bindex) begin
            btb_btype_54 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_55 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h37 == fb_wire_bindex) begin
            btb_btype_55 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_56 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h38 == fb_wire_bindex) begin
            btb_btype_56 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_57 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h39 == fb_wire_bindex) begin
            btb_btype_57 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_58 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3a == fb_wire_bindex) begin
            btb_btype_58 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_59 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3b == fb_wire_bindex) begin
            btb_btype_59 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_60 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3c == fb_wire_bindex) begin
            btb_btype_60 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_61 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3d == fb_wire_bindex) begin
            btb_btype_61 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_62 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3e == fb_wire_bindex) begin
            btb_btype_62 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      btb_btype_63 <= 2'h0;
    end else begin
      if (fb_reg_valid) begin
        if (fb_reg_redirect) begin
          if (6'h3f == fb_wire_bindex) begin
            btb_btype_63 <= fb_reg_btype;
          end
        end
      end
    end
    if (reset) begin
      fb_reg_valid <= 1'h0;
    end else begin
      fb_reg_valid <= io_feedBack_valid;
    end
    if (reset) begin
      fb_reg_redirect <= 1'h0;
    end else begin
      fb_reg_redirect <= io_feedBack_bits_redirect;
    end
    if (reset) begin
      fb_reg_lfsr <= 6'h1;
    end else begin
      fb_reg_lfsr <= _T_1386;
    end
    if (reset) begin
      fb_reg_pc <= 32'h0;
    end else begin
      fb_reg_pc <= io_fb_pc;
    end
    if (reset) begin
      fb_reg_target <= 32'h0;
    end else begin
      fb_reg_target <= io_feedBack_bits_tgt;
    end
    if (reset) begin
      fb_reg_btype <= 2'h0;
    end else begin
      fb_reg_btype <= io_fb_type;
    end
  end
endmodule
module RAS( // @[:@2524.2]
  input         clock, // @[:@2525.4]
  input         reset, // @[:@2526.4]
  input         io_push_valid, // @[:@2527.4]
  input  [31:0] io_push_bits, // @[:@2527.4]
  input         io_pop, // @[:@2527.4]
  output [31:0] io_peek // @[:@2527.4]
);
  reg [31:0] stack [0:15]; // @[RAS.scala 13:18:@2529.4]
  reg [31:0] _RAND_0;
  wire [31:0] stack__T_23_data; // @[RAS.scala 13:18:@2529.4]
  wire [3:0] stack__T_23_addr; // @[RAS.scala 13:18:@2529.4]
  wire [31:0] stack__T_24_data; // @[RAS.scala 13:18:@2529.4]
  wire [3:0] stack__T_24_addr; // @[RAS.scala 13:18:@2529.4]
  wire  stack__T_24_mask; // @[RAS.scala 13:18:@2529.4]
  wire  stack__T_24_en; // @[RAS.scala 13:18:@2529.4]
  wire [31:0] stack__T_25_data; // @[RAS.scala 13:18:@2529.4]
  wire [3:0] stack__T_25_addr; // @[RAS.scala 13:18:@2529.4]
  wire  stack__T_25_mask; // @[RAS.scala 13:18:@2529.4]
  wire  stack__T_25_en; // @[RAS.scala 13:18:@2529.4]
  reg [3:0] pos; // @[RAS.scala 14:22:@2530.4]
  reg [31:0] _RAND_1;
  reg [3:0] next; // @[RAS.scala 15:22:@2531.4]
  reg [31:0] _RAND_2;
  wire  _GEN_7; // @[RAS.scala 19:18:@2535.6]
  wire  _T_27; // @[RAS.scala 26:26:@2544.4]
  wire  _T_28; // @[RAS.scala 26:23:@2545.4]
  wire [4:0] _T_30; // @[RAS.scala 27:16:@2547.6]
  wire [3:0] _T_31; // @[RAS.scala 27:16:@2548.6]
  wire [4:0] _T_33; // @[RAS.scala 28:18:@2550.6]
  wire [3:0] _T_34; // @[RAS.scala 28:18:@2551.6]
  wire [4:0] _T_36; // @[RAS.scala 31:16:@2556.8]
  wire [4:0] _T_37; // @[RAS.scala 31:16:@2557.8]
  wire [3:0] _T_38; // @[RAS.scala 31:16:@2558.8]
  wire [4:0] _T_40; // @[RAS.scala 32:18:@2560.8]
  wire [4:0] _T_41; // @[RAS.scala 32:18:@2561.8]
  wire [3:0] _T_42; // @[RAS.scala 32:18:@2562.8]
  wire [3:0] _GEN_20; // @[RAS.scala 29:22:@2555.6]
  wire [3:0] _GEN_21; // @[RAS.scala 29:22:@2555.6]
  wire [3:0] _GEN_22; // @[RAS.scala 26:35:@2546.4]
  wire [3:0] _GEN_23; // @[RAS.scala 26:35:@2546.4]
  assign stack__T_23_addr = pos;
  assign stack__T_23_data = stack[stack__T_23_addr]; // @[RAS.scala 13:18:@2529.4]
  assign stack__T_24_data = io_push_bits;
  assign stack__T_24_addr = pos;
  assign stack__T_24_mask = 1'h1;
  assign stack__T_24_en = io_push_valid ? io_pop : 1'h0;
  assign stack__T_25_data = io_push_bits;
  assign stack__T_25_addr = next;
  assign stack__T_25_mask = 1'h1;
  assign stack__T_25_en = io_push_valid ? _GEN_7 : 1'h0;
  assign _GEN_7 = io_pop ? 1'h0 : 1'h1; // @[RAS.scala 19:18:@2535.6]
  assign _T_27 = io_pop == 1'h0; // @[RAS.scala 26:26:@2544.4]
  assign _T_28 = io_push_valid & _T_27; // @[RAS.scala 26:23:@2545.4]
  assign _T_30 = pos + 4'h1; // @[RAS.scala 27:16:@2547.6]
  assign _T_31 = pos + 4'h1; // @[RAS.scala 27:16:@2548.6]
  assign _T_33 = next + 4'h1; // @[RAS.scala 28:18:@2550.6]
  assign _T_34 = next + 4'h1; // @[RAS.scala 28:18:@2551.6]
  assign _T_36 = pos - 4'h1; // @[RAS.scala 31:16:@2556.8]
  assign _T_37 = $unsigned(_T_36); // @[RAS.scala 31:16:@2557.8]
  assign _T_38 = _T_37[3:0]; // @[RAS.scala 31:16:@2558.8]
  assign _T_40 = next - 4'h1; // @[RAS.scala 32:18:@2560.8]
  assign _T_41 = $unsigned(_T_40); // @[RAS.scala 32:18:@2561.8]
  assign _T_42 = _T_41[3:0]; // @[RAS.scala 32:18:@2562.8]
  assign _GEN_20 = io_pop ? _T_38 : pos; // @[RAS.scala 29:22:@2555.6]
  assign _GEN_21 = io_pop ? _T_42 : next; // @[RAS.scala 29:22:@2555.6]
  assign _GEN_22 = _T_28 ? _T_31 : _GEN_20; // @[RAS.scala 26:35:@2546.4]
  assign _GEN_23 = _T_28 ? _T_34 : _GEN_21; // @[RAS.scala 26:35:@2546.4]
  assign io_peek = stack__T_23_data; // @[RAS.scala 16:11:@2533.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 16; initvar = initvar+1)
    stack[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  pos = _RAND_1[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  next = _RAND_2[3:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(stack__T_24_en & stack__T_24_mask) begin
      stack[stack__T_24_addr] <= stack__T_24_data; // @[RAS.scala 13:18:@2529.4]
    end
    if(stack__T_25_en & stack__T_25_mask) begin
      stack[stack__T_25_addr] <= stack__T_25_data; // @[RAS.scala 13:18:@2529.4]
    end
    if (reset) begin
      pos <= 4'hf;
    end else begin
      if (_T_28) begin
        pos <= _T_31;
      end else begin
        if (io_pop) begin
          pos <= _T_38;
        end
      end
    end
    if (reset) begin
      next <= 4'h0;
    end else begin
      if (_T_28) begin
        next <= _T_34;
      end else begin
        if (io_pop) begin
          next <= _T_42;
        end
      end
    end
  end
endmodule
module FrontEnd( // @[:@2566.2]
  input         clock, // @[:@2567.4]
  input         reset, // @[:@2568.4]
  input  [31:0] io_cyc, // @[:@2569.4]
  output        io_mem_req_valid, // @[:@2569.4]
  output [31:0] io_mem_req_bits_addr, // @[:@2569.4]
  input         io_mem_resp_valid, // @[:@2569.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@2569.4]
  input         io_back_xcpt_valid, // @[:@2569.4]
  input  [31:0] io_back_xcpt_bits, // @[:@2569.4]
  input         io_back_kill, // @[:@2569.4]
  input         io_back_fence, // @[:@2569.4]
  input         io_back_forward, // @[:@2569.4]
  input         io_back_ras_pop, // @[:@2569.4]
  input         io_back_ras_push_valid, // @[:@2569.4]
  input  [31:0] io_back_ras_push_bits, // @[:@2569.4]
  input  [31:0] io_back_fb_pc, // @[:@2569.4]
  input  [1:0]  io_back_fb_type, // @[:@2569.4]
  input         io_back_feedBack_valid, // @[:@2569.4]
  input         io_back_feedBack_bits_redirect, // @[:@2569.4]
  input  [31:0] io_back_feedBack_bits_tgt, // @[:@2569.4]
  output        io_back_inst_valid, // @[:@2569.4]
  output [31:0] io_back_inst_bits, // @[:@2569.4]
  output [31:0] io_back_pc, // @[:@2569.4]
  output [31:0] io_back_pred // @[:@2569.4]
);
  wire  FetchInst_clock; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_reset; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_mem_req_valid; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_mem_req_bits_addr; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_mem_resp_valid; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_mem_resp_bits_data; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_if_kill; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_if_fence; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_dec_forward; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_dec_kill; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_if_target; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_btb_target; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_if_forward; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_if_pc; // @[FrontEnd.scala 12:22:@2571.4]
  wire  FetchInst_io_dec_inst_valid; // @[FrontEnd.scala 12:22:@2571.4]
  wire [31:0] FetchInst_io_dec_inst_bits; // @[FrontEnd.scala 12:22:@2571.4]
  wire  BTB_clock; // @[FrontEnd.scala 14:22:@2575.4]
  wire  BTB_reset; // @[FrontEnd.scala 14:22:@2575.4]
  wire [31:0] BTB_io_if_pc; // @[FrontEnd.scala 14:22:@2575.4]
  wire [31:0] BTB_io_ras_peek; // @[FrontEnd.scala 14:22:@2575.4]
  wire [31:0] BTB_io_pred_pc; // @[FrontEnd.scala 14:22:@2575.4]
  wire [31:0] BTB_io_fb_pc; // @[FrontEnd.scala 14:22:@2575.4]
  wire [1:0] BTB_io_fb_type; // @[FrontEnd.scala 14:22:@2575.4]
  wire  BTB_io_feedBack_valid; // @[FrontEnd.scala 14:22:@2575.4]
  wire  BTB_io_feedBack_bits_redirect; // @[FrontEnd.scala 14:22:@2575.4]
  wire [31:0] BTB_io_feedBack_bits_tgt; // @[FrontEnd.scala 14:22:@2575.4]
  wire  RAS_clock; // @[FrontEnd.scala 16:22:@2579.4]
  wire  RAS_reset; // @[FrontEnd.scala 16:22:@2579.4]
  wire  RAS_io_push_valid; // @[FrontEnd.scala 16:22:@2579.4]
  wire [31:0] RAS_io_push_bits; // @[FrontEnd.scala 16:22:@2579.4]
  wire  RAS_io_pop; // @[FrontEnd.scala 16:22:@2579.4]
  wire [31:0] RAS_io_peek; // @[FrontEnd.scala 16:22:@2579.4]
  reg [31:0] dec_reg_pc; // @[FrontEnd.scala 35:23:@2608.4]
  reg [31:0] _RAND_0;
  reg [31:0] dec_reg_pred; // @[FrontEnd.scala 36:25:@2609.4]
  reg [31:0] _RAND_1;
  wire  _T_96; // @[FrontEnd.scala 46:9:@2618.4]
  wire  _T_97; // @[FrontEnd.scala 46:26:@2619.4]
  wire  _T_100; // @[FrontEnd.scala 47:11:@2622.6]
  FetchInst FetchInst ( // @[FrontEnd.scala 12:22:@2571.4]
    .clock(FetchInst_clock),
    .reset(FetchInst_reset),
    .io_mem_req_valid(FetchInst_io_mem_req_valid),
    .io_mem_req_bits_addr(FetchInst_io_mem_req_bits_addr),
    .io_mem_resp_valid(FetchInst_io_mem_resp_valid),
    .io_mem_resp_bits_data(FetchInst_io_mem_resp_bits_data),
    .io_if_kill(FetchInst_io_if_kill),
    .io_if_fence(FetchInst_io_if_fence),
    .io_dec_forward(FetchInst_io_dec_forward),
    .io_dec_kill(FetchInst_io_dec_kill),
    .io_if_target(FetchInst_io_if_target),
    .io_btb_target(FetchInst_io_btb_target),
    .io_if_forward(FetchInst_io_if_forward),
    .io_if_pc(FetchInst_io_if_pc),
    .io_dec_inst_valid(FetchInst_io_dec_inst_valid),
    .io_dec_inst_bits(FetchInst_io_dec_inst_bits)
  );
  BTB BTB ( // @[FrontEnd.scala 14:22:@2575.4]
    .clock(BTB_clock),
    .reset(BTB_reset),
    .io_if_pc(BTB_io_if_pc),
    .io_ras_peek(BTB_io_ras_peek),
    .io_pred_pc(BTB_io_pred_pc),
    .io_fb_pc(BTB_io_fb_pc),
    .io_fb_type(BTB_io_fb_type),
    .io_feedBack_valid(BTB_io_feedBack_valid),
    .io_feedBack_bits_redirect(BTB_io_feedBack_bits_redirect),
    .io_feedBack_bits_tgt(BTB_io_feedBack_bits_tgt)
  );
  RAS RAS ( // @[FrontEnd.scala 16:22:@2579.4]
    .clock(RAS_clock),
    .reset(RAS_reset),
    .io_push_valid(RAS_io_push_valid),
    .io_push_bits(RAS_io_push_bits),
    .io_pop(RAS_io_pop),
    .io_peek(RAS_io_peek)
  );
  assign _T_96 = io_back_forward == 1'h0; // @[FrontEnd.scala 46:9:@2618.4]
  assign _T_97 = _T_96 & io_back_inst_valid; // @[FrontEnd.scala 46:26:@2619.4]
  assign _T_100 = reset == 1'h0; // @[FrontEnd.scala 47:11:@2622.6]
  assign io_mem_req_valid = FetchInst_io_mem_req_valid; // @[FrontEnd.scala 18:14:@2588.4]
  assign io_mem_req_bits_addr = FetchInst_io_mem_req_bits_addr; // @[FrontEnd.scala 18:14:@2587.4]
  assign io_back_inst_valid = FetchInst_io_dec_inst_valid; // @[FrontEnd.scala 44:16:@2617.4]
  assign io_back_inst_bits = FetchInst_io_dec_inst_bits; // @[FrontEnd.scala 44:16:@2616.4]
  assign io_back_pc = dec_reg_pc; // @[FrontEnd.scala 42:16:@2614.4]
  assign io_back_pred = dec_reg_pred; // @[FrontEnd.scala 43:16:@2615.4]
  assign FetchInst_clock = clock; // @[:@2572.4]
  assign FetchInst_reset = reset; // @[:@2573.4]
  assign FetchInst_io_mem_resp_valid = io_mem_resp_valid; // @[FrontEnd.scala 18:14:@2583.4]
  assign FetchInst_io_mem_resp_bits_data = io_mem_resp_bits_data; // @[FrontEnd.scala 18:14:@2582.4]
  assign FetchInst_io_if_kill = FetchInst_io_dec_kill; // @[FrontEnd.scala 21:18:@2593.4]
  assign FetchInst_io_if_fence = io_back_fence; // @[FrontEnd.scala 24:19:@2597.4]
  assign FetchInst_io_dec_forward = io_back_forward; // @[FrontEnd.scala 23:22:@2596.4]
  assign FetchInst_io_dec_kill = io_back_kill | io_back_xcpt_valid; // @[FrontEnd.scala 22:19:@2595.4]
  assign FetchInst_io_if_target = io_back_xcpt_valid ? io_back_xcpt_bits : io_back_feedBack_bits_tgt; // @[FrontEnd.scala 20:20:@2592.4]
  assign FetchInst_io_btb_target = BTB_io_pred_pc; // @[FrontEnd.scala 19:21:@2590.4]
  assign BTB_clock = clock; // @[:@2576.4]
  assign BTB_reset = reset; // @[:@2577.4]
  assign BTB_io_if_pc = FetchInst_io_if_pc; // @[FrontEnd.scala 29:16:@2601.4]
  assign BTB_io_ras_peek = RAS_io_peek; // @[FrontEnd.scala 30:16:@2602.4]
  assign BTB_io_fb_pc = io_back_fb_pc; // @[FrontEnd.scala 31:16:@2603.4]
  assign BTB_io_fb_type = io_back_fb_type; // @[FrontEnd.scala 32:16:@2604.4]
  assign BTB_io_feedBack_valid = io_back_feedBack_valid; // @[FrontEnd.scala 33:16:@2607.4]
  assign BTB_io_feedBack_bits_redirect = io_back_feedBack_bits_redirect; // @[FrontEnd.scala 33:16:@2606.4]
  assign BTB_io_feedBack_bits_tgt = io_back_feedBack_bits_tgt; // @[FrontEnd.scala 33:16:@2605.4]
  assign RAS_clock = clock; // @[:@2580.4]
  assign RAS_reset = reset; // @[:@2581.4]
  assign RAS_io_push_valid = io_back_ras_push_valid; // @[FrontEnd.scala 27:12:@2600.4]
  assign RAS_io_push_bits = io_back_ras_push_bits; // @[FrontEnd.scala 27:12:@2599.4]
  assign RAS_io_pop = io_back_ras_pop; // @[FrontEnd.scala 26:12:@2598.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  dec_reg_pc = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  dec_reg_pred = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (FetchInst_io_if_forward) begin
      dec_reg_pc <= FetchInst_io_if_pc;
    end
    if (FetchInst_io_if_forward) begin
      dec_reg_pred <= BTB_io_pred_pc;
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_97 & _T_100) begin
          $fwrite(32'h80000002,"STALL Cyc= %d\n",io_cyc); // @[FrontEnd.scala 47:11:@2624.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module CSRFile( // @[:@2628.2]
  input         clock, // @[:@2629.4]
  input         reset, // @[:@2630.4]
  input  [2:0]  io_rw_cmd, // @[:@2631.4]
  input  [11:0] io_rw_addr, // @[:@2631.4]
  output [31:0] io_rw_rdata, // @[:@2631.4]
  input  [31:0] io_rw_wdata, // @[:@2631.4]
  output        io_eret, // @[:@2631.4]
  output [1:0]  io_status_prv, // @[:@2631.4]
  output [13:0] io_status_unimp5, // @[:@2631.4]
  output        io_status_mprv, // @[:@2631.4]
  output [1:0]  io_status_unimp4, // @[:@2631.4]
  output [1:0]  io_status_mpp, // @[:@2631.4]
  output [2:0]  io_status_unimp3, // @[:@2631.4]
  output        io_status_mpie, // @[:@2631.4]
  output [2:0]  io_status_unimp2, // @[:@2631.4]
  output        io_status_mie, // @[:@2631.4]
  output [2:0]  io_status_unimp1, // @[:@2631.4]
  input         io_xcpt, // @[:@2631.4]
  input  [31:0] io_cause, // @[:@2631.4]
  input  [31:0] io_tval, // @[:@2631.4]
  output [31:0] io_evec, // @[:@2631.4]
  input         io_illegal, // @[:@2631.4]
  input  [1:0]  io_retire, // @[:@2631.4]
  input  [31:0] io_pc, // @[:@2631.4]
  output [31:0] io_time // @[:@2631.4]
);
  reg [1:0] reg_mstatus_prv; // @[CSR.scala 112:28:@2758.4]
  reg [31:0] _RAND_0;
  reg  reg_mstatus_mpie; // @[CSR.scala 112:28:@2758.4]
  reg [31:0] _RAND_1;
  reg  reg_mstatus_mie; // @[CSR.scala 112:28:@2758.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_mepc; // @[CSR.scala 113:21:@2759.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_mcause; // @[CSR.scala 114:23:@2760.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_mtval; // @[CSR.scala 115:22:@2761.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_mscratch; // @[CSR.scala 116:25:@2762.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_medeleg; // @[CSR.scala 118:24:@2764.4]
  reg [31:0] _RAND_7;
  reg  reg_mip_mtip; // @[CSR.scala 120:24:@2782.4]
  reg [31:0] _RAND_8;
  reg  reg_mip_msip; // @[CSR.scala 120:24:@2782.4]
  reg [31:0] _RAND_9;
  reg  reg_mie_mtip; // @[CSR.scala 121:24:@2800.4]
  reg [31:0] _RAND_10;
  reg  reg_mie_msip; // @[CSR.scala 121:24:@2800.4]
  reg [31:0] _RAND_11;
  reg [5:0] _T_240; // @[Util.scala 112:41:@2803.4]
  reg [31:0] _RAND_12;
  wire [6:0] _T_241; // @[Util.scala 113:33:@2804.4]
  reg [57:0] _T_244; // @[Util.scala 117:31:@2806.4]
  reg [63:0] _RAND_13;
  wire  _T_245; // @[Util.scala 118:20:@2807.4]
  wire [58:0] _T_247; // @[Util.scala 118:43:@2809.6]
  wire [57:0] _T_248; // @[Util.scala 118:43:@2810.6]
  wire [57:0] _GEN_0; // @[Util.scala 118:34:@2808.4]
  wire [63:0] _T_249; // @[Cat.scala 30:58:@2813.4]
  reg [5:0] _T_252; // @[Util.scala 112:41:@2814.4]
  reg [31:0] _RAND_14;
  wire [5:0] _GEN_147; // @[Util.scala 113:33:@2815.4]
  wire [6:0] _T_253; // @[Util.scala 113:33:@2815.4]
  reg [57:0] _T_256; // @[Util.scala 117:31:@2817.4]
  reg [63:0] _RAND_15;
  wire  _T_257; // @[Util.scala 118:20:@2818.4]
  wire [58:0] _T_259; // @[Util.scala 118:43:@2820.6]
  wire [57:0] _T_260; // @[Util.scala 118:43:@2821.6]
  wire [57:0] _GEN_1; // @[Util.scala 118:34:@2819.4]
  wire [63:0] _T_261; // @[Cat.scala 30:58:@2824.4]
  reg [39:0] _T_264; // @[Util.scala 112:74:@2826.4]
  reg [63:0] _RAND_16;
  wire [40:0] _T_265; // @[Util.scala 113:33:@2827.4]
  reg [39:0] _T_267; // @[Util.scala 112:74:@2829.4]
  reg [63:0] _RAND_17;
  wire [40:0] _T_268; // @[Util.scala 113:33:@2830.4]
  reg [39:0] _T_270; // @[Util.scala 112:74:@2832.4]
  reg [63:0] _RAND_18;
  wire [40:0] _T_271; // @[Util.scala 113:33:@2833.4]
  reg [39:0] _T_273; // @[Util.scala 112:74:@2835.4]
  reg [63:0] _RAND_19;
  wire [40:0] _T_274; // @[Util.scala 113:33:@2836.4]
  reg [39:0] _T_276; // @[Util.scala 112:74:@2838.4]
  reg [63:0] _RAND_20;
  wire [40:0] _T_277; // @[Util.scala 113:33:@2839.4]
  reg [39:0] _T_279; // @[Util.scala 112:74:@2841.4]
  reg [63:0] _RAND_21;
  wire [40:0] _T_280; // @[Util.scala 113:33:@2842.4]
  reg [39:0] _T_282; // @[Util.scala 112:74:@2844.4]
  reg [63:0] _RAND_22;
  wire [40:0] _T_283; // @[Util.scala 113:33:@2845.4]
  reg [39:0] _T_285; // @[Util.scala 112:74:@2847.4]
  reg [63:0] _RAND_23;
  wire [40:0] _T_286; // @[Util.scala 113:33:@2848.4]
  reg [39:0] _T_288; // @[Util.scala 112:74:@2850.4]
  reg [63:0] _RAND_24;
  wire [40:0] _T_289; // @[Util.scala 113:33:@2851.4]
  reg [39:0] _T_291; // @[Util.scala 112:74:@2853.4]
  reg [63:0] _RAND_25;
  wire [40:0] _T_292; // @[Util.scala 113:33:@2854.4]
  reg [39:0] _T_294; // @[Util.scala 112:74:@2856.4]
  reg [63:0] _RAND_26;
  wire [40:0] _T_295; // @[Util.scala 113:33:@2857.4]
  reg [39:0] _T_297; // @[Util.scala 112:74:@2859.4]
  reg [63:0] _RAND_27;
  wire [40:0] _T_298; // @[Util.scala 113:33:@2860.4]
  reg [39:0] _T_300; // @[Util.scala 112:74:@2862.4]
  reg [63:0] _RAND_28;
  wire [40:0] _T_301; // @[Util.scala 113:33:@2863.4]
  reg [39:0] _T_303; // @[Util.scala 112:74:@2865.4]
  reg [63:0] _RAND_29;
  wire [40:0] _T_304; // @[Util.scala 113:33:@2866.4]
  reg [39:0] _T_306; // @[Util.scala 112:74:@2868.4]
  reg [63:0] _RAND_30;
  wire [40:0] _T_307; // @[Util.scala 113:33:@2869.4]
  reg [39:0] _T_309; // @[Util.scala 112:74:@2871.4]
  reg [63:0] _RAND_31;
  wire [40:0] _T_310; // @[Util.scala 113:33:@2872.4]
  reg [39:0] _T_312; // @[Util.scala 112:74:@2874.4]
  reg [63:0] _RAND_32;
  wire [40:0] _T_313; // @[Util.scala 113:33:@2875.4]
  reg [39:0] _T_315; // @[Util.scala 112:74:@2877.4]
  reg [63:0] _RAND_33;
  wire [40:0] _T_316; // @[Util.scala 113:33:@2878.4]
  reg [39:0] _T_318; // @[Util.scala 112:74:@2880.4]
  reg [63:0] _RAND_34;
  wire [40:0] _T_319; // @[Util.scala 113:33:@2881.4]
  reg [39:0] _T_321; // @[Util.scala 112:74:@2883.4]
  reg [63:0] _RAND_35;
  wire [40:0] _T_322; // @[Util.scala 113:33:@2884.4]
  reg [39:0] _T_324; // @[Util.scala 112:74:@2886.4]
  reg [63:0] _RAND_36;
  wire [40:0] _T_325; // @[Util.scala 113:33:@2887.4]
  reg [39:0] _T_327; // @[Util.scala 112:74:@2889.4]
  reg [63:0] _RAND_37;
  wire [40:0] _T_328; // @[Util.scala 113:33:@2890.4]
  reg [39:0] _T_330; // @[Util.scala 112:74:@2892.4]
  reg [63:0] _RAND_38;
  wire [40:0] _T_331; // @[Util.scala 113:33:@2893.4]
  reg [39:0] _T_333; // @[Util.scala 112:74:@2895.4]
  reg [63:0] _RAND_39;
  wire [40:0] _T_334; // @[Util.scala 113:33:@2896.4]
  reg [39:0] _T_336; // @[Util.scala 112:74:@2898.4]
  reg [63:0] _RAND_40;
  wire [40:0] _T_337; // @[Util.scala 113:33:@2899.4]
  reg [39:0] _T_339; // @[Util.scala 112:74:@2901.4]
  reg [63:0] _RAND_41;
  wire [40:0] _T_340; // @[Util.scala 113:33:@2902.4]
  reg [39:0] _T_342; // @[Util.scala 112:74:@2904.4]
  reg [63:0] _RAND_42;
  wire [40:0] _T_343; // @[Util.scala 113:33:@2905.4]
  reg [39:0] _T_345; // @[Util.scala 112:74:@2907.4]
  reg [63:0] _RAND_43;
  wire [40:0] _T_346; // @[Util.scala 113:33:@2908.4]
  reg [39:0] _T_348; // @[Util.scala 112:74:@2910.4]
  reg [63:0] _RAND_44;
  wire [40:0] _T_349; // @[Util.scala 113:33:@2911.4]
  reg [39:0] _T_351; // @[Util.scala 112:74:@2913.4]
  reg [63:0] _RAND_45;
  wire [40:0] _T_352; // @[Util.scala 113:33:@2914.4]
  reg [39:0] _T_354; // @[Util.scala 112:74:@2916.4]
  reg [63:0] _RAND_46;
  wire [40:0] _T_355; // @[Util.scala 113:33:@2917.4]
  reg [39:0] _T_357; // @[Util.scala 112:74:@2919.4]
  reg [63:0] _RAND_47;
  wire [40:0] _T_358; // @[Util.scala 113:33:@2920.4]
  reg [31:0] reg_dscratch; // @[CSR.scala 134:25:@3009.4]
  reg [31:0] _RAND_48;
  wire  system_insn; // @[CSR.scala 137:31:@3011.4]
  wire  _T_446; // @[CSR.scala 138:27:@3012.4]
  wire  _T_448; // @[CSR.scala 138:40:@3013.4]
  wire  cpu_ren; // @[CSR.scala 138:37:@3014.4]
  wire [31:0] read_mstatus; // @[CSR.scala 140:32:@3023.4]
  wire [15:0] _T_468; // @[CSR.scala 156:25:@3029.4]
  wire [15:0] _T_474; // @[CSR.scala 157:25:@3035.4]
  wire  _T_478; // @[CSR.scala 177:73:@3036.4]
  wire  _T_480; // @[CSR.scala 177:73:@3037.4]
  wire  _T_482; // @[CSR.scala 177:73:@3038.4]
  wire  _T_488; // @[CSR.scala 177:73:@3041.4]
  wire  _T_490; // @[CSR.scala 177:73:@3042.4]
  wire  _T_492; // @[CSR.scala 177:73:@3043.4]
  wire  _T_494; // @[CSR.scala 177:73:@3044.4]
  wire  _T_496; // @[CSR.scala 177:73:@3045.4]
  wire  _T_498; // @[CSR.scala 177:73:@3046.4]
  wire  _T_500; // @[CSR.scala 177:73:@3047.4]
  wire  _T_502; // @[CSR.scala 177:73:@3048.4]
  wire  _T_504; // @[CSR.scala 177:73:@3049.4]
  wire  _T_508; // @[CSR.scala 177:73:@3051.4]
  wire  _T_510; // @[CSR.scala 177:73:@3052.4]
  wire  _T_512; // @[CSR.scala 177:73:@3053.4]
  wire  _T_514; // @[CSR.scala 177:73:@3054.4]
  wire  _T_516; // @[CSR.scala 177:73:@3055.4]
  wire  _T_518; // @[CSR.scala 177:73:@3056.4]
  wire  _T_520; // @[CSR.scala 177:73:@3057.4]
  wire  _T_522; // @[CSR.scala 177:73:@3058.4]
  wire  _T_524; // @[CSR.scala 177:73:@3059.4]
  wire  _T_526; // @[CSR.scala 177:73:@3060.4]
  wire  _T_528; // @[CSR.scala 177:73:@3061.4]
  wire  _T_530; // @[CSR.scala 177:73:@3062.4]
  wire  _T_532; // @[CSR.scala 177:73:@3063.4]
  wire  _T_534; // @[CSR.scala 177:73:@3064.4]
  wire  _T_536; // @[CSR.scala 177:73:@3065.4]
  wire  _T_538; // @[CSR.scala 177:73:@3066.4]
  wire  _T_540; // @[CSR.scala 177:73:@3067.4]
  wire  _T_542; // @[CSR.scala 177:73:@3068.4]
  wire  _T_544; // @[CSR.scala 177:73:@3069.4]
  wire  _T_546; // @[CSR.scala 177:73:@3070.4]
  wire  _T_548; // @[CSR.scala 177:73:@3071.4]
  wire  _T_550; // @[CSR.scala 177:73:@3072.4]
  wire  _T_552; // @[CSR.scala 177:73:@3073.4]
  wire  _T_554; // @[CSR.scala 177:73:@3074.4]
  wire  _T_556; // @[CSR.scala 177:73:@3075.4]
  wire  _T_558; // @[CSR.scala 177:73:@3076.4]
  wire  _T_560; // @[CSR.scala 177:73:@3077.4]
  wire  _T_562; // @[CSR.scala 177:73:@3078.4]
  wire  _T_564; // @[CSR.scala 177:73:@3079.4]
  wire  _T_566; // @[CSR.scala 177:73:@3080.4]
  wire  _T_568; // @[CSR.scala 177:73:@3081.4]
  wire  _T_570; // @[CSR.scala 177:73:@3082.4]
  wire  _T_572; // @[CSR.scala 177:73:@3083.4]
  wire  _T_574; // @[CSR.scala 177:73:@3084.4]
  wire  _T_576; // @[CSR.scala 177:73:@3085.4]
  wire  _T_578; // @[CSR.scala 177:73:@3086.4]
  wire  _T_580; // @[CSR.scala 177:73:@3087.4]
  wire  _T_582; // @[CSR.scala 177:73:@3088.4]
  wire  _T_584; // @[CSR.scala 177:73:@3089.4]
  wire  _T_586; // @[CSR.scala 177:73:@3090.4]
  wire  _T_588; // @[CSR.scala 177:73:@3091.4]
  wire  _T_590; // @[CSR.scala 177:73:@3092.4]
  wire  _T_592; // @[CSR.scala 177:73:@3093.4]
  wire  _T_594; // @[CSR.scala 177:73:@3094.4]
  wire  _T_596; // @[CSR.scala 177:73:@3095.4]
  wire  _T_598; // @[CSR.scala 177:73:@3096.4]
  wire  _T_600; // @[CSR.scala 177:73:@3097.4]
  wire  _T_602; // @[CSR.scala 177:73:@3098.4]
  wire  _T_604; // @[CSR.scala 177:73:@3099.4]
  wire  _T_606; // @[CSR.scala 177:73:@3100.4]
  wire  _T_608; // @[CSR.scala 177:73:@3101.4]
  wire  _T_610; // @[CSR.scala 177:73:@3102.4]
  wire  _T_612; // @[CSR.scala 177:73:@3103.4]
  wire  _T_614; // @[CSR.scala 177:73:@3104.4]
  wire  _T_616; // @[CSR.scala 177:73:@3105.4]
  wire  _T_618; // @[CSR.scala 177:73:@3106.4]
  wire  _T_620; // @[CSR.scala 177:73:@3107.4]
  wire  _T_622; // @[CSR.scala 177:73:@3108.4]
  wire  _T_624; // @[CSR.scala 177:73:@3109.4]
  wire  _T_626; // @[CSR.scala 177:73:@3110.4]
  wire  _T_628; // @[CSR.scala 177:73:@3111.4]
  wire  _T_630; // @[CSR.scala 177:73:@3112.4]
  wire  _T_632; // @[CSR.scala 177:73:@3113.4]
  wire  _T_634; // @[CSR.scala 177:73:@3114.4]
  wire  _T_636; // @[CSR.scala 177:73:@3115.4]
  wire  _T_638; // @[CSR.scala 177:73:@3116.4]
  wire  _T_640; // @[CSR.scala 177:73:@3117.4]
  wire  _T_642; // @[CSR.scala 177:73:@3118.4]
  wire [1:0] _T_643; // @[CSR.scala 179:54:@3119.4]
  wire  priv_sufficient; // @[CSR.scala 179:41:@3120.4]
  wire [1:0] _T_644; // @[CSR.scala 180:29:@3121.4]
  wire [1:0] _T_645; // @[CSR.scala 180:37:@3122.4]
  wire  read_only; // @[CSR.scala 180:37:@3123.4]
  wire  _T_647; // @[CSR.scala 181:38:@3124.4]
  wire  _T_648; // @[CSR.scala 181:25:@3125.4]
  wire  cpu_wen; // @[CSR.scala 181:48:@3126.4]
  wire  _T_650; // @[CSR.scala 182:24:@3127.4]
  wire  wen; // @[CSR.scala 182:21:@3128.4]
  wire  _T_651; // @[Util.scala 23:47:@3129.4]
  wire  _T_652; // @[Util.scala 23:47:@3130.4]
  wire  _T_653; // @[Util.scala 23:62:@3131.4]
  wire [31:0] _T_655; // @[CSR.scala 281:9:@3132.4]
  wire [31:0] _T_656; // @[CSR.scala 281:49:@3133.4]
  wire [31:0] _T_659; // @[CSR.scala 281:64:@3135.4]
  wire [31:0] _T_660; // @[CSR.scala 281:60:@3136.4]
  wire [31:0] wdata; // @[CSR.scala 281:58:@3137.4]
  wire [2:0] _T_662; // @[CSR.scala 185:33:@3138.4]
  wire [7:0] opcode; // @[CSR.scala 185:20:@3139.4]
  wire  _T_663; // @[CSR.scala 186:40:@3140.4]
  wire  insn_call; // @[CSR.scala 186:31:@3141.4]
  wire  _T_664; // @[CSR.scala 187:41:@3142.4]
  wire  insn_break; // @[CSR.scala 187:32:@3143.4]
  wire  _T_665; // @[CSR.scala 188:39:@3144.4]
  wire  _T_666; // @[CSR.scala 188:30:@3145.4]
  wire  insn_ret; // @[CSR.scala 188:43:@3146.4]
  wire  _T_940; // @[CSR.scala 199:24:@3345.4]
  wire [1:0] _T_942; // @[Bitwise.scala 48:55:@3348.4]
  wire  _T_944; // @[CSR.scala 201:50:@3349.4]
  wire  _T_946; // @[CSR.scala 201:9:@3351.4]
  wire  _T_948; // @[CSR.scala 201:9:@3352.4]
  wire  _T_951; // @[CSR.scala 208:32:@3361.4]
  wire  _T_953; // @[CSR.scala 208:21:@3362.4]
  wire  _T_954; // @[CSR.scala 208:18:@3363.4]
  wire  _GEN_3; // @[CSR.scala 208:38:@3364.4]
  wire  _GEN_4; // @[CSR.scala 208:38:@3364.4]
  wire [1:0] new_prv; // @[CSR.scala 208:38:@3364.4]
  wire [3:0] _GEN_148; // @[CSR.scala 218:35:@3372.6]
  wire [4:0] _T_958; // @[CSR.scala 218:35:@3372.6]
  wire [3:0] _T_959; // @[CSR.scala 218:35:@3373.6]
  wire [31:0] _GEN_7; // @[CSR.scala 216:18:@3370.4]
  wire [31:0] _GEN_8; // @[CSR.scala 216:18:@3370.4]
  wire [31:0] _GEN_9; // @[CSR.scala 216:18:@3370.4]
  wire [31:0] _GEN_10; // @[CSR.scala 223:19:@3377.4]
  wire [31:0] _GEN_11; // @[CSR.scala 223:19:@3377.4]
  wire [31:0] _GEN_12; // @[CSR.scala 223:19:@3377.4]
  wire [31:0] _GEN_14; // @[CSR.scala 229:17:@3382.4]
  wire [31:0] _GEN_15; // @[CSR.scala 229:17:@3382.4]
  wire [31:0] _GEN_16; // @[CSR.scala 229:17:@3382.4]
  wire [63:0] _T_965; // @[Mux.scala 19:72:@3390.4]
  wire [63:0] _T_967; // @[Mux.scala 19:72:@3391.4]
  wire [15:0] _T_969; // @[Mux.scala 19:72:@3392.4]
  wire [30:0] _T_975; // @[Mux.scala 19:72:@3395.4]
  wire [31:0] _T_977; // @[Mux.scala 19:72:@3396.4]
  wire [8:0] _T_979; // @[Mux.scala 19:72:@3397.4]
  wire [15:0] _T_981; // @[Mux.scala 19:72:@3398.4]
  wire [15:0] _T_983; // @[Mux.scala 19:72:@3399.4]
  wire [31:0] _T_985; // @[Mux.scala 19:72:@3400.4]
  wire [31:0] _T_987; // @[Mux.scala 19:72:@3401.4]
  wire [31:0] _T_989; // @[Mux.scala 19:72:@3402.4]
  wire [31:0] _T_991; // @[Mux.scala 19:72:@3403.4]
  wire [31:0] _T_995; // @[Mux.scala 19:72:@3405.4]
  wire [31:0] _T_997; // @[Mux.scala 19:72:@3406.4]
  wire [39:0] _T_999; // @[Mux.scala 19:72:@3407.4]
  wire [39:0] _T_1001; // @[Mux.scala 19:72:@3408.4]
  wire [39:0] _T_1003; // @[Mux.scala 19:72:@3409.4]
  wire [39:0] _T_1005; // @[Mux.scala 19:72:@3410.4]
  wire [39:0] _T_1007; // @[Mux.scala 19:72:@3411.4]
  wire [39:0] _T_1009; // @[Mux.scala 19:72:@3412.4]
  wire [39:0] _T_1011; // @[Mux.scala 19:72:@3413.4]
  wire [39:0] _T_1013; // @[Mux.scala 19:72:@3414.4]
  wire [39:0] _T_1015; // @[Mux.scala 19:72:@3415.4]
  wire [39:0] _T_1017; // @[Mux.scala 19:72:@3416.4]
  wire [39:0] _T_1019; // @[Mux.scala 19:72:@3417.4]
  wire [39:0] _T_1021; // @[Mux.scala 19:72:@3418.4]
  wire [39:0] _T_1023; // @[Mux.scala 19:72:@3419.4]
  wire [39:0] _T_1025; // @[Mux.scala 19:72:@3420.4]
  wire [39:0] _T_1027; // @[Mux.scala 19:72:@3421.4]
  wire [39:0] _T_1029; // @[Mux.scala 19:72:@3422.4]
  wire [39:0] _T_1031; // @[Mux.scala 19:72:@3423.4]
  wire [39:0] _T_1033; // @[Mux.scala 19:72:@3424.4]
  wire [39:0] _T_1035; // @[Mux.scala 19:72:@3425.4]
  wire [39:0] _T_1037; // @[Mux.scala 19:72:@3426.4]
  wire [39:0] _T_1039; // @[Mux.scala 19:72:@3427.4]
  wire [39:0] _T_1041; // @[Mux.scala 19:72:@3428.4]
  wire [39:0] _T_1043; // @[Mux.scala 19:72:@3429.4]
  wire [39:0] _T_1045; // @[Mux.scala 19:72:@3430.4]
  wire [39:0] _T_1047; // @[Mux.scala 19:72:@3431.4]
  wire [39:0] _T_1049; // @[Mux.scala 19:72:@3432.4]
  wire [39:0] _T_1051; // @[Mux.scala 19:72:@3433.4]
  wire [39:0] _T_1053; // @[Mux.scala 19:72:@3434.4]
  wire [39:0] _T_1055; // @[Mux.scala 19:72:@3435.4]
  wire [39:0] _T_1057; // @[Mux.scala 19:72:@3436.4]
  wire [39:0] _T_1059; // @[Mux.scala 19:72:@3437.4]
  wire [39:0] _T_1061; // @[Mux.scala 19:72:@3438.4]
  wire [39:0] _T_1063; // @[Mux.scala 19:72:@3439.4]
  wire [39:0] _T_1065; // @[Mux.scala 19:72:@3440.4]
  wire [39:0] _T_1067; // @[Mux.scala 19:72:@3441.4]
  wire [39:0] _T_1069; // @[Mux.scala 19:72:@3442.4]
  wire [39:0] _T_1071; // @[Mux.scala 19:72:@3443.4]
  wire [39:0] _T_1073; // @[Mux.scala 19:72:@3444.4]
  wire [39:0] _T_1075; // @[Mux.scala 19:72:@3445.4]
  wire [39:0] _T_1077; // @[Mux.scala 19:72:@3446.4]
  wire [39:0] _T_1079; // @[Mux.scala 19:72:@3447.4]
  wire [39:0] _T_1081; // @[Mux.scala 19:72:@3448.4]
  wire [39:0] _T_1083; // @[Mux.scala 19:72:@3449.4]
  wire [39:0] _T_1085; // @[Mux.scala 19:72:@3450.4]
  wire [39:0] _T_1087; // @[Mux.scala 19:72:@3451.4]
  wire [39:0] _T_1089; // @[Mux.scala 19:72:@3452.4]
  wire [39:0] _T_1091; // @[Mux.scala 19:72:@3453.4]
  wire [39:0] _T_1093; // @[Mux.scala 19:72:@3454.4]
  wire [39:0] _T_1095; // @[Mux.scala 19:72:@3455.4]
  wire [39:0] _T_1097; // @[Mux.scala 19:72:@3456.4]
  wire [39:0] _T_1099; // @[Mux.scala 19:72:@3457.4]
  wire [39:0] _T_1101; // @[Mux.scala 19:72:@3458.4]
  wire [39:0] _T_1103; // @[Mux.scala 19:72:@3459.4]
  wire [39:0] _T_1105; // @[Mux.scala 19:72:@3460.4]
  wire [39:0] _T_1107; // @[Mux.scala 19:72:@3461.4]
  wire [39:0] _T_1109; // @[Mux.scala 19:72:@3462.4]
  wire [39:0] _T_1111; // @[Mux.scala 19:72:@3463.4]
  wire [39:0] _T_1113; // @[Mux.scala 19:72:@3464.4]
  wire [39:0] _T_1115; // @[Mux.scala 19:72:@3465.4]
  wire [39:0] _T_1117; // @[Mux.scala 19:72:@3466.4]
  wire [39:0] _T_1119; // @[Mux.scala 19:72:@3467.4]
  wire [39:0] _T_1121; // @[Mux.scala 19:72:@3468.4]
  wire [39:0] _T_1123; // @[Mux.scala 19:72:@3469.4]
  wire [39:0] _T_1125; // @[Mux.scala 19:72:@3470.4]
  wire [63:0] _T_1130; // @[Mux.scala 19:72:@3473.4]
  wire [63:0] _GEN_149; // @[Mux.scala 19:72:@3474.4]
  wire [63:0] _T_1131; // @[Mux.scala 19:72:@3474.4]
  wire [63:0] _GEN_150; // @[Mux.scala 19:72:@3477.4]
  wire [63:0] _T_1134; // @[Mux.scala 19:72:@3477.4]
  wire [63:0] _GEN_151; // @[Mux.scala 19:72:@3478.4]
  wire [63:0] _T_1135; // @[Mux.scala 19:72:@3478.4]
  wire [63:0] _GEN_152; // @[Mux.scala 19:72:@3479.4]
  wire [63:0] _T_1136; // @[Mux.scala 19:72:@3479.4]
  wire [63:0] _GEN_153; // @[Mux.scala 19:72:@3480.4]
  wire [63:0] _T_1137; // @[Mux.scala 19:72:@3480.4]
  wire [63:0] _GEN_154; // @[Mux.scala 19:72:@3481.4]
  wire [63:0] _T_1138; // @[Mux.scala 19:72:@3481.4]
  wire [63:0] _GEN_155; // @[Mux.scala 19:72:@3482.4]
  wire [63:0] _T_1139; // @[Mux.scala 19:72:@3482.4]
  wire [63:0] _GEN_156; // @[Mux.scala 19:72:@3483.4]
  wire [63:0] _T_1140; // @[Mux.scala 19:72:@3483.4]
  wire [63:0] _GEN_157; // @[Mux.scala 19:72:@3484.4]
  wire [63:0] _T_1141; // @[Mux.scala 19:72:@3484.4]
  wire [63:0] _GEN_158; // @[Mux.scala 19:72:@3485.4]
  wire [63:0] _T_1142; // @[Mux.scala 19:72:@3485.4]
  wire [63:0] _GEN_159; // @[Mux.scala 19:72:@3487.4]
  wire [63:0] _T_1144; // @[Mux.scala 19:72:@3487.4]
  wire [63:0] _GEN_160; // @[Mux.scala 19:72:@3488.4]
  wire [63:0] _T_1145; // @[Mux.scala 19:72:@3488.4]
  wire [63:0] _GEN_161; // @[Mux.scala 19:72:@3489.4]
  wire [63:0] _T_1146; // @[Mux.scala 19:72:@3489.4]
  wire [63:0] _GEN_162; // @[Mux.scala 19:72:@3490.4]
  wire [63:0] _T_1147; // @[Mux.scala 19:72:@3490.4]
  wire [63:0] _GEN_163; // @[Mux.scala 19:72:@3491.4]
  wire [63:0] _T_1148; // @[Mux.scala 19:72:@3491.4]
  wire [63:0] _GEN_164; // @[Mux.scala 19:72:@3492.4]
  wire [63:0] _T_1149; // @[Mux.scala 19:72:@3492.4]
  wire [63:0] _GEN_165; // @[Mux.scala 19:72:@3493.4]
  wire [63:0] _T_1150; // @[Mux.scala 19:72:@3493.4]
  wire [63:0] _GEN_166; // @[Mux.scala 19:72:@3494.4]
  wire [63:0] _T_1151; // @[Mux.scala 19:72:@3494.4]
  wire [63:0] _GEN_167; // @[Mux.scala 19:72:@3495.4]
  wire [63:0] _T_1152; // @[Mux.scala 19:72:@3495.4]
  wire [63:0] _GEN_168; // @[Mux.scala 19:72:@3496.4]
  wire [63:0] _T_1153; // @[Mux.scala 19:72:@3496.4]
  wire [63:0] _GEN_169; // @[Mux.scala 19:72:@3497.4]
  wire [63:0] _T_1154; // @[Mux.scala 19:72:@3497.4]
  wire [63:0] _GEN_170; // @[Mux.scala 19:72:@3498.4]
  wire [63:0] _T_1155; // @[Mux.scala 19:72:@3498.4]
  wire [63:0] _GEN_171; // @[Mux.scala 19:72:@3499.4]
  wire [63:0] _T_1156; // @[Mux.scala 19:72:@3499.4]
  wire [63:0] _GEN_172; // @[Mux.scala 19:72:@3500.4]
  wire [63:0] _T_1157; // @[Mux.scala 19:72:@3500.4]
  wire [63:0] _GEN_173; // @[Mux.scala 19:72:@3501.4]
  wire [63:0] _T_1158; // @[Mux.scala 19:72:@3501.4]
  wire [63:0] _GEN_174; // @[Mux.scala 19:72:@3502.4]
  wire [63:0] _T_1159; // @[Mux.scala 19:72:@3502.4]
  wire [63:0] _GEN_175; // @[Mux.scala 19:72:@3503.4]
  wire [63:0] _T_1160; // @[Mux.scala 19:72:@3503.4]
  wire [63:0] _GEN_176; // @[Mux.scala 19:72:@3504.4]
  wire [63:0] _T_1161; // @[Mux.scala 19:72:@3504.4]
  wire [63:0] _GEN_177; // @[Mux.scala 19:72:@3505.4]
  wire [63:0] _T_1162; // @[Mux.scala 19:72:@3505.4]
  wire [63:0] _GEN_178; // @[Mux.scala 19:72:@3506.4]
  wire [63:0] _T_1163; // @[Mux.scala 19:72:@3506.4]
  wire [63:0] _GEN_179; // @[Mux.scala 19:72:@3507.4]
  wire [63:0] _T_1164; // @[Mux.scala 19:72:@3507.4]
  wire [63:0] _GEN_180; // @[Mux.scala 19:72:@3508.4]
  wire [63:0] _T_1165; // @[Mux.scala 19:72:@3508.4]
  wire [63:0] _GEN_181; // @[Mux.scala 19:72:@3509.4]
  wire [63:0] _T_1166; // @[Mux.scala 19:72:@3509.4]
  wire [63:0] _GEN_182; // @[Mux.scala 19:72:@3510.4]
  wire [63:0] _T_1167; // @[Mux.scala 19:72:@3510.4]
  wire [63:0] _GEN_183; // @[Mux.scala 19:72:@3511.4]
  wire [63:0] _T_1168; // @[Mux.scala 19:72:@3511.4]
  wire [63:0] _GEN_184; // @[Mux.scala 19:72:@3512.4]
  wire [63:0] _T_1169; // @[Mux.scala 19:72:@3512.4]
  wire [63:0] _GEN_185; // @[Mux.scala 19:72:@3513.4]
  wire [63:0] _T_1170; // @[Mux.scala 19:72:@3513.4]
  wire [63:0] _GEN_186; // @[Mux.scala 19:72:@3514.4]
  wire [63:0] _T_1171; // @[Mux.scala 19:72:@3514.4]
  wire [63:0] _GEN_187; // @[Mux.scala 19:72:@3515.4]
  wire [63:0] _T_1172; // @[Mux.scala 19:72:@3515.4]
  wire [63:0] _GEN_188; // @[Mux.scala 19:72:@3516.4]
  wire [63:0] _T_1173; // @[Mux.scala 19:72:@3516.4]
  wire [63:0] _GEN_189; // @[Mux.scala 19:72:@3517.4]
  wire [63:0] _T_1174; // @[Mux.scala 19:72:@3517.4]
  wire [63:0] _GEN_190; // @[Mux.scala 19:72:@3518.4]
  wire [63:0] _T_1175; // @[Mux.scala 19:72:@3518.4]
  wire [63:0] _GEN_191; // @[Mux.scala 19:72:@3519.4]
  wire [63:0] _T_1176; // @[Mux.scala 19:72:@3519.4]
  wire [63:0] _GEN_192; // @[Mux.scala 19:72:@3520.4]
  wire [63:0] _T_1177; // @[Mux.scala 19:72:@3520.4]
  wire [63:0] _GEN_193; // @[Mux.scala 19:72:@3521.4]
  wire [63:0] _T_1178; // @[Mux.scala 19:72:@3521.4]
  wire [63:0] _GEN_194; // @[Mux.scala 19:72:@3522.4]
  wire [63:0] _T_1179; // @[Mux.scala 19:72:@3522.4]
  wire [63:0] _GEN_195; // @[Mux.scala 19:72:@3523.4]
  wire [63:0] _T_1180; // @[Mux.scala 19:72:@3523.4]
  wire [63:0] _GEN_196; // @[Mux.scala 19:72:@3524.4]
  wire [63:0] _T_1181; // @[Mux.scala 19:72:@3524.4]
  wire [63:0] _GEN_197; // @[Mux.scala 19:72:@3525.4]
  wire [63:0] _T_1182; // @[Mux.scala 19:72:@3525.4]
  wire [63:0] _GEN_198; // @[Mux.scala 19:72:@3526.4]
  wire [63:0] _T_1183; // @[Mux.scala 19:72:@3526.4]
  wire [63:0] _GEN_199; // @[Mux.scala 19:72:@3527.4]
  wire [63:0] _T_1184; // @[Mux.scala 19:72:@3527.4]
  wire [63:0] _GEN_200; // @[Mux.scala 19:72:@3528.4]
  wire [63:0] _T_1185; // @[Mux.scala 19:72:@3528.4]
  wire [63:0] _GEN_201; // @[Mux.scala 19:72:@3529.4]
  wire [63:0] _T_1186; // @[Mux.scala 19:72:@3529.4]
  wire [63:0] _GEN_202; // @[Mux.scala 19:72:@3530.4]
  wire [63:0] _T_1187; // @[Mux.scala 19:72:@3530.4]
  wire [63:0] _GEN_203; // @[Mux.scala 19:72:@3531.4]
  wire [63:0] _T_1188; // @[Mux.scala 19:72:@3531.4]
  wire [63:0] _GEN_204; // @[Mux.scala 19:72:@3532.4]
  wire [63:0] _T_1189; // @[Mux.scala 19:72:@3532.4]
  wire [63:0] _GEN_205; // @[Mux.scala 19:72:@3533.4]
  wire [63:0] _T_1190; // @[Mux.scala 19:72:@3533.4]
  wire [63:0] _GEN_206; // @[Mux.scala 19:72:@3534.4]
  wire [63:0] _T_1191; // @[Mux.scala 19:72:@3534.4]
  wire [63:0] _GEN_207; // @[Mux.scala 19:72:@3535.4]
  wire [63:0] _T_1192; // @[Mux.scala 19:72:@3535.4]
  wire [63:0] _GEN_208; // @[Mux.scala 19:72:@3536.4]
  wire [63:0] _T_1193; // @[Mux.scala 19:72:@3536.4]
  wire [63:0] _GEN_209; // @[Mux.scala 19:72:@3537.4]
  wire [63:0] _T_1194; // @[Mux.scala 19:72:@3537.4]
  wire [63:0] _GEN_210; // @[Mux.scala 19:72:@3538.4]
  wire [63:0] _T_1195; // @[Mux.scala 19:72:@3538.4]
  wire [63:0] _GEN_211; // @[Mux.scala 19:72:@3539.4]
  wire [63:0] _T_1196; // @[Mux.scala 19:72:@3539.4]
  wire [63:0] _GEN_212; // @[Mux.scala 19:72:@3540.4]
  wire [63:0] _T_1197; // @[Mux.scala 19:72:@3540.4]
  wire [63:0] _GEN_213; // @[Mux.scala 19:72:@3541.4]
  wire [63:0] _T_1198; // @[Mux.scala 19:72:@3541.4]
  wire [63:0] _GEN_214; // @[Mux.scala 19:72:@3542.4]
  wire [63:0] _T_1199; // @[Mux.scala 19:72:@3542.4]
  wire [63:0] _GEN_215; // @[Mux.scala 19:72:@3543.4]
  wire [63:0] _T_1200; // @[Mux.scala 19:72:@3543.4]
  wire [63:0] _GEN_216; // @[Mux.scala 19:72:@3544.4]
  wire [63:0] _T_1201; // @[Mux.scala 19:72:@3544.4]
  wire [63:0] _GEN_217; // @[Mux.scala 19:72:@3545.4]
  wire [63:0] _T_1202; // @[Mux.scala 19:72:@3545.4]
  wire [63:0] _GEN_218; // @[Mux.scala 19:72:@3546.4]
  wire [63:0] _T_1203; // @[Mux.scala 19:72:@3546.4]
  wire [63:0] _GEN_219; // @[Mux.scala 19:72:@3547.4]
  wire [63:0] _T_1204; // @[Mux.scala 19:72:@3547.4]
  wire [63:0] _GEN_220; // @[Mux.scala 19:72:@3548.4]
  wire [63:0] _T_1205; // @[Mux.scala 19:72:@3548.4]
  wire [63:0] _GEN_221; // @[Mux.scala 19:72:@3549.4]
  wire [63:0] _T_1206; // @[Mux.scala 19:72:@3549.4]
  wire [63:0] _GEN_222; // @[Mux.scala 19:72:@3550.4]
  wire [63:0] _T_1207; // @[Mux.scala 19:72:@3550.4]
  wire [63:0] _GEN_223; // @[Mux.scala 19:72:@3551.4]
  wire [63:0] _T_1208; // @[Mux.scala 19:72:@3551.4]
  wire [63:0] _GEN_224; // @[Mux.scala 19:72:@3552.4]
  wire [63:0] _T_1209; // @[Mux.scala 19:72:@3552.4]
  wire  _T_1220; // @[CSR.scala 245:39:@3565.8]
  wire  _T_1222; // @[CSR.scala 245:39:@3569.8]
  wire  _GEN_17; // @[CSR.scala 244:39:@3559.6]
  wire  _GEN_18; // @[CSR.scala 244:39:@3559.6]
  wire [15:0] _T_1233; // @[:@3588.8 :@3589.8]
  wire  _T_1235; // @[CSR.scala 250:35:@3592.8]
  wire  _T_1237; // @[CSR.scala 250:35:@3596.8]
  wire  _GEN_19; // @[CSR.scala 249:35:@3586.6]
  wire  _GEN_20; // @[CSR.scala 253:35:@3606.6]
  wire  _GEN_21; // @[CSR.scala 253:35:@3606.6]
  wire [7:0] _T_1253; // @[CSR.scala 277:47:@3628.8]
  wire [31:0] _T_1254; // @[CSR.scala 277:72:@3629.8]
  wire [39:0] _T_1255; // @[Cat.scala 30:58:@3630.8]
  wire [40:0] _GEN_22; // @[CSR.scala 277:29:@3627.6]
  wire [7:0] _T_1256; // @[CSR.scala 278:45:@3634.8]
  wire [39:0] _T_1257; // @[Cat.scala 30:58:@3635.8]
  wire [40:0] _GEN_23; // @[CSR.scala 278:29:@3633.6]
  wire [31:0] _T_1259; // @[CSR.scala 277:72:@3640.8]
  wire [39:0] _T_1260; // @[Cat.scala 30:58:@3641.8]
  wire [40:0] _GEN_24; // @[CSR.scala 277:29:@3638.6]
  wire [7:0] _T_1261; // @[CSR.scala 278:45:@3645.8]
  wire [39:0] _T_1262; // @[Cat.scala 30:58:@3646.8]
  wire [40:0] _GEN_25; // @[CSR.scala 278:29:@3644.6]
  wire [31:0] _T_1264; // @[CSR.scala 277:72:@3651.8]
  wire [39:0] _T_1265; // @[Cat.scala 30:58:@3652.8]
  wire [40:0] _GEN_26; // @[CSR.scala 277:29:@3649.6]
  wire [7:0] _T_1266; // @[CSR.scala 278:45:@3656.8]
  wire [39:0] _T_1267; // @[Cat.scala 30:58:@3657.8]
  wire [40:0] _GEN_27; // @[CSR.scala 278:29:@3655.6]
  wire [31:0] _T_1269; // @[CSR.scala 277:72:@3662.8]
  wire [39:0] _T_1270; // @[Cat.scala 30:58:@3663.8]
  wire [40:0] _GEN_28; // @[CSR.scala 277:29:@3660.6]
  wire [7:0] _T_1271; // @[CSR.scala 278:45:@3667.8]
  wire [39:0] _T_1272; // @[Cat.scala 30:58:@3668.8]
  wire [40:0] _GEN_29; // @[CSR.scala 278:29:@3666.6]
  wire [31:0] _T_1274; // @[CSR.scala 277:72:@3673.8]
  wire [39:0] _T_1275; // @[Cat.scala 30:58:@3674.8]
  wire [40:0] _GEN_30; // @[CSR.scala 277:29:@3671.6]
  wire [7:0] _T_1276; // @[CSR.scala 278:45:@3678.8]
  wire [39:0] _T_1277; // @[Cat.scala 30:58:@3679.8]
  wire [40:0] _GEN_31; // @[CSR.scala 278:29:@3677.6]
  wire [31:0] _T_1279; // @[CSR.scala 277:72:@3684.8]
  wire [39:0] _T_1280; // @[Cat.scala 30:58:@3685.8]
  wire [40:0] _GEN_32; // @[CSR.scala 277:29:@3682.6]
  wire [7:0] _T_1281; // @[CSR.scala 278:45:@3689.8]
  wire [39:0] _T_1282; // @[Cat.scala 30:58:@3690.8]
  wire [40:0] _GEN_33; // @[CSR.scala 278:29:@3688.6]
  wire [31:0] _T_1284; // @[CSR.scala 277:72:@3695.8]
  wire [39:0] _T_1285; // @[Cat.scala 30:58:@3696.8]
  wire [40:0] _GEN_34; // @[CSR.scala 277:29:@3693.6]
  wire [7:0] _T_1286; // @[CSR.scala 278:45:@3700.8]
  wire [39:0] _T_1287; // @[Cat.scala 30:58:@3701.8]
  wire [40:0] _GEN_35; // @[CSR.scala 278:29:@3699.6]
  wire [31:0] _T_1289; // @[CSR.scala 277:72:@3706.8]
  wire [39:0] _T_1290; // @[Cat.scala 30:58:@3707.8]
  wire [40:0] _GEN_36; // @[CSR.scala 277:29:@3704.6]
  wire [7:0] _T_1291; // @[CSR.scala 278:45:@3711.8]
  wire [39:0] _T_1292; // @[Cat.scala 30:58:@3712.8]
  wire [40:0] _GEN_37; // @[CSR.scala 278:29:@3710.6]
  wire [31:0] _T_1294; // @[CSR.scala 277:72:@3717.8]
  wire [39:0] _T_1295; // @[Cat.scala 30:58:@3718.8]
  wire [40:0] _GEN_38; // @[CSR.scala 277:29:@3715.6]
  wire [7:0] _T_1296; // @[CSR.scala 278:45:@3722.8]
  wire [39:0] _T_1297; // @[Cat.scala 30:58:@3723.8]
  wire [40:0] _GEN_39; // @[CSR.scala 278:29:@3721.6]
  wire [31:0] _T_1299; // @[CSR.scala 277:72:@3728.8]
  wire [39:0] _T_1300; // @[Cat.scala 30:58:@3729.8]
  wire [40:0] _GEN_40; // @[CSR.scala 277:29:@3726.6]
  wire [7:0] _T_1301; // @[CSR.scala 278:45:@3733.8]
  wire [39:0] _T_1302; // @[Cat.scala 30:58:@3734.8]
  wire [40:0] _GEN_41; // @[CSR.scala 278:29:@3732.6]
  wire [31:0] _T_1304; // @[CSR.scala 277:72:@3739.8]
  wire [39:0] _T_1305; // @[Cat.scala 30:58:@3740.8]
  wire [40:0] _GEN_42; // @[CSR.scala 277:29:@3737.6]
  wire [7:0] _T_1306; // @[CSR.scala 278:45:@3744.8]
  wire [39:0] _T_1307; // @[Cat.scala 30:58:@3745.8]
  wire [40:0] _GEN_43; // @[CSR.scala 278:29:@3743.6]
  wire [31:0] _T_1309; // @[CSR.scala 277:72:@3750.8]
  wire [39:0] _T_1310; // @[Cat.scala 30:58:@3751.8]
  wire [40:0] _GEN_44; // @[CSR.scala 277:29:@3748.6]
  wire [7:0] _T_1311; // @[CSR.scala 278:45:@3755.8]
  wire [39:0] _T_1312; // @[Cat.scala 30:58:@3756.8]
  wire [40:0] _GEN_45; // @[CSR.scala 278:29:@3754.6]
  wire [31:0] _T_1314; // @[CSR.scala 277:72:@3761.8]
  wire [39:0] _T_1315; // @[Cat.scala 30:58:@3762.8]
  wire [40:0] _GEN_46; // @[CSR.scala 277:29:@3759.6]
  wire [7:0] _T_1316; // @[CSR.scala 278:45:@3766.8]
  wire [39:0] _T_1317; // @[Cat.scala 30:58:@3767.8]
  wire [40:0] _GEN_47; // @[CSR.scala 278:29:@3765.6]
  wire [31:0] _T_1319; // @[CSR.scala 277:72:@3772.8]
  wire [39:0] _T_1320; // @[Cat.scala 30:58:@3773.8]
  wire [40:0] _GEN_48; // @[CSR.scala 277:29:@3770.6]
  wire [7:0] _T_1321; // @[CSR.scala 278:45:@3777.8]
  wire [39:0] _T_1322; // @[Cat.scala 30:58:@3778.8]
  wire [40:0] _GEN_49; // @[CSR.scala 278:29:@3776.6]
  wire [31:0] _T_1324; // @[CSR.scala 277:72:@3783.8]
  wire [39:0] _T_1325; // @[Cat.scala 30:58:@3784.8]
  wire [40:0] _GEN_50; // @[CSR.scala 277:29:@3781.6]
  wire [7:0] _T_1326; // @[CSR.scala 278:45:@3788.8]
  wire [39:0] _T_1327; // @[Cat.scala 30:58:@3789.8]
  wire [40:0] _GEN_51; // @[CSR.scala 278:29:@3787.6]
  wire [31:0] _T_1329; // @[CSR.scala 277:72:@3794.8]
  wire [39:0] _T_1330; // @[Cat.scala 30:58:@3795.8]
  wire [40:0] _GEN_52; // @[CSR.scala 277:29:@3792.6]
  wire [7:0] _T_1331; // @[CSR.scala 278:45:@3799.8]
  wire [39:0] _T_1332; // @[Cat.scala 30:58:@3800.8]
  wire [40:0] _GEN_53; // @[CSR.scala 278:29:@3798.6]
  wire [31:0] _T_1334; // @[CSR.scala 277:72:@3805.8]
  wire [39:0] _T_1335; // @[Cat.scala 30:58:@3806.8]
  wire [40:0] _GEN_54; // @[CSR.scala 277:29:@3803.6]
  wire [7:0] _T_1336; // @[CSR.scala 278:45:@3810.8]
  wire [39:0] _T_1337; // @[Cat.scala 30:58:@3811.8]
  wire [40:0] _GEN_55; // @[CSR.scala 278:29:@3809.6]
  wire [31:0] _T_1339; // @[CSR.scala 277:72:@3816.8]
  wire [39:0] _T_1340; // @[Cat.scala 30:58:@3817.8]
  wire [40:0] _GEN_56; // @[CSR.scala 277:29:@3814.6]
  wire [7:0] _T_1341; // @[CSR.scala 278:45:@3821.8]
  wire [39:0] _T_1342; // @[Cat.scala 30:58:@3822.8]
  wire [40:0] _GEN_57; // @[CSR.scala 278:29:@3820.6]
  wire [31:0] _T_1344; // @[CSR.scala 277:72:@3827.8]
  wire [39:0] _T_1345; // @[Cat.scala 30:58:@3828.8]
  wire [40:0] _GEN_58; // @[CSR.scala 277:29:@3825.6]
  wire [7:0] _T_1346; // @[CSR.scala 278:45:@3832.8]
  wire [39:0] _T_1347; // @[Cat.scala 30:58:@3833.8]
  wire [40:0] _GEN_59; // @[CSR.scala 278:29:@3831.6]
  wire [31:0] _T_1349; // @[CSR.scala 277:72:@3838.8]
  wire [39:0] _T_1350; // @[Cat.scala 30:58:@3839.8]
  wire [40:0] _GEN_60; // @[CSR.scala 277:29:@3836.6]
  wire [7:0] _T_1351; // @[CSR.scala 278:45:@3843.8]
  wire [39:0] _T_1352; // @[Cat.scala 30:58:@3844.8]
  wire [40:0] _GEN_61; // @[CSR.scala 278:29:@3842.6]
  wire [31:0] _T_1354; // @[CSR.scala 277:72:@3849.8]
  wire [39:0] _T_1355; // @[Cat.scala 30:58:@3850.8]
  wire [40:0] _GEN_62; // @[CSR.scala 277:29:@3847.6]
  wire [7:0] _T_1356; // @[CSR.scala 278:45:@3854.8]
  wire [39:0] _T_1357; // @[Cat.scala 30:58:@3855.8]
  wire [40:0] _GEN_63; // @[CSR.scala 278:29:@3853.6]
  wire [31:0] _T_1359; // @[CSR.scala 277:72:@3860.8]
  wire [39:0] _T_1360; // @[Cat.scala 30:58:@3861.8]
  wire [40:0] _GEN_64; // @[CSR.scala 277:29:@3858.6]
  wire [7:0] _T_1361; // @[CSR.scala 278:45:@3865.8]
  wire [39:0] _T_1362; // @[Cat.scala 30:58:@3866.8]
  wire [40:0] _GEN_65; // @[CSR.scala 278:29:@3864.6]
  wire [31:0] _T_1364; // @[CSR.scala 277:72:@3871.8]
  wire [39:0] _T_1365; // @[Cat.scala 30:58:@3872.8]
  wire [40:0] _GEN_66; // @[CSR.scala 277:29:@3869.6]
  wire [7:0] _T_1366; // @[CSR.scala 278:45:@3876.8]
  wire [39:0] _T_1367; // @[Cat.scala 30:58:@3877.8]
  wire [40:0] _GEN_67; // @[CSR.scala 278:29:@3875.6]
  wire [31:0] _T_1369; // @[CSR.scala 277:72:@3882.8]
  wire [39:0] _T_1370; // @[Cat.scala 30:58:@3883.8]
  wire [40:0] _GEN_68; // @[CSR.scala 277:29:@3880.6]
  wire [7:0] _T_1371; // @[CSR.scala 278:45:@3887.8]
  wire [39:0] _T_1372; // @[Cat.scala 30:58:@3888.8]
  wire [40:0] _GEN_69; // @[CSR.scala 278:29:@3886.6]
  wire [31:0] _T_1374; // @[CSR.scala 277:72:@3893.8]
  wire [39:0] _T_1375; // @[Cat.scala 30:58:@3894.8]
  wire [40:0] _GEN_70; // @[CSR.scala 277:29:@3891.6]
  wire [7:0] _T_1376; // @[CSR.scala 278:45:@3898.8]
  wire [39:0] _T_1377; // @[Cat.scala 30:58:@3899.8]
  wire [40:0] _GEN_71; // @[CSR.scala 278:29:@3897.6]
  wire [31:0] _T_1379; // @[CSR.scala 277:72:@3904.8]
  wire [39:0] _T_1380; // @[Cat.scala 30:58:@3905.8]
  wire [40:0] _GEN_72; // @[CSR.scala 277:29:@3902.6]
  wire [7:0] _T_1381; // @[CSR.scala 278:45:@3909.8]
  wire [39:0] _T_1382; // @[Cat.scala 30:58:@3910.8]
  wire [40:0] _GEN_73; // @[CSR.scala 278:29:@3908.6]
  wire [31:0] _T_1384; // @[CSR.scala 277:72:@3915.8]
  wire [39:0] _T_1385; // @[Cat.scala 30:58:@3916.8]
  wire [40:0] _GEN_74; // @[CSR.scala 277:29:@3913.6]
  wire [7:0] _T_1386; // @[CSR.scala 278:45:@3920.8]
  wire [39:0] _T_1387; // @[Cat.scala 30:58:@3921.8]
  wire [40:0] _GEN_75; // @[CSR.scala 278:29:@3919.6]
  wire [31:0] _T_1389; // @[CSR.scala 277:72:@3926.8]
  wire [39:0] _T_1390; // @[Cat.scala 30:58:@3927.8]
  wire [40:0] _GEN_76; // @[CSR.scala 277:29:@3924.6]
  wire [7:0] _T_1391; // @[CSR.scala 278:45:@3931.8]
  wire [39:0] _T_1392; // @[Cat.scala 30:58:@3932.8]
  wire [40:0] _GEN_77; // @[CSR.scala 278:29:@3930.6]
  wire [31:0] _T_1394; // @[CSR.scala 277:72:@3937.8]
  wire [39:0] _T_1395; // @[Cat.scala 30:58:@3938.8]
  wire [40:0] _GEN_78; // @[CSR.scala 277:29:@3935.6]
  wire [7:0] _T_1396; // @[CSR.scala 278:45:@3942.8]
  wire [39:0] _T_1397; // @[Cat.scala 30:58:@3943.8]
  wire [40:0] _GEN_79; // @[CSR.scala 278:29:@3941.6]
  wire [31:0] _T_1399; // @[CSR.scala 277:72:@3948.8]
  wire [39:0] _T_1400; // @[Cat.scala 30:58:@3949.8]
  wire [40:0] _GEN_80; // @[CSR.scala 277:29:@3946.6]
  wire [7:0] _T_1401; // @[CSR.scala 278:45:@3953.8]
  wire [39:0] _T_1402; // @[Cat.scala 30:58:@3954.8]
  wire [40:0] _GEN_81; // @[CSR.scala 278:29:@3952.6]
  wire [31:0] _T_1404; // @[CSR.scala 277:72:@3959.8]
  wire [39:0] _T_1405; // @[Cat.scala 30:58:@3960.8]
  wire [40:0] _GEN_82; // @[CSR.scala 277:29:@3957.6]
  wire [7:0] _T_1406; // @[CSR.scala 278:45:@3964.8]
  wire [39:0] _T_1407; // @[Cat.scala 30:58:@3965.8]
  wire [40:0] _GEN_83; // @[CSR.scala 278:29:@3963.6]
  wire [31:0] _T_1409; // @[CSR.scala 277:72:@3970.8]
  wire [39:0] _T_1410; // @[Cat.scala 30:58:@3971.8]
  wire [40:0] _GEN_84; // @[CSR.scala 277:29:@3968.6]
  wire [7:0] _T_1411; // @[CSR.scala 278:45:@3975.8]
  wire [39:0] _T_1412; // @[Cat.scala 30:58:@3976.8]
  wire [40:0] _GEN_85; // @[CSR.scala 278:29:@3974.6]
  wire [31:0] _T_1414; // @[CSR.scala 277:72:@3981.8]
  wire [63:0] _T_1415; // @[Cat.scala 30:58:@3982.8]
  wire [57:0] _T_1416; // @[Util.scala 133:28:@3984.8]
  wire [63:0] _GEN_86; // @[CSR.scala 277:29:@3979.6]
  wire [57:0] _GEN_87; // @[CSR.scala 277:29:@3979.6]
  wire [31:0] _T_1417; // @[CSR.scala 278:45:@3988.8]
  wire [63:0] _T_1418; // @[Cat.scala 30:58:@3989.8]
  wire [57:0] _T_1419; // @[Util.scala 133:28:@3991.8]
  wire [63:0] _GEN_88; // @[CSR.scala 278:29:@3987.6]
  wire [57:0] _GEN_89; // @[CSR.scala 278:29:@3987.6]
  wire [31:0] _T_1421; // @[CSR.scala 277:72:@3996.8]
  wire [63:0] _T_1422; // @[Cat.scala 30:58:@3997.8]
  wire [57:0] _T_1423; // @[Util.scala 133:28:@3999.8]
  wire [63:0] _GEN_90; // @[CSR.scala 277:29:@3994.6]
  wire [57:0] _GEN_91; // @[CSR.scala 277:29:@3994.6]
  wire [31:0] _T_1424; // @[CSR.scala 278:45:@4003.8]
  wire [63:0] _T_1425; // @[Cat.scala 30:58:@4004.8]
  wire [57:0] _T_1426; // @[Util.scala 133:28:@4006.8]
  wire [63:0] _GEN_92; // @[CSR.scala 278:29:@4002.6]
  wire [57:0] _GEN_93; // @[CSR.scala 278:29:@4002.6]
  wire [31:0] _GEN_94; // @[CSR.scala 265:40:@4009.6]
  wire [31:0] _T_1429; // @[CSR.scala 267:78:@4014.8]
  wire [34:0] _GEN_225; // @[CSR.scala 267:86:@4015.8]
  wire [34:0] _T_1431; // @[CSR.scala 267:86:@4015.8]
  wire [34:0] _GEN_95; // @[CSR.scala 267:40:@4012.6]
  wire [31:0] _GEN_96; // @[CSR.scala 268:40:@4018.6]
  wire [31:0] _T_1433; // @[CSR.scala 269:62:@4022.8]
  wire [31:0] _GEN_97; // @[CSR.scala 269:40:@4021.6]
  wire [31:0] _GEN_98; // @[CSR.scala 270:40:@4025.6]
  wire [31:0] _GEN_99; // @[CSR.scala 271:42:@4029.6]
  wire  _GEN_100; // @[CSR.scala 242:14:@3558.4]
  wire  _GEN_101; // @[CSR.scala 242:14:@3558.4]
  wire  _GEN_102; // @[CSR.scala 242:14:@3558.4]
  wire  _GEN_103; // @[CSR.scala 242:14:@3558.4]
  wire  _GEN_104; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_105; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_106; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_107; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_108; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_109; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_110; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_111; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_112; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_113; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_114; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_115; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_116; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_117; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_118; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_119; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_120; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_121; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_122; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_123; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_124; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_125; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_126; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_127; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_128; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_129; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_130; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_131; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_132; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_133; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_134; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_135; // @[CSR.scala 242:14:@3558.4]
  wire [40:0] _GEN_136; // @[CSR.scala 242:14:@3558.4]
  wire [63:0] _GEN_137; // @[CSR.scala 242:14:@3558.4]
  wire [57:0] _GEN_138; // @[CSR.scala 242:14:@3558.4]
  wire [63:0] _GEN_139; // @[CSR.scala 242:14:@3558.4]
  wire [57:0] _GEN_140; // @[CSR.scala 242:14:@3558.4]
  wire [34:0] _GEN_142; // @[CSR.scala 242:14:@3558.4]
  assign _T_241 = _T_240 + 6'h1; // @[Util.scala 113:33:@2804.4]
  assign _T_245 = _T_241[6]; // @[Util.scala 118:20:@2807.4]
  assign _T_247 = _T_244 + 58'h1; // @[Util.scala 118:43:@2809.6]
  assign _T_248 = _T_244 + 58'h1; // @[Util.scala 118:43:@2810.6]
  assign _GEN_0 = _T_245 ? _T_248 : _T_244; // @[Util.scala 118:34:@2808.4]
  assign _T_249 = {_T_244,_T_240}; // @[Cat.scala 30:58:@2813.4]
  assign _GEN_147 = {{4'd0}, io_retire}; // @[Util.scala 113:33:@2815.4]
  assign _T_253 = _T_252 + _GEN_147; // @[Util.scala 113:33:@2815.4]
  assign _T_257 = _T_253[6]; // @[Util.scala 118:20:@2818.4]
  assign _T_259 = _T_256 + 58'h1; // @[Util.scala 118:43:@2820.6]
  assign _T_260 = _T_256 + 58'h1; // @[Util.scala 118:43:@2821.6]
  assign _GEN_1 = _T_257 ? _T_260 : _T_256; // @[Util.scala 118:34:@2819.4]
  assign _T_261 = {_T_256,_T_252}; // @[Cat.scala 30:58:@2824.4]
  assign _T_265 = {{1'd0}, _T_264}; // @[Util.scala 113:33:@2827.4]
  assign _T_268 = {{1'd0}, _T_267}; // @[Util.scala 113:33:@2830.4]
  assign _T_271 = {{1'd0}, _T_270}; // @[Util.scala 113:33:@2833.4]
  assign _T_274 = {{1'd0}, _T_273}; // @[Util.scala 113:33:@2836.4]
  assign _T_277 = {{1'd0}, _T_276}; // @[Util.scala 113:33:@2839.4]
  assign _T_280 = {{1'd0}, _T_279}; // @[Util.scala 113:33:@2842.4]
  assign _T_283 = {{1'd0}, _T_282}; // @[Util.scala 113:33:@2845.4]
  assign _T_286 = {{1'd0}, _T_285}; // @[Util.scala 113:33:@2848.4]
  assign _T_289 = {{1'd0}, _T_288}; // @[Util.scala 113:33:@2851.4]
  assign _T_292 = {{1'd0}, _T_291}; // @[Util.scala 113:33:@2854.4]
  assign _T_295 = {{1'd0}, _T_294}; // @[Util.scala 113:33:@2857.4]
  assign _T_298 = {{1'd0}, _T_297}; // @[Util.scala 113:33:@2860.4]
  assign _T_301 = {{1'd0}, _T_300}; // @[Util.scala 113:33:@2863.4]
  assign _T_304 = {{1'd0}, _T_303}; // @[Util.scala 113:33:@2866.4]
  assign _T_307 = {{1'd0}, _T_306}; // @[Util.scala 113:33:@2869.4]
  assign _T_310 = {{1'd0}, _T_309}; // @[Util.scala 113:33:@2872.4]
  assign _T_313 = {{1'd0}, _T_312}; // @[Util.scala 113:33:@2875.4]
  assign _T_316 = {{1'd0}, _T_315}; // @[Util.scala 113:33:@2878.4]
  assign _T_319 = {{1'd0}, _T_318}; // @[Util.scala 113:33:@2881.4]
  assign _T_322 = {{1'd0}, _T_321}; // @[Util.scala 113:33:@2884.4]
  assign _T_325 = {{1'd0}, _T_324}; // @[Util.scala 113:33:@2887.4]
  assign _T_328 = {{1'd0}, _T_327}; // @[Util.scala 113:33:@2890.4]
  assign _T_331 = {{1'd0}, _T_330}; // @[Util.scala 113:33:@2893.4]
  assign _T_334 = {{1'd0}, _T_333}; // @[Util.scala 113:33:@2896.4]
  assign _T_337 = {{1'd0}, _T_336}; // @[Util.scala 113:33:@2899.4]
  assign _T_340 = {{1'd0}, _T_339}; // @[Util.scala 113:33:@2902.4]
  assign _T_343 = {{1'd0}, _T_342}; // @[Util.scala 113:33:@2905.4]
  assign _T_346 = {{1'd0}, _T_345}; // @[Util.scala 113:33:@2908.4]
  assign _T_349 = {{1'd0}, _T_348}; // @[Util.scala 113:33:@2911.4]
  assign _T_352 = {{1'd0}, _T_351}; // @[Util.scala 113:33:@2914.4]
  assign _T_355 = {{1'd0}, _T_354}; // @[Util.scala 113:33:@2917.4]
  assign _T_358 = {{1'd0}, _T_357}; // @[Util.scala 113:33:@2920.4]
  assign system_insn = io_rw_cmd == 3'h4; // @[CSR.scala 137:31:@3011.4]
  assign _T_446 = io_rw_cmd != 3'h0; // @[CSR.scala 138:27:@3012.4]
  assign _T_448 = system_insn == 1'h0; // @[CSR.scala 138:40:@3013.4]
  assign cpu_ren = _T_446 & _T_448; // @[CSR.scala 138:37:@3014.4]
  assign read_mstatus = {io_status_prv,io_status_unimp5,io_status_mprv,io_status_unimp4,io_status_mpp,io_status_unimp3,io_status_mpie,io_status_unimp2,io_status_mie,io_status_unimp1}; // @[CSR.scala 140:32:@3023.4]
  assign _T_468 = {5'h0,3'h0,reg_mip_mtip,3'h0,reg_mip_msip,3'h0}; // @[CSR.scala 156:25:@3029.4]
  assign _T_474 = {5'h0,3'h0,reg_mie_mtip,3'h0,reg_mie_msip,3'h0}; // @[CSR.scala 157:25:@3035.4]
  assign _T_478 = io_rw_addr == 12'hb00; // @[CSR.scala 177:73:@3036.4]
  assign _T_480 = io_rw_addr == 12'hb02; // @[CSR.scala 177:73:@3037.4]
  assign _T_482 = io_rw_addr == 12'hf13; // @[CSR.scala 177:73:@3038.4]
  assign _T_488 = io_rw_addr == 12'h301; // @[CSR.scala 177:73:@3041.4]
  assign _T_490 = io_rw_addr == 12'h300; // @[CSR.scala 177:73:@3042.4]
  assign _T_492 = io_rw_addr == 12'h305; // @[CSR.scala 177:73:@3043.4]
  assign _T_494 = io_rw_addr == 12'h344; // @[CSR.scala 177:73:@3044.4]
  assign _T_496 = io_rw_addr == 12'h304; // @[CSR.scala 177:73:@3045.4]
  assign _T_498 = io_rw_addr == 12'h340; // @[CSR.scala 177:73:@3046.4]
  assign _T_500 = io_rw_addr == 12'h341; // @[CSR.scala 177:73:@3047.4]
  assign _T_502 = io_rw_addr == 12'h343; // @[CSR.scala 177:73:@3048.4]
  assign _T_504 = io_rw_addr == 12'h342; // @[CSR.scala 177:73:@3049.4]
  assign _T_508 = io_rw_addr == 12'h7b2; // @[CSR.scala 177:73:@3051.4]
  assign _T_510 = io_rw_addr == 12'h302; // @[CSR.scala 177:73:@3052.4]
  assign _T_512 = io_rw_addr == 12'hb03; // @[CSR.scala 177:73:@3053.4]
  assign _T_514 = io_rw_addr == 12'hb83; // @[CSR.scala 177:73:@3054.4]
  assign _T_516 = io_rw_addr == 12'hb04; // @[CSR.scala 177:73:@3055.4]
  assign _T_518 = io_rw_addr == 12'hb84; // @[CSR.scala 177:73:@3056.4]
  assign _T_520 = io_rw_addr == 12'hb05; // @[CSR.scala 177:73:@3057.4]
  assign _T_522 = io_rw_addr == 12'hb85; // @[CSR.scala 177:73:@3058.4]
  assign _T_524 = io_rw_addr == 12'hb06; // @[CSR.scala 177:73:@3059.4]
  assign _T_526 = io_rw_addr == 12'hb86; // @[CSR.scala 177:73:@3060.4]
  assign _T_528 = io_rw_addr == 12'hb07; // @[CSR.scala 177:73:@3061.4]
  assign _T_530 = io_rw_addr == 12'hb87; // @[CSR.scala 177:73:@3062.4]
  assign _T_532 = io_rw_addr == 12'hb08; // @[CSR.scala 177:73:@3063.4]
  assign _T_534 = io_rw_addr == 12'hb88; // @[CSR.scala 177:73:@3064.4]
  assign _T_536 = io_rw_addr == 12'hb09; // @[CSR.scala 177:73:@3065.4]
  assign _T_538 = io_rw_addr == 12'hb89; // @[CSR.scala 177:73:@3066.4]
  assign _T_540 = io_rw_addr == 12'hb0a; // @[CSR.scala 177:73:@3067.4]
  assign _T_542 = io_rw_addr == 12'hb8a; // @[CSR.scala 177:73:@3068.4]
  assign _T_544 = io_rw_addr == 12'hb0b; // @[CSR.scala 177:73:@3069.4]
  assign _T_546 = io_rw_addr == 12'hb8b; // @[CSR.scala 177:73:@3070.4]
  assign _T_548 = io_rw_addr == 12'hb0c; // @[CSR.scala 177:73:@3071.4]
  assign _T_550 = io_rw_addr == 12'hb8c; // @[CSR.scala 177:73:@3072.4]
  assign _T_552 = io_rw_addr == 12'hb0d; // @[CSR.scala 177:73:@3073.4]
  assign _T_554 = io_rw_addr == 12'hb8d; // @[CSR.scala 177:73:@3074.4]
  assign _T_556 = io_rw_addr == 12'hb0e; // @[CSR.scala 177:73:@3075.4]
  assign _T_558 = io_rw_addr == 12'hb8e; // @[CSR.scala 177:73:@3076.4]
  assign _T_560 = io_rw_addr == 12'hb0f; // @[CSR.scala 177:73:@3077.4]
  assign _T_562 = io_rw_addr == 12'hb8f; // @[CSR.scala 177:73:@3078.4]
  assign _T_564 = io_rw_addr == 12'hb10; // @[CSR.scala 177:73:@3079.4]
  assign _T_566 = io_rw_addr == 12'hb90; // @[CSR.scala 177:73:@3080.4]
  assign _T_568 = io_rw_addr == 12'hb11; // @[CSR.scala 177:73:@3081.4]
  assign _T_570 = io_rw_addr == 12'hb91; // @[CSR.scala 177:73:@3082.4]
  assign _T_572 = io_rw_addr == 12'hb12; // @[CSR.scala 177:73:@3083.4]
  assign _T_574 = io_rw_addr == 12'hb92; // @[CSR.scala 177:73:@3084.4]
  assign _T_576 = io_rw_addr == 12'hb13; // @[CSR.scala 177:73:@3085.4]
  assign _T_578 = io_rw_addr == 12'hb93; // @[CSR.scala 177:73:@3086.4]
  assign _T_580 = io_rw_addr == 12'hb14; // @[CSR.scala 177:73:@3087.4]
  assign _T_582 = io_rw_addr == 12'hb94; // @[CSR.scala 177:73:@3088.4]
  assign _T_584 = io_rw_addr == 12'hb15; // @[CSR.scala 177:73:@3089.4]
  assign _T_586 = io_rw_addr == 12'hb95; // @[CSR.scala 177:73:@3090.4]
  assign _T_588 = io_rw_addr == 12'hb16; // @[CSR.scala 177:73:@3091.4]
  assign _T_590 = io_rw_addr == 12'hb96; // @[CSR.scala 177:73:@3092.4]
  assign _T_592 = io_rw_addr == 12'hb17; // @[CSR.scala 177:73:@3093.4]
  assign _T_594 = io_rw_addr == 12'hb97; // @[CSR.scala 177:73:@3094.4]
  assign _T_596 = io_rw_addr == 12'hb18; // @[CSR.scala 177:73:@3095.4]
  assign _T_598 = io_rw_addr == 12'hb98; // @[CSR.scala 177:73:@3096.4]
  assign _T_600 = io_rw_addr == 12'hb19; // @[CSR.scala 177:73:@3097.4]
  assign _T_602 = io_rw_addr == 12'hb99; // @[CSR.scala 177:73:@3098.4]
  assign _T_604 = io_rw_addr == 12'hb1a; // @[CSR.scala 177:73:@3099.4]
  assign _T_606 = io_rw_addr == 12'hb9a; // @[CSR.scala 177:73:@3100.4]
  assign _T_608 = io_rw_addr == 12'hb1b; // @[CSR.scala 177:73:@3101.4]
  assign _T_610 = io_rw_addr == 12'hb9b; // @[CSR.scala 177:73:@3102.4]
  assign _T_612 = io_rw_addr == 12'hb1c; // @[CSR.scala 177:73:@3103.4]
  assign _T_614 = io_rw_addr == 12'hb9c; // @[CSR.scala 177:73:@3104.4]
  assign _T_616 = io_rw_addr == 12'hb1d; // @[CSR.scala 177:73:@3105.4]
  assign _T_618 = io_rw_addr == 12'hb9d; // @[CSR.scala 177:73:@3106.4]
  assign _T_620 = io_rw_addr == 12'hb1e; // @[CSR.scala 177:73:@3107.4]
  assign _T_622 = io_rw_addr == 12'hb9e; // @[CSR.scala 177:73:@3108.4]
  assign _T_624 = io_rw_addr == 12'hb1f; // @[CSR.scala 177:73:@3109.4]
  assign _T_626 = io_rw_addr == 12'hb9f; // @[CSR.scala 177:73:@3110.4]
  assign _T_628 = io_rw_addr == 12'hb20; // @[CSR.scala 177:73:@3111.4]
  assign _T_630 = io_rw_addr == 12'hba0; // @[CSR.scala 177:73:@3112.4]
  assign _T_632 = io_rw_addr == 12'hb21; // @[CSR.scala 177:73:@3113.4]
  assign _T_634 = io_rw_addr == 12'hba1; // @[CSR.scala 177:73:@3114.4]
  assign _T_636 = io_rw_addr == 12'hb22; // @[CSR.scala 177:73:@3115.4]
  assign _T_638 = io_rw_addr == 12'hba2; // @[CSR.scala 177:73:@3116.4]
  assign _T_640 = io_rw_addr == 12'hb80; // @[CSR.scala 177:73:@3117.4]
  assign _T_642 = io_rw_addr == 12'hb82; // @[CSR.scala 177:73:@3118.4]
  assign _T_643 = io_rw_addr[9:8]; // @[CSR.scala 179:54:@3119.4]
  assign priv_sufficient = reg_mstatus_prv >= _T_643; // @[CSR.scala 179:41:@3120.4]
  assign _T_644 = io_rw_addr[11:10]; // @[CSR.scala 180:29:@3121.4]
  assign _T_645 = ~ _T_644; // @[CSR.scala 180:37:@3122.4]
  assign read_only = _T_645 == 2'h0; // @[CSR.scala 180:37:@3123.4]
  assign _T_647 = io_rw_cmd != 3'h5; // @[CSR.scala 181:38:@3124.4]
  assign _T_648 = cpu_ren & _T_647; // @[CSR.scala 181:25:@3125.4]
  assign cpu_wen = _T_648 & priv_sufficient; // @[CSR.scala 181:48:@3126.4]
  assign _T_650 = read_only == 1'h0; // @[CSR.scala 182:24:@3127.4]
  assign wen = cpu_wen & _T_650; // @[CSR.scala 182:21:@3128.4]
  assign _T_651 = io_rw_cmd == 3'h2; // @[Util.scala 23:47:@3129.4]
  assign _T_652 = io_rw_cmd == 3'h3; // @[Util.scala 23:47:@3130.4]
  assign _T_653 = _T_651 | _T_652; // @[Util.scala 23:62:@3131.4]
  assign _T_655 = _T_653 ? io_rw_rdata : 32'h0; // @[CSR.scala 281:9:@3132.4]
  assign _T_656 = _T_655 | io_rw_wdata; // @[CSR.scala 281:49:@3133.4]
  assign _T_659 = _T_652 ? io_rw_wdata : 32'h0; // @[CSR.scala 281:64:@3135.4]
  assign _T_660 = ~ _T_659; // @[CSR.scala 281:60:@3136.4]
  assign wdata = _T_656 & _T_660; // @[CSR.scala 281:58:@3137.4]
  assign _T_662 = io_rw_addr[2:0]; // @[CSR.scala 185:33:@3138.4]
  assign opcode = 8'h1 << _T_662; // @[CSR.scala 185:20:@3139.4]
  assign _T_663 = opcode[0]; // @[CSR.scala 186:40:@3140.4]
  assign insn_call = system_insn & _T_663; // @[CSR.scala 186:31:@3141.4]
  assign _T_664 = opcode[1]; // @[CSR.scala 187:41:@3142.4]
  assign insn_break = system_insn & _T_664; // @[CSR.scala 187:32:@3143.4]
  assign _T_665 = opcode[2]; // @[CSR.scala 188:39:@3144.4]
  assign _T_666 = system_insn & _T_665; // @[CSR.scala 188:30:@3145.4]
  assign insn_ret = _T_666 & priv_sufficient; // @[CSR.scala 188:43:@3146.4]
  assign _T_940 = insn_call | insn_break; // @[CSR.scala 199:24:@3345.4]
  assign _T_942 = {{1'd0}, insn_ret}; // @[Bitwise.scala 48:55:@3348.4]
  assign _T_944 = _T_942 <= 2'h1; // @[CSR.scala 201:50:@3349.4]
  assign _T_946 = _T_944 | reset; // @[CSR.scala 201:9:@3351.4]
  assign _T_948 = _T_946 == 1'h0; // @[CSR.scala 201:9:@3352.4]
  assign _T_951 = io_rw_addr[10]; // @[CSR.scala 208:32:@3361.4]
  assign _T_953 = _T_951 == 1'h0; // @[CSR.scala 208:21:@3362.4]
  assign _T_954 = insn_ret & _T_953; // @[CSR.scala 208:18:@3363.4]
  assign _GEN_3 = _T_954 ? reg_mstatus_mpie : reg_mstatus_mie; // @[CSR.scala 208:38:@3364.4]
  assign _GEN_4 = _T_954 ? 1'h1 : reg_mstatus_mpie; // @[CSR.scala 208:38:@3364.4]
  assign new_prv = _T_954 ? 2'h3 : reg_mstatus_prv; // @[CSR.scala 208:38:@3364.4]
  assign _GEN_148 = {{2'd0}, reg_mstatus_prv}; // @[CSR.scala 218:35:@3372.6]
  assign _T_958 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3372.6]
  assign _T_959 = _GEN_148 + 4'h8; // @[CSR.scala 218:35:@3373.6]
  assign _GEN_7 = insn_call ? 32'h80000004 : reg_mepc; // @[CSR.scala 216:18:@3370.4]
  assign _GEN_8 = insn_call ? {{28'd0}, _T_959} : reg_mcause; // @[CSR.scala 216:18:@3370.4]
  assign _GEN_9 = insn_call ? io_pc : reg_mepc; // @[CSR.scala 216:18:@3370.4]
  assign _GEN_10 = insn_break ? 32'h80000004 : _GEN_7; // @[CSR.scala 223:19:@3377.4]
  assign _GEN_11 = insn_break ? 32'h3 : _GEN_8; // @[CSR.scala 223:19:@3377.4]
  assign _GEN_12 = insn_break ? io_pc : _GEN_9; // @[CSR.scala 223:19:@3377.4]
  assign _GEN_14 = io_xcpt ? io_cause : _GEN_11; // @[CSR.scala 229:17:@3382.4]
  assign _GEN_15 = io_xcpt ? io_pc : _GEN_12; // @[CSR.scala 229:17:@3382.4]
  assign _GEN_16 = io_xcpt ? io_tval : reg_mtval; // @[CSR.scala 229:17:@3382.4]
  assign _T_965 = _T_478 ? _T_249 : 64'h0; // @[Mux.scala 19:72:@3390.4]
  assign _T_967 = _T_480 ? _T_261 : 64'h0; // @[Mux.scala 19:72:@3391.4]
  assign _T_969 = _T_482 ? 16'h8000 : 16'h0; // @[Mux.scala 19:72:@3392.4]
  assign _T_975 = _T_488 ? 31'h40000100 : 31'h0; // @[Mux.scala 19:72:@3395.4]
  assign _T_977 = _T_490 ? read_mstatus : 32'h0; // @[Mux.scala 19:72:@3396.4]
  assign _T_979 = _T_492 ? 9'h100 : 9'h0; // @[Mux.scala 19:72:@3397.4]
  assign _T_981 = _T_494 ? _T_468 : 16'h0; // @[Mux.scala 19:72:@3398.4]
  assign _T_983 = _T_496 ? _T_474 : 16'h0; // @[Mux.scala 19:72:@3399.4]
  assign _T_985 = _T_498 ? reg_mscratch : 32'h0; // @[Mux.scala 19:72:@3400.4]
  assign _T_987 = _T_500 ? reg_mepc : 32'h0; // @[Mux.scala 19:72:@3401.4]
  assign _T_989 = _T_502 ? reg_mtval : 32'h0; // @[Mux.scala 19:72:@3402.4]
  assign _T_991 = _T_504 ? reg_mcause : 32'h0; // @[Mux.scala 19:72:@3403.4]
  assign _T_995 = _T_508 ? reg_dscratch : 32'h0; // @[Mux.scala 19:72:@3405.4]
  assign _T_997 = _T_510 ? reg_medeleg : 32'h0; // @[Mux.scala 19:72:@3406.4]
  assign _T_999 = _T_512 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3407.4]
  assign _T_1001 = _T_514 ? _T_264 : 40'h0; // @[Mux.scala 19:72:@3408.4]
  assign _T_1003 = _T_516 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3409.4]
  assign _T_1005 = _T_518 ? _T_267 : 40'h0; // @[Mux.scala 19:72:@3410.4]
  assign _T_1007 = _T_520 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3411.4]
  assign _T_1009 = _T_522 ? _T_270 : 40'h0; // @[Mux.scala 19:72:@3412.4]
  assign _T_1011 = _T_524 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3413.4]
  assign _T_1013 = _T_526 ? _T_273 : 40'h0; // @[Mux.scala 19:72:@3414.4]
  assign _T_1015 = _T_528 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3415.4]
  assign _T_1017 = _T_530 ? _T_276 : 40'h0; // @[Mux.scala 19:72:@3416.4]
  assign _T_1019 = _T_532 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3417.4]
  assign _T_1021 = _T_534 ? _T_279 : 40'h0; // @[Mux.scala 19:72:@3418.4]
  assign _T_1023 = _T_536 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3419.4]
  assign _T_1025 = _T_538 ? _T_282 : 40'h0; // @[Mux.scala 19:72:@3420.4]
  assign _T_1027 = _T_540 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3421.4]
  assign _T_1029 = _T_542 ? _T_285 : 40'h0; // @[Mux.scala 19:72:@3422.4]
  assign _T_1031 = _T_544 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3423.4]
  assign _T_1033 = _T_546 ? _T_288 : 40'h0; // @[Mux.scala 19:72:@3424.4]
  assign _T_1035 = _T_548 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3425.4]
  assign _T_1037 = _T_550 ? _T_291 : 40'h0; // @[Mux.scala 19:72:@3426.4]
  assign _T_1039 = _T_552 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3427.4]
  assign _T_1041 = _T_554 ? _T_294 : 40'h0; // @[Mux.scala 19:72:@3428.4]
  assign _T_1043 = _T_556 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3429.4]
  assign _T_1045 = _T_558 ? _T_297 : 40'h0; // @[Mux.scala 19:72:@3430.4]
  assign _T_1047 = _T_560 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3431.4]
  assign _T_1049 = _T_562 ? _T_300 : 40'h0; // @[Mux.scala 19:72:@3432.4]
  assign _T_1051 = _T_564 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3433.4]
  assign _T_1053 = _T_566 ? _T_303 : 40'h0; // @[Mux.scala 19:72:@3434.4]
  assign _T_1055 = _T_568 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3435.4]
  assign _T_1057 = _T_570 ? _T_306 : 40'h0; // @[Mux.scala 19:72:@3436.4]
  assign _T_1059 = _T_572 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3437.4]
  assign _T_1061 = _T_574 ? _T_309 : 40'h0; // @[Mux.scala 19:72:@3438.4]
  assign _T_1063 = _T_576 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3439.4]
  assign _T_1065 = _T_578 ? _T_312 : 40'h0; // @[Mux.scala 19:72:@3440.4]
  assign _T_1067 = _T_580 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3441.4]
  assign _T_1069 = _T_582 ? _T_315 : 40'h0; // @[Mux.scala 19:72:@3442.4]
  assign _T_1071 = _T_584 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3443.4]
  assign _T_1073 = _T_586 ? _T_318 : 40'h0; // @[Mux.scala 19:72:@3444.4]
  assign _T_1075 = _T_588 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3445.4]
  assign _T_1077 = _T_590 ? _T_321 : 40'h0; // @[Mux.scala 19:72:@3446.4]
  assign _T_1079 = _T_592 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3447.4]
  assign _T_1081 = _T_594 ? _T_324 : 40'h0; // @[Mux.scala 19:72:@3448.4]
  assign _T_1083 = _T_596 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3449.4]
  assign _T_1085 = _T_598 ? _T_327 : 40'h0; // @[Mux.scala 19:72:@3450.4]
  assign _T_1087 = _T_600 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3451.4]
  assign _T_1089 = _T_602 ? _T_330 : 40'h0; // @[Mux.scala 19:72:@3452.4]
  assign _T_1091 = _T_604 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3453.4]
  assign _T_1093 = _T_606 ? _T_333 : 40'h0; // @[Mux.scala 19:72:@3454.4]
  assign _T_1095 = _T_608 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3455.4]
  assign _T_1097 = _T_610 ? _T_336 : 40'h0; // @[Mux.scala 19:72:@3456.4]
  assign _T_1099 = _T_612 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3457.4]
  assign _T_1101 = _T_614 ? _T_339 : 40'h0; // @[Mux.scala 19:72:@3458.4]
  assign _T_1103 = _T_616 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3459.4]
  assign _T_1105 = _T_618 ? _T_342 : 40'h0; // @[Mux.scala 19:72:@3460.4]
  assign _T_1107 = _T_620 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3461.4]
  assign _T_1109 = _T_622 ? _T_345 : 40'h0; // @[Mux.scala 19:72:@3462.4]
  assign _T_1111 = _T_624 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3463.4]
  assign _T_1113 = _T_626 ? _T_348 : 40'h0; // @[Mux.scala 19:72:@3464.4]
  assign _T_1115 = _T_628 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@3465.4]
  assign _T_1117 = _T_630 ? _T_351 : 40'h0; // @[Mux.scala 19:72:@3466.4]
  assign _T_1119 = _T_632 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@3467.4]
  assign _T_1121 = _T_634 ? _T_354 : 40'h0; // @[Mux.scala 19:72:@3468.4]
  assign _T_1123 = _T_636 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@3469.4]
  assign _T_1125 = _T_638 ? _T_357 : 40'h0; // @[Mux.scala 19:72:@3470.4]
  assign _T_1130 = _T_965 | _T_967; // @[Mux.scala 19:72:@3473.4]
  assign _GEN_149 = {{48'd0}, _T_969}; // @[Mux.scala 19:72:@3474.4]
  assign _T_1131 = _T_1130 | _GEN_149; // @[Mux.scala 19:72:@3474.4]
  assign _GEN_150 = {{33'd0}, _T_975}; // @[Mux.scala 19:72:@3477.4]
  assign _T_1134 = _T_1131 | _GEN_150; // @[Mux.scala 19:72:@3477.4]
  assign _GEN_151 = {{32'd0}, _T_977}; // @[Mux.scala 19:72:@3478.4]
  assign _T_1135 = _T_1134 | _GEN_151; // @[Mux.scala 19:72:@3478.4]
  assign _GEN_152 = {{55'd0}, _T_979}; // @[Mux.scala 19:72:@3479.4]
  assign _T_1136 = _T_1135 | _GEN_152; // @[Mux.scala 19:72:@3479.4]
  assign _GEN_153 = {{48'd0}, _T_981}; // @[Mux.scala 19:72:@3480.4]
  assign _T_1137 = _T_1136 | _GEN_153; // @[Mux.scala 19:72:@3480.4]
  assign _GEN_154 = {{48'd0}, _T_983}; // @[Mux.scala 19:72:@3481.4]
  assign _T_1138 = _T_1137 | _GEN_154; // @[Mux.scala 19:72:@3481.4]
  assign _GEN_155 = {{32'd0}, _T_985}; // @[Mux.scala 19:72:@3482.4]
  assign _T_1139 = _T_1138 | _GEN_155; // @[Mux.scala 19:72:@3482.4]
  assign _GEN_156 = {{32'd0}, _T_987}; // @[Mux.scala 19:72:@3483.4]
  assign _T_1140 = _T_1139 | _GEN_156; // @[Mux.scala 19:72:@3483.4]
  assign _GEN_157 = {{32'd0}, _T_989}; // @[Mux.scala 19:72:@3484.4]
  assign _T_1141 = _T_1140 | _GEN_157; // @[Mux.scala 19:72:@3484.4]
  assign _GEN_158 = {{32'd0}, _T_991}; // @[Mux.scala 19:72:@3485.4]
  assign _T_1142 = _T_1141 | _GEN_158; // @[Mux.scala 19:72:@3485.4]
  assign _GEN_159 = {{32'd0}, _T_995}; // @[Mux.scala 19:72:@3487.4]
  assign _T_1144 = _T_1142 | _GEN_159; // @[Mux.scala 19:72:@3487.4]
  assign _GEN_160 = {{32'd0}, _T_997}; // @[Mux.scala 19:72:@3488.4]
  assign _T_1145 = _T_1144 | _GEN_160; // @[Mux.scala 19:72:@3488.4]
  assign _GEN_161 = {{24'd0}, _T_999}; // @[Mux.scala 19:72:@3489.4]
  assign _T_1146 = _T_1145 | _GEN_161; // @[Mux.scala 19:72:@3489.4]
  assign _GEN_162 = {{24'd0}, _T_1001}; // @[Mux.scala 19:72:@3490.4]
  assign _T_1147 = _T_1146 | _GEN_162; // @[Mux.scala 19:72:@3490.4]
  assign _GEN_163 = {{24'd0}, _T_1003}; // @[Mux.scala 19:72:@3491.4]
  assign _T_1148 = _T_1147 | _GEN_163; // @[Mux.scala 19:72:@3491.4]
  assign _GEN_164 = {{24'd0}, _T_1005}; // @[Mux.scala 19:72:@3492.4]
  assign _T_1149 = _T_1148 | _GEN_164; // @[Mux.scala 19:72:@3492.4]
  assign _GEN_165 = {{24'd0}, _T_1007}; // @[Mux.scala 19:72:@3493.4]
  assign _T_1150 = _T_1149 | _GEN_165; // @[Mux.scala 19:72:@3493.4]
  assign _GEN_166 = {{24'd0}, _T_1009}; // @[Mux.scala 19:72:@3494.4]
  assign _T_1151 = _T_1150 | _GEN_166; // @[Mux.scala 19:72:@3494.4]
  assign _GEN_167 = {{24'd0}, _T_1011}; // @[Mux.scala 19:72:@3495.4]
  assign _T_1152 = _T_1151 | _GEN_167; // @[Mux.scala 19:72:@3495.4]
  assign _GEN_168 = {{24'd0}, _T_1013}; // @[Mux.scala 19:72:@3496.4]
  assign _T_1153 = _T_1152 | _GEN_168; // @[Mux.scala 19:72:@3496.4]
  assign _GEN_169 = {{24'd0}, _T_1015}; // @[Mux.scala 19:72:@3497.4]
  assign _T_1154 = _T_1153 | _GEN_169; // @[Mux.scala 19:72:@3497.4]
  assign _GEN_170 = {{24'd0}, _T_1017}; // @[Mux.scala 19:72:@3498.4]
  assign _T_1155 = _T_1154 | _GEN_170; // @[Mux.scala 19:72:@3498.4]
  assign _GEN_171 = {{24'd0}, _T_1019}; // @[Mux.scala 19:72:@3499.4]
  assign _T_1156 = _T_1155 | _GEN_171; // @[Mux.scala 19:72:@3499.4]
  assign _GEN_172 = {{24'd0}, _T_1021}; // @[Mux.scala 19:72:@3500.4]
  assign _T_1157 = _T_1156 | _GEN_172; // @[Mux.scala 19:72:@3500.4]
  assign _GEN_173 = {{24'd0}, _T_1023}; // @[Mux.scala 19:72:@3501.4]
  assign _T_1158 = _T_1157 | _GEN_173; // @[Mux.scala 19:72:@3501.4]
  assign _GEN_174 = {{24'd0}, _T_1025}; // @[Mux.scala 19:72:@3502.4]
  assign _T_1159 = _T_1158 | _GEN_174; // @[Mux.scala 19:72:@3502.4]
  assign _GEN_175 = {{24'd0}, _T_1027}; // @[Mux.scala 19:72:@3503.4]
  assign _T_1160 = _T_1159 | _GEN_175; // @[Mux.scala 19:72:@3503.4]
  assign _GEN_176 = {{24'd0}, _T_1029}; // @[Mux.scala 19:72:@3504.4]
  assign _T_1161 = _T_1160 | _GEN_176; // @[Mux.scala 19:72:@3504.4]
  assign _GEN_177 = {{24'd0}, _T_1031}; // @[Mux.scala 19:72:@3505.4]
  assign _T_1162 = _T_1161 | _GEN_177; // @[Mux.scala 19:72:@3505.4]
  assign _GEN_178 = {{24'd0}, _T_1033}; // @[Mux.scala 19:72:@3506.4]
  assign _T_1163 = _T_1162 | _GEN_178; // @[Mux.scala 19:72:@3506.4]
  assign _GEN_179 = {{24'd0}, _T_1035}; // @[Mux.scala 19:72:@3507.4]
  assign _T_1164 = _T_1163 | _GEN_179; // @[Mux.scala 19:72:@3507.4]
  assign _GEN_180 = {{24'd0}, _T_1037}; // @[Mux.scala 19:72:@3508.4]
  assign _T_1165 = _T_1164 | _GEN_180; // @[Mux.scala 19:72:@3508.4]
  assign _GEN_181 = {{24'd0}, _T_1039}; // @[Mux.scala 19:72:@3509.4]
  assign _T_1166 = _T_1165 | _GEN_181; // @[Mux.scala 19:72:@3509.4]
  assign _GEN_182 = {{24'd0}, _T_1041}; // @[Mux.scala 19:72:@3510.4]
  assign _T_1167 = _T_1166 | _GEN_182; // @[Mux.scala 19:72:@3510.4]
  assign _GEN_183 = {{24'd0}, _T_1043}; // @[Mux.scala 19:72:@3511.4]
  assign _T_1168 = _T_1167 | _GEN_183; // @[Mux.scala 19:72:@3511.4]
  assign _GEN_184 = {{24'd0}, _T_1045}; // @[Mux.scala 19:72:@3512.4]
  assign _T_1169 = _T_1168 | _GEN_184; // @[Mux.scala 19:72:@3512.4]
  assign _GEN_185 = {{24'd0}, _T_1047}; // @[Mux.scala 19:72:@3513.4]
  assign _T_1170 = _T_1169 | _GEN_185; // @[Mux.scala 19:72:@3513.4]
  assign _GEN_186 = {{24'd0}, _T_1049}; // @[Mux.scala 19:72:@3514.4]
  assign _T_1171 = _T_1170 | _GEN_186; // @[Mux.scala 19:72:@3514.4]
  assign _GEN_187 = {{24'd0}, _T_1051}; // @[Mux.scala 19:72:@3515.4]
  assign _T_1172 = _T_1171 | _GEN_187; // @[Mux.scala 19:72:@3515.4]
  assign _GEN_188 = {{24'd0}, _T_1053}; // @[Mux.scala 19:72:@3516.4]
  assign _T_1173 = _T_1172 | _GEN_188; // @[Mux.scala 19:72:@3516.4]
  assign _GEN_189 = {{24'd0}, _T_1055}; // @[Mux.scala 19:72:@3517.4]
  assign _T_1174 = _T_1173 | _GEN_189; // @[Mux.scala 19:72:@3517.4]
  assign _GEN_190 = {{24'd0}, _T_1057}; // @[Mux.scala 19:72:@3518.4]
  assign _T_1175 = _T_1174 | _GEN_190; // @[Mux.scala 19:72:@3518.4]
  assign _GEN_191 = {{24'd0}, _T_1059}; // @[Mux.scala 19:72:@3519.4]
  assign _T_1176 = _T_1175 | _GEN_191; // @[Mux.scala 19:72:@3519.4]
  assign _GEN_192 = {{24'd0}, _T_1061}; // @[Mux.scala 19:72:@3520.4]
  assign _T_1177 = _T_1176 | _GEN_192; // @[Mux.scala 19:72:@3520.4]
  assign _GEN_193 = {{24'd0}, _T_1063}; // @[Mux.scala 19:72:@3521.4]
  assign _T_1178 = _T_1177 | _GEN_193; // @[Mux.scala 19:72:@3521.4]
  assign _GEN_194 = {{24'd0}, _T_1065}; // @[Mux.scala 19:72:@3522.4]
  assign _T_1179 = _T_1178 | _GEN_194; // @[Mux.scala 19:72:@3522.4]
  assign _GEN_195 = {{24'd0}, _T_1067}; // @[Mux.scala 19:72:@3523.4]
  assign _T_1180 = _T_1179 | _GEN_195; // @[Mux.scala 19:72:@3523.4]
  assign _GEN_196 = {{24'd0}, _T_1069}; // @[Mux.scala 19:72:@3524.4]
  assign _T_1181 = _T_1180 | _GEN_196; // @[Mux.scala 19:72:@3524.4]
  assign _GEN_197 = {{24'd0}, _T_1071}; // @[Mux.scala 19:72:@3525.4]
  assign _T_1182 = _T_1181 | _GEN_197; // @[Mux.scala 19:72:@3525.4]
  assign _GEN_198 = {{24'd0}, _T_1073}; // @[Mux.scala 19:72:@3526.4]
  assign _T_1183 = _T_1182 | _GEN_198; // @[Mux.scala 19:72:@3526.4]
  assign _GEN_199 = {{24'd0}, _T_1075}; // @[Mux.scala 19:72:@3527.4]
  assign _T_1184 = _T_1183 | _GEN_199; // @[Mux.scala 19:72:@3527.4]
  assign _GEN_200 = {{24'd0}, _T_1077}; // @[Mux.scala 19:72:@3528.4]
  assign _T_1185 = _T_1184 | _GEN_200; // @[Mux.scala 19:72:@3528.4]
  assign _GEN_201 = {{24'd0}, _T_1079}; // @[Mux.scala 19:72:@3529.4]
  assign _T_1186 = _T_1185 | _GEN_201; // @[Mux.scala 19:72:@3529.4]
  assign _GEN_202 = {{24'd0}, _T_1081}; // @[Mux.scala 19:72:@3530.4]
  assign _T_1187 = _T_1186 | _GEN_202; // @[Mux.scala 19:72:@3530.4]
  assign _GEN_203 = {{24'd0}, _T_1083}; // @[Mux.scala 19:72:@3531.4]
  assign _T_1188 = _T_1187 | _GEN_203; // @[Mux.scala 19:72:@3531.4]
  assign _GEN_204 = {{24'd0}, _T_1085}; // @[Mux.scala 19:72:@3532.4]
  assign _T_1189 = _T_1188 | _GEN_204; // @[Mux.scala 19:72:@3532.4]
  assign _GEN_205 = {{24'd0}, _T_1087}; // @[Mux.scala 19:72:@3533.4]
  assign _T_1190 = _T_1189 | _GEN_205; // @[Mux.scala 19:72:@3533.4]
  assign _GEN_206 = {{24'd0}, _T_1089}; // @[Mux.scala 19:72:@3534.4]
  assign _T_1191 = _T_1190 | _GEN_206; // @[Mux.scala 19:72:@3534.4]
  assign _GEN_207 = {{24'd0}, _T_1091}; // @[Mux.scala 19:72:@3535.4]
  assign _T_1192 = _T_1191 | _GEN_207; // @[Mux.scala 19:72:@3535.4]
  assign _GEN_208 = {{24'd0}, _T_1093}; // @[Mux.scala 19:72:@3536.4]
  assign _T_1193 = _T_1192 | _GEN_208; // @[Mux.scala 19:72:@3536.4]
  assign _GEN_209 = {{24'd0}, _T_1095}; // @[Mux.scala 19:72:@3537.4]
  assign _T_1194 = _T_1193 | _GEN_209; // @[Mux.scala 19:72:@3537.4]
  assign _GEN_210 = {{24'd0}, _T_1097}; // @[Mux.scala 19:72:@3538.4]
  assign _T_1195 = _T_1194 | _GEN_210; // @[Mux.scala 19:72:@3538.4]
  assign _GEN_211 = {{24'd0}, _T_1099}; // @[Mux.scala 19:72:@3539.4]
  assign _T_1196 = _T_1195 | _GEN_211; // @[Mux.scala 19:72:@3539.4]
  assign _GEN_212 = {{24'd0}, _T_1101}; // @[Mux.scala 19:72:@3540.4]
  assign _T_1197 = _T_1196 | _GEN_212; // @[Mux.scala 19:72:@3540.4]
  assign _GEN_213 = {{24'd0}, _T_1103}; // @[Mux.scala 19:72:@3541.4]
  assign _T_1198 = _T_1197 | _GEN_213; // @[Mux.scala 19:72:@3541.4]
  assign _GEN_214 = {{24'd0}, _T_1105}; // @[Mux.scala 19:72:@3542.4]
  assign _T_1199 = _T_1198 | _GEN_214; // @[Mux.scala 19:72:@3542.4]
  assign _GEN_215 = {{24'd0}, _T_1107}; // @[Mux.scala 19:72:@3543.4]
  assign _T_1200 = _T_1199 | _GEN_215; // @[Mux.scala 19:72:@3543.4]
  assign _GEN_216 = {{24'd0}, _T_1109}; // @[Mux.scala 19:72:@3544.4]
  assign _T_1201 = _T_1200 | _GEN_216; // @[Mux.scala 19:72:@3544.4]
  assign _GEN_217 = {{24'd0}, _T_1111}; // @[Mux.scala 19:72:@3545.4]
  assign _T_1202 = _T_1201 | _GEN_217; // @[Mux.scala 19:72:@3545.4]
  assign _GEN_218 = {{24'd0}, _T_1113}; // @[Mux.scala 19:72:@3546.4]
  assign _T_1203 = _T_1202 | _GEN_218; // @[Mux.scala 19:72:@3546.4]
  assign _GEN_219 = {{24'd0}, _T_1115}; // @[Mux.scala 19:72:@3547.4]
  assign _T_1204 = _T_1203 | _GEN_219; // @[Mux.scala 19:72:@3547.4]
  assign _GEN_220 = {{24'd0}, _T_1117}; // @[Mux.scala 19:72:@3548.4]
  assign _T_1205 = _T_1204 | _GEN_220; // @[Mux.scala 19:72:@3548.4]
  assign _GEN_221 = {{24'd0}, _T_1119}; // @[Mux.scala 19:72:@3549.4]
  assign _T_1206 = _T_1205 | _GEN_221; // @[Mux.scala 19:72:@3549.4]
  assign _GEN_222 = {{24'd0}, _T_1121}; // @[Mux.scala 19:72:@3550.4]
  assign _T_1207 = _T_1206 | _GEN_222; // @[Mux.scala 19:72:@3550.4]
  assign _GEN_223 = {{24'd0}, _T_1123}; // @[Mux.scala 19:72:@3551.4]
  assign _T_1208 = _T_1207 | _GEN_223; // @[Mux.scala 19:72:@3551.4]
  assign _GEN_224 = {{24'd0}, _T_1125}; // @[Mux.scala 19:72:@3552.4]
  assign _T_1209 = _T_1208 | _GEN_224; // @[Mux.scala 19:72:@3552.4]
  assign _T_1220 = wdata[3]; // @[CSR.scala 245:39:@3565.8]
  assign _T_1222 = wdata[7]; // @[CSR.scala 245:39:@3569.8]
  assign _GEN_17 = _T_490 ? _T_1220 : _GEN_3; // @[CSR.scala 244:39:@3559.6]
  assign _GEN_18 = _T_490 ? _T_1222 : _GEN_4; // @[CSR.scala 244:39:@3559.6]
  assign _T_1233 = wdata[15:0]; // @[:@3588.8 :@3589.8]
  assign _T_1235 = _T_1233[3]; // @[CSR.scala 250:35:@3592.8]
  assign _T_1237 = _T_1233[7]; // @[CSR.scala 250:35:@3596.8]
  assign _GEN_19 = _T_494 ? _T_1235 : reg_mip_msip; // @[CSR.scala 249:35:@3586.6]
  assign _GEN_20 = _T_496 ? _T_1235 : reg_mie_msip; // @[CSR.scala 253:35:@3606.6]
  assign _GEN_21 = _T_496 ? _T_1237 : reg_mie_mtip; // @[CSR.scala 253:35:@3606.6]
  assign _T_1253 = wdata[7:0]; // @[CSR.scala 277:47:@3628.8]
  assign _T_1254 = _T_264[31:0]; // @[CSR.scala 277:72:@3629.8]
  assign _T_1255 = {_T_1253,_T_1254}; // @[Cat.scala 30:58:@3630.8]
  assign _GEN_22 = _T_514 ? {{1'd0}, _T_1255} : _T_265; // @[CSR.scala 277:29:@3627.6]
  assign _T_1256 = _T_264[39:32]; // @[CSR.scala 278:45:@3634.8]
  assign _T_1257 = {_T_1256,wdata}; // @[Cat.scala 30:58:@3635.8]
  assign _GEN_23 = _T_512 ? {{1'd0}, _T_1257} : _GEN_22; // @[CSR.scala 278:29:@3633.6]
  assign _T_1259 = _T_267[31:0]; // @[CSR.scala 277:72:@3640.8]
  assign _T_1260 = {_T_1253,_T_1259}; // @[Cat.scala 30:58:@3641.8]
  assign _GEN_24 = _T_518 ? {{1'd0}, _T_1260} : _T_268; // @[CSR.scala 277:29:@3638.6]
  assign _T_1261 = _T_267[39:32]; // @[CSR.scala 278:45:@3645.8]
  assign _T_1262 = {_T_1261,wdata}; // @[Cat.scala 30:58:@3646.8]
  assign _GEN_25 = _T_516 ? {{1'd0}, _T_1262} : _GEN_24; // @[CSR.scala 278:29:@3644.6]
  assign _T_1264 = _T_270[31:0]; // @[CSR.scala 277:72:@3651.8]
  assign _T_1265 = {_T_1253,_T_1264}; // @[Cat.scala 30:58:@3652.8]
  assign _GEN_26 = _T_522 ? {{1'd0}, _T_1265} : _T_271; // @[CSR.scala 277:29:@3649.6]
  assign _T_1266 = _T_270[39:32]; // @[CSR.scala 278:45:@3656.8]
  assign _T_1267 = {_T_1266,wdata}; // @[Cat.scala 30:58:@3657.8]
  assign _GEN_27 = _T_520 ? {{1'd0}, _T_1267} : _GEN_26; // @[CSR.scala 278:29:@3655.6]
  assign _T_1269 = _T_273[31:0]; // @[CSR.scala 277:72:@3662.8]
  assign _T_1270 = {_T_1253,_T_1269}; // @[Cat.scala 30:58:@3663.8]
  assign _GEN_28 = _T_526 ? {{1'd0}, _T_1270} : _T_274; // @[CSR.scala 277:29:@3660.6]
  assign _T_1271 = _T_273[39:32]; // @[CSR.scala 278:45:@3667.8]
  assign _T_1272 = {_T_1271,wdata}; // @[Cat.scala 30:58:@3668.8]
  assign _GEN_29 = _T_524 ? {{1'd0}, _T_1272} : _GEN_28; // @[CSR.scala 278:29:@3666.6]
  assign _T_1274 = _T_276[31:0]; // @[CSR.scala 277:72:@3673.8]
  assign _T_1275 = {_T_1253,_T_1274}; // @[Cat.scala 30:58:@3674.8]
  assign _GEN_30 = _T_530 ? {{1'd0}, _T_1275} : _T_277; // @[CSR.scala 277:29:@3671.6]
  assign _T_1276 = _T_276[39:32]; // @[CSR.scala 278:45:@3678.8]
  assign _T_1277 = {_T_1276,wdata}; // @[Cat.scala 30:58:@3679.8]
  assign _GEN_31 = _T_528 ? {{1'd0}, _T_1277} : _GEN_30; // @[CSR.scala 278:29:@3677.6]
  assign _T_1279 = _T_279[31:0]; // @[CSR.scala 277:72:@3684.8]
  assign _T_1280 = {_T_1253,_T_1279}; // @[Cat.scala 30:58:@3685.8]
  assign _GEN_32 = _T_534 ? {{1'd0}, _T_1280} : _T_280; // @[CSR.scala 277:29:@3682.6]
  assign _T_1281 = _T_279[39:32]; // @[CSR.scala 278:45:@3689.8]
  assign _T_1282 = {_T_1281,wdata}; // @[Cat.scala 30:58:@3690.8]
  assign _GEN_33 = _T_532 ? {{1'd0}, _T_1282} : _GEN_32; // @[CSR.scala 278:29:@3688.6]
  assign _T_1284 = _T_282[31:0]; // @[CSR.scala 277:72:@3695.8]
  assign _T_1285 = {_T_1253,_T_1284}; // @[Cat.scala 30:58:@3696.8]
  assign _GEN_34 = _T_538 ? {{1'd0}, _T_1285} : _T_283; // @[CSR.scala 277:29:@3693.6]
  assign _T_1286 = _T_282[39:32]; // @[CSR.scala 278:45:@3700.8]
  assign _T_1287 = {_T_1286,wdata}; // @[Cat.scala 30:58:@3701.8]
  assign _GEN_35 = _T_536 ? {{1'd0}, _T_1287} : _GEN_34; // @[CSR.scala 278:29:@3699.6]
  assign _T_1289 = _T_285[31:0]; // @[CSR.scala 277:72:@3706.8]
  assign _T_1290 = {_T_1253,_T_1289}; // @[Cat.scala 30:58:@3707.8]
  assign _GEN_36 = _T_542 ? {{1'd0}, _T_1290} : _T_286; // @[CSR.scala 277:29:@3704.6]
  assign _T_1291 = _T_285[39:32]; // @[CSR.scala 278:45:@3711.8]
  assign _T_1292 = {_T_1291,wdata}; // @[Cat.scala 30:58:@3712.8]
  assign _GEN_37 = _T_540 ? {{1'd0}, _T_1292} : _GEN_36; // @[CSR.scala 278:29:@3710.6]
  assign _T_1294 = _T_288[31:0]; // @[CSR.scala 277:72:@3717.8]
  assign _T_1295 = {_T_1253,_T_1294}; // @[Cat.scala 30:58:@3718.8]
  assign _GEN_38 = _T_546 ? {{1'd0}, _T_1295} : _T_289; // @[CSR.scala 277:29:@3715.6]
  assign _T_1296 = _T_288[39:32]; // @[CSR.scala 278:45:@3722.8]
  assign _T_1297 = {_T_1296,wdata}; // @[Cat.scala 30:58:@3723.8]
  assign _GEN_39 = _T_544 ? {{1'd0}, _T_1297} : _GEN_38; // @[CSR.scala 278:29:@3721.6]
  assign _T_1299 = _T_291[31:0]; // @[CSR.scala 277:72:@3728.8]
  assign _T_1300 = {_T_1253,_T_1299}; // @[Cat.scala 30:58:@3729.8]
  assign _GEN_40 = _T_550 ? {{1'd0}, _T_1300} : _T_292; // @[CSR.scala 277:29:@3726.6]
  assign _T_1301 = _T_291[39:32]; // @[CSR.scala 278:45:@3733.8]
  assign _T_1302 = {_T_1301,wdata}; // @[Cat.scala 30:58:@3734.8]
  assign _GEN_41 = _T_548 ? {{1'd0}, _T_1302} : _GEN_40; // @[CSR.scala 278:29:@3732.6]
  assign _T_1304 = _T_294[31:0]; // @[CSR.scala 277:72:@3739.8]
  assign _T_1305 = {_T_1253,_T_1304}; // @[Cat.scala 30:58:@3740.8]
  assign _GEN_42 = _T_554 ? {{1'd0}, _T_1305} : _T_295; // @[CSR.scala 277:29:@3737.6]
  assign _T_1306 = _T_294[39:32]; // @[CSR.scala 278:45:@3744.8]
  assign _T_1307 = {_T_1306,wdata}; // @[Cat.scala 30:58:@3745.8]
  assign _GEN_43 = _T_552 ? {{1'd0}, _T_1307} : _GEN_42; // @[CSR.scala 278:29:@3743.6]
  assign _T_1309 = _T_297[31:0]; // @[CSR.scala 277:72:@3750.8]
  assign _T_1310 = {_T_1253,_T_1309}; // @[Cat.scala 30:58:@3751.8]
  assign _GEN_44 = _T_558 ? {{1'd0}, _T_1310} : _T_298; // @[CSR.scala 277:29:@3748.6]
  assign _T_1311 = _T_297[39:32]; // @[CSR.scala 278:45:@3755.8]
  assign _T_1312 = {_T_1311,wdata}; // @[Cat.scala 30:58:@3756.8]
  assign _GEN_45 = _T_556 ? {{1'd0}, _T_1312} : _GEN_44; // @[CSR.scala 278:29:@3754.6]
  assign _T_1314 = _T_300[31:0]; // @[CSR.scala 277:72:@3761.8]
  assign _T_1315 = {_T_1253,_T_1314}; // @[Cat.scala 30:58:@3762.8]
  assign _GEN_46 = _T_562 ? {{1'd0}, _T_1315} : _T_301; // @[CSR.scala 277:29:@3759.6]
  assign _T_1316 = _T_300[39:32]; // @[CSR.scala 278:45:@3766.8]
  assign _T_1317 = {_T_1316,wdata}; // @[Cat.scala 30:58:@3767.8]
  assign _GEN_47 = _T_560 ? {{1'd0}, _T_1317} : _GEN_46; // @[CSR.scala 278:29:@3765.6]
  assign _T_1319 = _T_303[31:0]; // @[CSR.scala 277:72:@3772.8]
  assign _T_1320 = {_T_1253,_T_1319}; // @[Cat.scala 30:58:@3773.8]
  assign _GEN_48 = _T_566 ? {{1'd0}, _T_1320} : _T_304; // @[CSR.scala 277:29:@3770.6]
  assign _T_1321 = _T_303[39:32]; // @[CSR.scala 278:45:@3777.8]
  assign _T_1322 = {_T_1321,wdata}; // @[Cat.scala 30:58:@3778.8]
  assign _GEN_49 = _T_564 ? {{1'd0}, _T_1322} : _GEN_48; // @[CSR.scala 278:29:@3776.6]
  assign _T_1324 = _T_306[31:0]; // @[CSR.scala 277:72:@3783.8]
  assign _T_1325 = {_T_1253,_T_1324}; // @[Cat.scala 30:58:@3784.8]
  assign _GEN_50 = _T_570 ? {{1'd0}, _T_1325} : _T_307; // @[CSR.scala 277:29:@3781.6]
  assign _T_1326 = _T_306[39:32]; // @[CSR.scala 278:45:@3788.8]
  assign _T_1327 = {_T_1326,wdata}; // @[Cat.scala 30:58:@3789.8]
  assign _GEN_51 = _T_568 ? {{1'd0}, _T_1327} : _GEN_50; // @[CSR.scala 278:29:@3787.6]
  assign _T_1329 = _T_309[31:0]; // @[CSR.scala 277:72:@3794.8]
  assign _T_1330 = {_T_1253,_T_1329}; // @[Cat.scala 30:58:@3795.8]
  assign _GEN_52 = _T_574 ? {{1'd0}, _T_1330} : _T_310; // @[CSR.scala 277:29:@3792.6]
  assign _T_1331 = _T_309[39:32]; // @[CSR.scala 278:45:@3799.8]
  assign _T_1332 = {_T_1331,wdata}; // @[Cat.scala 30:58:@3800.8]
  assign _GEN_53 = _T_572 ? {{1'd0}, _T_1332} : _GEN_52; // @[CSR.scala 278:29:@3798.6]
  assign _T_1334 = _T_312[31:0]; // @[CSR.scala 277:72:@3805.8]
  assign _T_1335 = {_T_1253,_T_1334}; // @[Cat.scala 30:58:@3806.8]
  assign _GEN_54 = _T_578 ? {{1'd0}, _T_1335} : _T_313; // @[CSR.scala 277:29:@3803.6]
  assign _T_1336 = _T_312[39:32]; // @[CSR.scala 278:45:@3810.8]
  assign _T_1337 = {_T_1336,wdata}; // @[Cat.scala 30:58:@3811.8]
  assign _GEN_55 = _T_576 ? {{1'd0}, _T_1337} : _GEN_54; // @[CSR.scala 278:29:@3809.6]
  assign _T_1339 = _T_315[31:0]; // @[CSR.scala 277:72:@3816.8]
  assign _T_1340 = {_T_1253,_T_1339}; // @[Cat.scala 30:58:@3817.8]
  assign _GEN_56 = _T_582 ? {{1'd0}, _T_1340} : _T_316; // @[CSR.scala 277:29:@3814.6]
  assign _T_1341 = _T_315[39:32]; // @[CSR.scala 278:45:@3821.8]
  assign _T_1342 = {_T_1341,wdata}; // @[Cat.scala 30:58:@3822.8]
  assign _GEN_57 = _T_580 ? {{1'd0}, _T_1342} : _GEN_56; // @[CSR.scala 278:29:@3820.6]
  assign _T_1344 = _T_318[31:0]; // @[CSR.scala 277:72:@3827.8]
  assign _T_1345 = {_T_1253,_T_1344}; // @[Cat.scala 30:58:@3828.8]
  assign _GEN_58 = _T_586 ? {{1'd0}, _T_1345} : _T_319; // @[CSR.scala 277:29:@3825.6]
  assign _T_1346 = _T_318[39:32]; // @[CSR.scala 278:45:@3832.8]
  assign _T_1347 = {_T_1346,wdata}; // @[Cat.scala 30:58:@3833.8]
  assign _GEN_59 = _T_584 ? {{1'd0}, _T_1347} : _GEN_58; // @[CSR.scala 278:29:@3831.6]
  assign _T_1349 = _T_321[31:0]; // @[CSR.scala 277:72:@3838.8]
  assign _T_1350 = {_T_1253,_T_1349}; // @[Cat.scala 30:58:@3839.8]
  assign _GEN_60 = _T_590 ? {{1'd0}, _T_1350} : _T_322; // @[CSR.scala 277:29:@3836.6]
  assign _T_1351 = _T_321[39:32]; // @[CSR.scala 278:45:@3843.8]
  assign _T_1352 = {_T_1351,wdata}; // @[Cat.scala 30:58:@3844.8]
  assign _GEN_61 = _T_588 ? {{1'd0}, _T_1352} : _GEN_60; // @[CSR.scala 278:29:@3842.6]
  assign _T_1354 = _T_324[31:0]; // @[CSR.scala 277:72:@3849.8]
  assign _T_1355 = {_T_1253,_T_1354}; // @[Cat.scala 30:58:@3850.8]
  assign _GEN_62 = _T_594 ? {{1'd0}, _T_1355} : _T_325; // @[CSR.scala 277:29:@3847.6]
  assign _T_1356 = _T_324[39:32]; // @[CSR.scala 278:45:@3854.8]
  assign _T_1357 = {_T_1356,wdata}; // @[Cat.scala 30:58:@3855.8]
  assign _GEN_63 = _T_592 ? {{1'd0}, _T_1357} : _GEN_62; // @[CSR.scala 278:29:@3853.6]
  assign _T_1359 = _T_327[31:0]; // @[CSR.scala 277:72:@3860.8]
  assign _T_1360 = {_T_1253,_T_1359}; // @[Cat.scala 30:58:@3861.8]
  assign _GEN_64 = _T_598 ? {{1'd0}, _T_1360} : _T_328; // @[CSR.scala 277:29:@3858.6]
  assign _T_1361 = _T_327[39:32]; // @[CSR.scala 278:45:@3865.8]
  assign _T_1362 = {_T_1361,wdata}; // @[Cat.scala 30:58:@3866.8]
  assign _GEN_65 = _T_596 ? {{1'd0}, _T_1362} : _GEN_64; // @[CSR.scala 278:29:@3864.6]
  assign _T_1364 = _T_330[31:0]; // @[CSR.scala 277:72:@3871.8]
  assign _T_1365 = {_T_1253,_T_1364}; // @[Cat.scala 30:58:@3872.8]
  assign _GEN_66 = _T_602 ? {{1'd0}, _T_1365} : _T_331; // @[CSR.scala 277:29:@3869.6]
  assign _T_1366 = _T_330[39:32]; // @[CSR.scala 278:45:@3876.8]
  assign _T_1367 = {_T_1366,wdata}; // @[Cat.scala 30:58:@3877.8]
  assign _GEN_67 = _T_600 ? {{1'd0}, _T_1367} : _GEN_66; // @[CSR.scala 278:29:@3875.6]
  assign _T_1369 = _T_333[31:0]; // @[CSR.scala 277:72:@3882.8]
  assign _T_1370 = {_T_1253,_T_1369}; // @[Cat.scala 30:58:@3883.8]
  assign _GEN_68 = _T_606 ? {{1'd0}, _T_1370} : _T_334; // @[CSR.scala 277:29:@3880.6]
  assign _T_1371 = _T_333[39:32]; // @[CSR.scala 278:45:@3887.8]
  assign _T_1372 = {_T_1371,wdata}; // @[Cat.scala 30:58:@3888.8]
  assign _GEN_69 = _T_604 ? {{1'd0}, _T_1372} : _GEN_68; // @[CSR.scala 278:29:@3886.6]
  assign _T_1374 = _T_336[31:0]; // @[CSR.scala 277:72:@3893.8]
  assign _T_1375 = {_T_1253,_T_1374}; // @[Cat.scala 30:58:@3894.8]
  assign _GEN_70 = _T_610 ? {{1'd0}, _T_1375} : _T_337; // @[CSR.scala 277:29:@3891.6]
  assign _T_1376 = _T_336[39:32]; // @[CSR.scala 278:45:@3898.8]
  assign _T_1377 = {_T_1376,wdata}; // @[Cat.scala 30:58:@3899.8]
  assign _GEN_71 = _T_608 ? {{1'd0}, _T_1377} : _GEN_70; // @[CSR.scala 278:29:@3897.6]
  assign _T_1379 = _T_339[31:0]; // @[CSR.scala 277:72:@3904.8]
  assign _T_1380 = {_T_1253,_T_1379}; // @[Cat.scala 30:58:@3905.8]
  assign _GEN_72 = _T_614 ? {{1'd0}, _T_1380} : _T_340; // @[CSR.scala 277:29:@3902.6]
  assign _T_1381 = _T_339[39:32]; // @[CSR.scala 278:45:@3909.8]
  assign _T_1382 = {_T_1381,wdata}; // @[Cat.scala 30:58:@3910.8]
  assign _GEN_73 = _T_612 ? {{1'd0}, _T_1382} : _GEN_72; // @[CSR.scala 278:29:@3908.6]
  assign _T_1384 = _T_342[31:0]; // @[CSR.scala 277:72:@3915.8]
  assign _T_1385 = {_T_1253,_T_1384}; // @[Cat.scala 30:58:@3916.8]
  assign _GEN_74 = _T_618 ? {{1'd0}, _T_1385} : _T_343; // @[CSR.scala 277:29:@3913.6]
  assign _T_1386 = _T_342[39:32]; // @[CSR.scala 278:45:@3920.8]
  assign _T_1387 = {_T_1386,wdata}; // @[Cat.scala 30:58:@3921.8]
  assign _GEN_75 = _T_616 ? {{1'd0}, _T_1387} : _GEN_74; // @[CSR.scala 278:29:@3919.6]
  assign _T_1389 = _T_345[31:0]; // @[CSR.scala 277:72:@3926.8]
  assign _T_1390 = {_T_1253,_T_1389}; // @[Cat.scala 30:58:@3927.8]
  assign _GEN_76 = _T_622 ? {{1'd0}, _T_1390} : _T_346; // @[CSR.scala 277:29:@3924.6]
  assign _T_1391 = _T_345[39:32]; // @[CSR.scala 278:45:@3931.8]
  assign _T_1392 = {_T_1391,wdata}; // @[Cat.scala 30:58:@3932.8]
  assign _GEN_77 = _T_620 ? {{1'd0}, _T_1392} : _GEN_76; // @[CSR.scala 278:29:@3930.6]
  assign _T_1394 = _T_348[31:0]; // @[CSR.scala 277:72:@3937.8]
  assign _T_1395 = {_T_1253,_T_1394}; // @[Cat.scala 30:58:@3938.8]
  assign _GEN_78 = _T_626 ? {{1'd0}, _T_1395} : _T_349; // @[CSR.scala 277:29:@3935.6]
  assign _T_1396 = _T_348[39:32]; // @[CSR.scala 278:45:@3942.8]
  assign _T_1397 = {_T_1396,wdata}; // @[Cat.scala 30:58:@3943.8]
  assign _GEN_79 = _T_624 ? {{1'd0}, _T_1397} : _GEN_78; // @[CSR.scala 278:29:@3941.6]
  assign _T_1399 = _T_351[31:0]; // @[CSR.scala 277:72:@3948.8]
  assign _T_1400 = {_T_1253,_T_1399}; // @[Cat.scala 30:58:@3949.8]
  assign _GEN_80 = _T_630 ? {{1'd0}, _T_1400} : _T_352; // @[CSR.scala 277:29:@3946.6]
  assign _T_1401 = _T_351[39:32]; // @[CSR.scala 278:45:@3953.8]
  assign _T_1402 = {_T_1401,wdata}; // @[Cat.scala 30:58:@3954.8]
  assign _GEN_81 = _T_628 ? {{1'd0}, _T_1402} : _GEN_80; // @[CSR.scala 278:29:@3952.6]
  assign _T_1404 = _T_354[31:0]; // @[CSR.scala 277:72:@3959.8]
  assign _T_1405 = {_T_1253,_T_1404}; // @[Cat.scala 30:58:@3960.8]
  assign _GEN_82 = _T_634 ? {{1'd0}, _T_1405} : _T_355; // @[CSR.scala 277:29:@3957.6]
  assign _T_1406 = _T_354[39:32]; // @[CSR.scala 278:45:@3964.8]
  assign _T_1407 = {_T_1406,wdata}; // @[Cat.scala 30:58:@3965.8]
  assign _GEN_83 = _T_632 ? {{1'd0}, _T_1407} : _GEN_82; // @[CSR.scala 278:29:@3963.6]
  assign _T_1409 = _T_357[31:0]; // @[CSR.scala 277:72:@3970.8]
  assign _T_1410 = {_T_1253,_T_1409}; // @[Cat.scala 30:58:@3971.8]
  assign _GEN_84 = _T_638 ? {{1'd0}, _T_1410} : _T_358; // @[CSR.scala 277:29:@3968.6]
  assign _T_1411 = _T_357[39:32]; // @[CSR.scala 278:45:@3975.8]
  assign _T_1412 = {_T_1411,wdata}; // @[Cat.scala 30:58:@3976.8]
  assign _GEN_85 = _T_636 ? {{1'd0}, _T_1412} : _GEN_84; // @[CSR.scala 278:29:@3974.6]
  assign _T_1414 = _T_249[31:0]; // @[CSR.scala 277:72:@3981.8]
  assign _T_1415 = {wdata,_T_1414}; // @[Cat.scala 30:58:@3982.8]
  assign _T_1416 = _T_1415[63:6]; // @[Util.scala 133:28:@3984.8]
  assign _GEN_86 = _T_640 ? _T_1415 : {{57'd0}, _T_241}; // @[CSR.scala 277:29:@3979.6]
  assign _GEN_87 = _T_640 ? _T_1416 : _GEN_0; // @[CSR.scala 277:29:@3979.6]
  assign _T_1417 = _T_249[63:32]; // @[CSR.scala 278:45:@3988.8]
  assign _T_1418 = {_T_1417,wdata}; // @[Cat.scala 30:58:@3989.8]
  assign _T_1419 = _T_1418[63:6]; // @[Util.scala 133:28:@3991.8]
  assign _GEN_88 = _T_478 ? _T_1418 : _GEN_86; // @[CSR.scala 278:29:@3987.6]
  assign _GEN_89 = _T_478 ? _T_1419 : _GEN_87; // @[CSR.scala 278:29:@3987.6]
  assign _T_1421 = _T_261[31:0]; // @[CSR.scala 277:72:@3996.8]
  assign _T_1422 = {wdata,_T_1421}; // @[Cat.scala 30:58:@3997.8]
  assign _T_1423 = _T_1422[63:6]; // @[Util.scala 133:28:@3999.8]
  assign _GEN_90 = _T_642 ? _T_1422 : {{57'd0}, _T_253}; // @[CSR.scala 277:29:@3994.6]
  assign _GEN_91 = _T_642 ? _T_1423 : _GEN_1; // @[CSR.scala 277:29:@3994.6]
  assign _T_1424 = _T_261[63:32]; // @[CSR.scala 278:45:@4003.8]
  assign _T_1425 = {_T_1424,wdata}; // @[Cat.scala 30:58:@4004.8]
  assign _T_1426 = _T_1425[63:6]; // @[Util.scala 133:28:@4006.8]
  assign _GEN_92 = _T_480 ? _T_1425 : _GEN_90; // @[CSR.scala 278:29:@4002.6]
  assign _GEN_93 = _T_480 ? _T_1426 : _GEN_91; // @[CSR.scala 278:29:@4002.6]
  assign _GEN_94 = _T_508 ? wdata : reg_dscratch; // @[CSR.scala 265:40:@4009.6]
  assign _T_1429 = wdata >> 2'h2; // @[CSR.scala 267:78:@4014.8]
  assign _GEN_225 = {{3'd0}, _T_1429}; // @[CSR.scala 267:86:@4015.8]
  assign _T_1431 = _GEN_225 << 2'h2; // @[CSR.scala 267:86:@4015.8]
  assign _GEN_95 = _T_500 ? _T_1431 : {{3'd0}, _GEN_15}; // @[CSR.scala 267:40:@4012.6]
  assign _GEN_96 = _T_498 ? wdata : reg_mscratch; // @[CSR.scala 268:40:@4018.6]
  assign _T_1433 = wdata & 32'h8000001f; // @[CSR.scala 269:62:@4022.8]
  assign _GEN_97 = _T_504 ? _T_1433 : _GEN_14; // @[CSR.scala 269:40:@4021.6]
  assign _GEN_98 = _T_502 ? wdata : _GEN_16; // @[CSR.scala 270:40:@4025.6]
  assign _GEN_99 = _T_510 ? wdata : reg_medeleg; // @[CSR.scala 271:42:@4029.6]
  assign _GEN_100 = wen ? _GEN_17 : _GEN_3; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_101 = wen ? _GEN_18 : _GEN_4; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_102 = wen ? _GEN_19 : reg_mip_msip; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_103 = wen ? _GEN_20 : reg_mie_msip; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_104 = wen ? _GEN_21 : reg_mie_mtip; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_105 = wen ? _GEN_23 : _T_265; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_106 = wen ? _GEN_25 : _T_268; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_107 = wen ? _GEN_27 : _T_271; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_108 = wen ? _GEN_29 : _T_274; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_109 = wen ? _GEN_31 : _T_277; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_110 = wen ? _GEN_33 : _T_280; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_111 = wen ? _GEN_35 : _T_283; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_112 = wen ? _GEN_37 : _T_286; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_113 = wen ? _GEN_39 : _T_289; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_114 = wen ? _GEN_41 : _T_292; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_115 = wen ? _GEN_43 : _T_295; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_116 = wen ? _GEN_45 : _T_298; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_117 = wen ? _GEN_47 : _T_301; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_118 = wen ? _GEN_49 : _T_304; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_119 = wen ? _GEN_51 : _T_307; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_120 = wen ? _GEN_53 : _T_310; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_121 = wen ? _GEN_55 : _T_313; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_122 = wen ? _GEN_57 : _T_316; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_123 = wen ? _GEN_59 : _T_319; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_124 = wen ? _GEN_61 : _T_322; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_125 = wen ? _GEN_63 : _T_325; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_126 = wen ? _GEN_65 : _T_328; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_127 = wen ? _GEN_67 : _T_331; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_128 = wen ? _GEN_69 : _T_334; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_129 = wen ? _GEN_71 : _T_337; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_130 = wen ? _GEN_73 : _T_340; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_131 = wen ? _GEN_75 : _T_343; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_132 = wen ? _GEN_77 : _T_346; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_133 = wen ? _GEN_79 : _T_349; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_134 = wen ? _GEN_81 : _T_352; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_135 = wen ? _GEN_83 : _T_355; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_136 = wen ? _GEN_85 : _T_358; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_137 = wen ? _GEN_88 : {{57'd0}, _T_241}; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_138 = wen ? _GEN_89 : _GEN_0; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_139 = wen ? _GEN_92 : {{57'd0}, _T_253}; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_140 = wen ? _GEN_93 : _GEN_1; // @[CSR.scala 242:14:@3558.4]
  assign _GEN_142 = wen ? _GEN_95 : {{3'd0}, _GEN_15}; // @[CSR.scala 242:14:@3558.4]
  assign io_rw_rdata = _T_1209[31:0]; // @[CSR.scala 240:15:@3557.4]
  assign io_eret = _T_940 | insn_ret; // @[CSR.scala 199:11:@3347.4]
  assign io_status_prv = reg_mstatus_prv; // @[CSR.scala 197:13:@3344.4]
  assign io_status_unimp5 = 14'h0; // @[CSR.scala 197:13:@3343.4]
  assign io_status_mprv = 1'h0; // @[CSR.scala 197:13:@3342.4]
  assign io_status_unimp4 = 2'h0; // @[CSR.scala 197:13:@3341.4]
  assign io_status_mpp = 2'h3; // @[CSR.scala 197:13:@3340.4]
  assign io_status_unimp3 = 3'h0; // @[CSR.scala 197:13:@3339.4]
  assign io_status_mpie = reg_mstatus_mpie; // @[CSR.scala 197:13:@3338.4]
  assign io_status_unimp2 = 3'h0; // @[CSR.scala 197:13:@3337.4]
  assign io_status_mie = reg_mstatus_mie; // @[CSR.scala 197:13:@3336.4]
  assign io_status_unimp1 = 3'h0; // @[CSR.scala 197:13:@3335.4]
  assign io_evec = io_xcpt ? 32'h80000004 : _GEN_10; // @[CSR.scala 212:13:@3368.6 CSR.scala 217:13:@3371.6 CSR.scala 224:13:@3378.6 CSR.scala 230:13:@3383.6]
  assign io_time = _T_249[31:0]; // @[CSR.scala 236:11:@3388.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  reg_mstatus_prv = _RAND_0[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  reg_mstatus_mpie = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  reg_mstatus_mie = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  reg_mepc = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  reg_mcause = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  reg_mtval = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  reg_mscratch = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  reg_medeleg = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  reg_mip_mtip = _RAND_8[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  reg_mip_msip = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  reg_mie_mtip = _RAND_10[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  reg_mie_msip = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  _T_240 = _RAND_12[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {2{`RANDOM}};
  _T_244 = _RAND_13[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  _T_252 = _RAND_14[5:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {2{`RANDOM}};
  _T_256 = _RAND_15[57:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {2{`RANDOM}};
  _T_264 = _RAND_16[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {2{`RANDOM}};
  _T_267 = _RAND_17[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {2{`RANDOM}};
  _T_270 = _RAND_18[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {2{`RANDOM}};
  _T_273 = _RAND_19[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {2{`RANDOM}};
  _T_276 = _RAND_20[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {2{`RANDOM}};
  _T_279 = _RAND_21[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {2{`RANDOM}};
  _T_282 = _RAND_22[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {2{`RANDOM}};
  _T_285 = _RAND_23[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {2{`RANDOM}};
  _T_288 = _RAND_24[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {2{`RANDOM}};
  _T_291 = _RAND_25[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {2{`RANDOM}};
  _T_294 = _RAND_26[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {2{`RANDOM}};
  _T_297 = _RAND_27[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {2{`RANDOM}};
  _T_300 = _RAND_28[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {2{`RANDOM}};
  _T_303 = _RAND_29[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {2{`RANDOM}};
  _T_306 = _RAND_30[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {2{`RANDOM}};
  _T_309 = _RAND_31[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {2{`RANDOM}};
  _T_312 = _RAND_32[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {2{`RANDOM}};
  _T_315 = _RAND_33[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {2{`RANDOM}};
  _T_318 = _RAND_34[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {2{`RANDOM}};
  _T_321 = _RAND_35[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {2{`RANDOM}};
  _T_324 = _RAND_36[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {2{`RANDOM}};
  _T_327 = _RAND_37[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {2{`RANDOM}};
  _T_330 = _RAND_38[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {2{`RANDOM}};
  _T_333 = _RAND_39[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {2{`RANDOM}};
  _T_336 = _RAND_40[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {2{`RANDOM}};
  _T_339 = _RAND_41[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {2{`RANDOM}};
  _T_342 = _RAND_42[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {2{`RANDOM}};
  _T_345 = _RAND_43[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {2{`RANDOM}};
  _T_348 = _RAND_44[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {2{`RANDOM}};
  _T_351 = _RAND_45[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {2{`RANDOM}};
  _T_354 = _RAND_46[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {2{`RANDOM}};
  _T_357 = _RAND_47[39:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{`RANDOM}};
  reg_dscratch = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_mstatus_prv <= 2'h3;
    end else begin
      if (_T_954) begin
        reg_mstatus_prv <= 2'h3;
      end
    end
    if (reset) begin
      reg_mstatus_mpie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mpie <= _T_1222;
        end else begin
          if (_T_954) begin
            reg_mstatus_mpie <= 1'h1;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mpie <= 1'h1;
        end
      end
    end
    if (reset) begin
      reg_mstatus_mie <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_490) begin
          reg_mstatus_mie <= _T_1220;
        end else begin
          if (_T_954) begin
            reg_mstatus_mie <= reg_mstatus_mpie;
          end
        end
      end else begin
        if (_T_954) begin
          reg_mstatus_mie <= reg_mstatus_mpie;
        end
      end
    end
    reg_mepc <= _GEN_142[31:0];
    if (wen) begin
      if (_T_504) begin
        reg_mcause <= _T_1433;
      end else begin
        if (io_xcpt) begin
          reg_mcause <= io_cause;
        end else begin
          if (insn_break) begin
            reg_mcause <= 32'h3;
          end else begin
            if (insn_call) begin
              reg_mcause <= {{28'd0}, _T_959};
            end
          end
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mcause <= io_cause;
      end else begin
        if (insn_break) begin
          reg_mcause <= 32'h3;
        end else begin
          if (insn_call) begin
            reg_mcause <= {{28'd0}, _T_959};
          end
        end
      end
    end
    if (wen) begin
      if (_T_502) begin
        reg_mtval <= wdata;
      end else begin
        if (io_xcpt) begin
          reg_mtval <= io_tval;
        end
      end
    end else begin
      if (io_xcpt) begin
        reg_mtval <= io_tval;
      end
    end
    if (wen) begin
      if (_T_498) begin
        reg_mscratch <= wdata;
      end
    end
    if (wen) begin
      if (_T_510) begin
        reg_medeleg <= wdata;
      end
    end
    if (reset) begin
      reg_mip_mtip <= 1'h0;
    end else begin
      reg_mip_mtip <= 1'h1;
    end
    if (reset) begin
      reg_mip_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_494) begin
          reg_mip_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      reg_mie_mtip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_mtip <= _T_1237;
        end
      end
    end
    if (reset) begin
      reg_mie_msip <= 1'h0;
    end else begin
      if (wen) begin
        if (_T_496) begin
          reg_mie_msip <= _T_1235;
        end
      end
    end
    if (reset) begin
      _T_240 <= 6'h0;
    end else begin
      _T_240 <= _GEN_137[5:0];
    end
    if (reset) begin
      _T_244 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_478) begin
          _T_244 <= _T_1419;
        end else begin
          if (_T_640) begin
            _T_244 <= _T_1416;
          end else begin
            if (_T_245) begin
              _T_244 <= _T_248;
            end
          end
        end
      end else begin
        if (_T_245) begin
          _T_244 <= _T_248;
        end
      end
    end
    if (reset) begin
      _T_252 <= 6'h0;
    end else begin
      _T_252 <= _GEN_139[5:0];
    end
    if (reset) begin
      _T_256 <= 58'h0;
    end else begin
      if (wen) begin
        if (_T_480) begin
          _T_256 <= _T_1426;
        end else begin
          if (_T_642) begin
            _T_256 <= _T_1423;
          end else begin
            if (_T_257) begin
              _T_256 <= _T_260;
            end
          end
        end
      end else begin
        if (_T_257) begin
          _T_256 <= _T_260;
        end
      end
    end
    _T_264 <= _GEN_105[39:0];
    _T_267 <= _GEN_106[39:0];
    _T_270 <= _GEN_107[39:0];
    _T_273 <= _GEN_108[39:0];
    _T_276 <= _GEN_109[39:0];
    _T_279 <= _GEN_110[39:0];
    _T_282 <= _GEN_111[39:0];
    _T_285 <= _GEN_112[39:0];
    _T_288 <= _GEN_113[39:0];
    _T_291 <= _GEN_114[39:0];
    _T_294 <= _GEN_115[39:0];
    _T_297 <= _GEN_116[39:0];
    _T_300 <= _GEN_117[39:0];
    _T_303 <= _GEN_118[39:0];
    _T_306 <= _GEN_119[39:0];
    _T_309 <= _GEN_120[39:0];
    _T_312 <= _GEN_121[39:0];
    _T_315 <= _GEN_122[39:0];
    _T_318 <= _GEN_123[39:0];
    _T_321 <= _GEN_124[39:0];
    _T_324 <= _GEN_125[39:0];
    _T_327 <= _GEN_126[39:0];
    _T_330 <= _GEN_127[39:0];
    _T_333 <= _GEN_128[39:0];
    _T_336 <= _GEN_129[39:0];
    _T_339 <= _GEN_130[39:0];
    _T_342 <= _GEN_131[39:0];
    _T_345 <= _GEN_132[39:0];
    _T_348 <= _GEN_133[39:0];
    _T_351 <= _GEN_134[39:0];
    _T_354 <= _GEN_135[39:0];
    _T_357 <= _GEN_136[39:0];
    if (wen) begin
      if (_T_508) begin
        reg_dscratch <= wdata;
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_948) begin
          $fwrite(32'h80000002,"Assertion failed: these conditions must be mutually exclusive\n    at CSR.scala:201 assert(PopCount(insn_ret :: io.illegal :: Nil) <= 1, \"these conditions must be mutually exclusive\")\n"); // @[CSR.scala 201:9:@3354.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef STOP_COND
      if (`STOP_COND) begin
    `endif
        if (_T_948) begin
          $fatal; // @[CSR.scala 201:9:@3355.6]
        end
    `ifdef STOP_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module InstDecoder( // @[:@4035.2]
  input  [31:0] io_inst, // @[:@4038.4]
  output [3:0]  io_cinfo_br_type, // @[:@4038.4]
  output [1:0]  io_cinfo_op1_sel, // @[:@4038.4]
  output [2:0]  io_cinfo_op2_sel, // @[:@4038.4]
  output        io_cinfo_rs1_oen, // @[:@4038.4]
  output        io_cinfo_rs2_oen, // @[:@4038.4]
  output [3:0]  io_cinfo_alu_fun, // @[:@4038.4]
  output [1:0]  io_cinfo_wb_sel, // @[:@4038.4]
  output        io_cinfo_rf_wen, // @[:@4038.4]
  output        io_cinfo_mem_en, // @[:@4038.4]
  output        io_cinfo_mem_fcn, // @[:@4038.4]
  output [2:0]  io_cinfo_mem_typ, // @[:@4038.4]
  output [2:0]  io_cinfo_csr_cmd, // @[:@4038.4]
  output        io_cinfo_illegal, // @[:@4038.4]
  output        io_cinfo_fencei, // @[:@4038.4]
  output        io_cinfo_is_branch, // @[:@4038.4]
  output        io_cinfo_push, // @[:@4038.4]
  output        io_cinfo_pop, // @[:@4038.4]
  output [4:0]  io_cinfo_rs1_addr, // @[:@4038.4]
  output [4:0]  io_cinfo_rs2_addr, // @[:@4038.4]
  output [4:0]  io_cinfo_wbaddr, // @[:@4038.4]
  output [31:0] io_dinfo_imm_i, // @[:@4038.4]
  output [31:0] io_dinfo_imm_s, // @[:@4038.4]
  output [31:0] io_dinfo_imm_sb, // @[:@4038.4]
  output [31:0] io_dinfo_imm_u, // @[:@4038.4]
  output [31:0] io_dinfo_imm_uj, // @[:@4038.4]
  output [31:0] io_dinfo_imm_z // @[:@4038.4]
);
  wire [31:0] _T_13; // @[Lookup.scala 9:38:@4040.4]
  wire  _T_14; // @[Lookup.scala 9:38:@4041.4]
  wire  _T_18; // @[Lookup.scala 9:38:@4043.4]
  wire  _T_22; // @[Lookup.scala 9:38:@4045.4]
  wire  _T_26; // @[Lookup.scala 9:38:@4047.4]
  wire  _T_30; // @[Lookup.scala 9:38:@4049.4]
  wire  _T_34; // @[Lookup.scala 9:38:@4051.4]
  wire  _T_38; // @[Lookup.scala 9:38:@4053.4]
  wire  _T_42; // @[Lookup.scala 9:38:@4055.4]
  wire [31:0] _T_45; // @[Lookup.scala 9:38:@4056.4]
  wire  _T_46; // @[Lookup.scala 9:38:@4057.4]
  wire  _T_50; // @[Lookup.scala 9:38:@4059.4]
  wire  _T_54; // @[Lookup.scala 9:38:@4061.4]
  wire  _T_58; // @[Lookup.scala 9:38:@4063.4]
  wire  _T_62; // @[Lookup.scala 9:38:@4065.4]
  wire  _T_66; // @[Lookup.scala 9:38:@4067.4]
  wire  _T_70; // @[Lookup.scala 9:38:@4069.4]
  wire  _T_74; // @[Lookup.scala 9:38:@4071.4]
  wire [31:0] _T_77; // @[Lookup.scala 9:38:@4072.4]
  wire  _T_78; // @[Lookup.scala 9:38:@4073.4]
  wire  _T_82; // @[Lookup.scala 9:38:@4075.4]
  wire  _T_86; // @[Lookup.scala 9:38:@4077.4]
  wire [31:0] _T_89; // @[Lookup.scala 9:38:@4078.4]
  wire  _T_90; // @[Lookup.scala 9:38:@4079.4]
  wire  _T_94; // @[Lookup.scala 9:38:@4081.4]
  wire  _T_98; // @[Lookup.scala 9:38:@4083.4]
  wire  _T_102; // @[Lookup.scala 9:38:@4085.4]
  wire  _T_106; // @[Lookup.scala 9:38:@4087.4]
  wire  _T_110; // @[Lookup.scala 9:38:@4089.4]
  wire  _T_114; // @[Lookup.scala 9:38:@4091.4]
  wire  _T_118; // @[Lookup.scala 9:38:@4093.4]
  wire  _T_122; // @[Lookup.scala 9:38:@4095.4]
  wire  _T_126; // @[Lookup.scala 9:38:@4097.4]
  wire  _T_130; // @[Lookup.scala 9:38:@4099.4]
  wire  _T_134; // @[Lookup.scala 9:38:@4101.4]
  wire  _T_138; // @[Lookup.scala 9:38:@4103.4]
  wire  _T_142; // @[Lookup.scala 9:38:@4105.4]
  wire  _T_146; // @[Lookup.scala 9:38:@4107.4]
  wire  _T_150; // @[Lookup.scala 9:38:@4109.4]
  wire  _T_154; // @[Lookup.scala 9:38:@4111.4]
  wire  _T_158; // @[Lookup.scala 9:38:@4113.4]
  wire  _T_162; // @[Lookup.scala 9:38:@4115.4]
  wire  _T_166; // @[Lookup.scala 9:38:@4117.4]
  wire  _T_170; // @[Lookup.scala 9:38:@4119.4]
  wire  _T_174; // @[Lookup.scala 9:38:@4121.4]
  wire  _T_178; // @[Lookup.scala 9:38:@4123.4]
  wire  _T_182; // @[Lookup.scala 9:38:@4125.4]
  wire  _T_186; // @[Lookup.scala 9:38:@4127.4]
  wire  _T_190; // @[Lookup.scala 9:38:@4129.4]
  wire  _T_194; // @[Lookup.scala 9:38:@4131.4]
  wire  _T_198; // @[Lookup.scala 9:38:@4133.4]
  wire  _T_202; // @[Lookup.scala 9:38:@4135.4]
  wire  _T_206; // @[Lookup.scala 9:38:@4137.4]
  wire  _T_210; // @[Lookup.scala 9:38:@4139.4]
  wire  _T_212; // @[Lookup.scala 11:37:@4141.4]
  wire  _T_213; // @[Lookup.scala 11:37:@4142.4]
  wire  _T_214; // @[Lookup.scala 11:37:@4143.4]
  wire  _T_215; // @[Lookup.scala 11:37:@4144.4]
  wire  _T_216; // @[Lookup.scala 11:37:@4145.4]
  wire  _T_217; // @[Lookup.scala 11:37:@4146.4]
  wire  _T_218; // @[Lookup.scala 11:37:@4147.4]
  wire  _T_219; // @[Lookup.scala 11:37:@4148.4]
  wire  _T_220; // @[Lookup.scala 11:37:@4149.4]
  wire  _T_221; // @[Lookup.scala 11:37:@4150.4]
  wire  _T_222; // @[Lookup.scala 11:37:@4151.4]
  wire  _T_223; // @[Lookup.scala 11:37:@4152.4]
  wire  _T_224; // @[Lookup.scala 11:37:@4153.4]
  wire  _T_225; // @[Lookup.scala 11:37:@4154.4]
  wire  _T_226; // @[Lookup.scala 11:37:@4155.4]
  wire  _T_227; // @[Lookup.scala 11:37:@4156.4]
  wire  _T_228; // @[Lookup.scala 11:37:@4157.4]
  wire  _T_229; // @[Lookup.scala 11:37:@4158.4]
  wire  _T_230; // @[Lookup.scala 11:37:@4159.4]
  wire  _T_231; // @[Lookup.scala 11:37:@4160.4]
  wire  _T_232; // @[Lookup.scala 11:37:@4161.4]
  wire  _T_233; // @[Lookup.scala 11:37:@4162.4]
  wire  _T_234; // @[Lookup.scala 11:37:@4163.4]
  wire  _T_235; // @[Lookup.scala 11:37:@4164.4]
  wire  _T_236; // @[Lookup.scala 11:37:@4165.4]
  wire  _T_237; // @[Lookup.scala 11:37:@4166.4]
  wire  _T_238; // @[Lookup.scala 11:37:@4167.4]
  wire  _T_239; // @[Lookup.scala 11:37:@4168.4]
  wire  _T_240; // @[Lookup.scala 11:37:@4169.4]
  wire  _T_241; // @[Lookup.scala 11:37:@4170.4]
  wire  _T_242; // @[Lookup.scala 11:37:@4171.4]
  wire  _T_243; // @[Lookup.scala 11:37:@4172.4]
  wire  _T_244; // @[Lookup.scala 11:37:@4173.4]
  wire  _T_245; // @[Lookup.scala 11:37:@4174.4]
  wire  _T_246; // @[Lookup.scala 11:37:@4175.4]
  wire  _T_247; // @[Lookup.scala 11:37:@4176.4]
  wire  _T_248; // @[Lookup.scala 11:37:@4177.4]
  wire  _T_249; // @[Lookup.scala 11:37:@4178.4]
  wire  _T_250; // @[Lookup.scala 11:37:@4179.4]
  wire  _T_251; // @[Lookup.scala 11:37:@4180.4]
  wire  _T_252; // @[Lookup.scala 11:37:@4181.4]
  wire  _T_253; // @[Lookup.scala 11:37:@4182.4]
  wire  _T_254; // @[Lookup.scala 11:37:@4183.4]
  wire  _T_255; // @[Lookup.scala 11:37:@4184.4]
  wire  _T_256; // @[Lookup.scala 11:37:@4185.4]
  wire  _T_257; // @[Lookup.scala 11:37:@4186.4]
  wire  _T_258; // @[Lookup.scala 11:37:@4187.4]
  wire  _T_259; // @[Lookup.scala 11:37:@4188.4]
  wire  signals_0; // @[Lookup.scala 11:37:@4189.4]
  wire [3:0] _T_273; // @[Lookup.scala 11:37:@4203.4]
  wire [3:0] _T_274; // @[Lookup.scala 11:37:@4204.4]
  wire [3:0] _T_275; // @[Lookup.scala 11:37:@4205.4]
  wire [3:0] _T_276; // @[Lookup.scala 11:37:@4206.4]
  wire [3:0] _T_277; // @[Lookup.scala 11:37:@4207.4]
  wire [3:0] _T_278; // @[Lookup.scala 11:37:@4208.4]
  wire [3:0] _T_279; // @[Lookup.scala 11:37:@4209.4]
  wire [3:0] _T_280; // @[Lookup.scala 11:37:@4210.4]
  wire [3:0] _T_281; // @[Lookup.scala 11:37:@4211.4]
  wire [3:0] _T_282; // @[Lookup.scala 11:37:@4212.4]
  wire [3:0] _T_283; // @[Lookup.scala 11:37:@4213.4]
  wire [3:0] _T_284; // @[Lookup.scala 11:37:@4214.4]
  wire [3:0] _T_285; // @[Lookup.scala 11:37:@4215.4]
  wire [3:0] _T_286; // @[Lookup.scala 11:37:@4216.4]
  wire [3:0] _T_287; // @[Lookup.scala 11:37:@4217.4]
  wire [3:0] _T_288; // @[Lookup.scala 11:37:@4218.4]
  wire [3:0] _T_289; // @[Lookup.scala 11:37:@4219.4]
  wire [3:0] _T_290; // @[Lookup.scala 11:37:@4220.4]
  wire [3:0] _T_291; // @[Lookup.scala 11:37:@4221.4]
  wire [3:0] _T_292; // @[Lookup.scala 11:37:@4222.4]
  wire [3:0] _T_293; // @[Lookup.scala 11:37:@4223.4]
  wire [3:0] _T_294; // @[Lookup.scala 11:37:@4224.4]
  wire [3:0] _T_295; // @[Lookup.scala 11:37:@4225.4]
  wire [3:0] _T_296; // @[Lookup.scala 11:37:@4226.4]
  wire [3:0] _T_297; // @[Lookup.scala 11:37:@4227.4]
  wire [3:0] _T_298; // @[Lookup.scala 11:37:@4228.4]
  wire [3:0] _T_299; // @[Lookup.scala 11:37:@4229.4]
  wire [3:0] _T_300; // @[Lookup.scala 11:37:@4230.4]
  wire [3:0] _T_301; // @[Lookup.scala 11:37:@4231.4]
  wire [3:0] _T_302; // @[Lookup.scala 11:37:@4232.4]
  wire [3:0] _T_303; // @[Lookup.scala 11:37:@4233.4]
  wire [3:0] _T_304; // @[Lookup.scala 11:37:@4234.4]
  wire [3:0] _T_305; // @[Lookup.scala 11:37:@4235.4]
  wire [3:0] _T_306; // @[Lookup.scala 11:37:@4236.4]
  wire [3:0] _T_307; // @[Lookup.scala 11:37:@4237.4]
  wire [3:0] _T_308; // @[Lookup.scala 11:37:@4238.4]
  wire [1:0] _T_316; // @[Lookup.scala 11:37:@4247.4]
  wire [1:0] _T_317; // @[Lookup.scala 11:37:@4248.4]
  wire [1:0] _T_318; // @[Lookup.scala 11:37:@4249.4]
  wire [1:0] _T_319; // @[Lookup.scala 11:37:@4250.4]
  wire [1:0] _T_320; // @[Lookup.scala 11:37:@4251.4]
  wire [1:0] _T_321; // @[Lookup.scala 11:37:@4252.4]
  wire [1:0] _T_322; // @[Lookup.scala 11:37:@4253.4]
  wire [1:0] _T_323; // @[Lookup.scala 11:37:@4254.4]
  wire [1:0] _T_324; // @[Lookup.scala 11:37:@4255.4]
  wire [1:0] _T_325; // @[Lookup.scala 11:37:@4256.4]
  wire [1:0] _T_326; // @[Lookup.scala 11:37:@4257.4]
  wire [1:0] _T_327; // @[Lookup.scala 11:37:@4258.4]
  wire [1:0] _T_328; // @[Lookup.scala 11:37:@4259.4]
  wire [1:0] _T_329; // @[Lookup.scala 11:37:@4260.4]
  wire [1:0] _T_330; // @[Lookup.scala 11:37:@4261.4]
  wire [1:0] _T_331; // @[Lookup.scala 11:37:@4262.4]
  wire [1:0] _T_332; // @[Lookup.scala 11:37:@4263.4]
  wire [1:0] _T_333; // @[Lookup.scala 11:37:@4264.4]
  wire [1:0] _T_334; // @[Lookup.scala 11:37:@4265.4]
  wire [1:0] _T_335; // @[Lookup.scala 11:37:@4266.4]
  wire [1:0] _T_336; // @[Lookup.scala 11:37:@4267.4]
  wire [1:0] _T_337; // @[Lookup.scala 11:37:@4268.4]
  wire [1:0] _T_338; // @[Lookup.scala 11:37:@4269.4]
  wire [1:0] _T_339; // @[Lookup.scala 11:37:@4270.4]
  wire [1:0] _T_340; // @[Lookup.scala 11:37:@4271.4]
  wire [1:0] _T_341; // @[Lookup.scala 11:37:@4272.4]
  wire [1:0] _T_342; // @[Lookup.scala 11:37:@4273.4]
  wire [1:0] _T_343; // @[Lookup.scala 11:37:@4274.4]
  wire [1:0] _T_344; // @[Lookup.scala 11:37:@4275.4]
  wire [1:0] _T_345; // @[Lookup.scala 11:37:@4276.4]
  wire [1:0] _T_346; // @[Lookup.scala 11:37:@4277.4]
  wire [1:0] _T_347; // @[Lookup.scala 11:37:@4278.4]
  wire [1:0] _T_348; // @[Lookup.scala 11:37:@4279.4]
  wire [1:0] _T_349; // @[Lookup.scala 11:37:@4280.4]
  wire [1:0] _T_350; // @[Lookup.scala 11:37:@4281.4]
  wire [1:0] _T_351; // @[Lookup.scala 11:37:@4282.4]
  wire [1:0] _T_352; // @[Lookup.scala 11:37:@4283.4]
  wire [1:0] _T_353; // @[Lookup.scala 11:37:@4284.4]
  wire [1:0] _T_354; // @[Lookup.scala 11:37:@4285.4]
  wire [1:0] _T_355; // @[Lookup.scala 11:37:@4286.4]
  wire [1:0] _T_356; // @[Lookup.scala 11:37:@4287.4]
  wire [1:0] _T_357; // @[Lookup.scala 11:37:@4288.4]
  wire [2:0] _T_371; // @[Lookup.scala 11:37:@4303.4]
  wire [2:0] _T_372; // @[Lookup.scala 11:37:@4304.4]
  wire [2:0] _T_373; // @[Lookup.scala 11:37:@4305.4]
  wire [2:0] _T_374; // @[Lookup.scala 11:37:@4306.4]
  wire [2:0] _T_375; // @[Lookup.scala 11:37:@4307.4]
  wire [2:0] _T_376; // @[Lookup.scala 11:37:@4308.4]
  wire [2:0] _T_377; // @[Lookup.scala 11:37:@4309.4]
  wire [2:0] _T_378; // @[Lookup.scala 11:37:@4310.4]
  wire [2:0] _T_379; // @[Lookup.scala 11:37:@4311.4]
  wire [2:0] _T_380; // @[Lookup.scala 11:37:@4312.4]
  wire [2:0] _T_381; // @[Lookup.scala 11:37:@4313.4]
  wire [2:0] _T_382; // @[Lookup.scala 11:37:@4314.4]
  wire [2:0] _T_383; // @[Lookup.scala 11:37:@4315.4]
  wire [2:0] _T_384; // @[Lookup.scala 11:37:@4316.4]
  wire [2:0] _T_385; // @[Lookup.scala 11:37:@4317.4]
  wire [2:0] _T_386; // @[Lookup.scala 11:37:@4318.4]
  wire [2:0] _T_387; // @[Lookup.scala 11:37:@4319.4]
  wire [2:0] _T_388; // @[Lookup.scala 11:37:@4320.4]
  wire [2:0] _T_389; // @[Lookup.scala 11:37:@4321.4]
  wire [2:0] _T_390; // @[Lookup.scala 11:37:@4322.4]
  wire [2:0] _T_391; // @[Lookup.scala 11:37:@4323.4]
  wire [2:0] _T_392; // @[Lookup.scala 11:37:@4324.4]
  wire [2:0] _T_393; // @[Lookup.scala 11:37:@4325.4]
  wire [2:0] _T_394; // @[Lookup.scala 11:37:@4326.4]
  wire [2:0] _T_395; // @[Lookup.scala 11:37:@4327.4]
  wire [2:0] _T_396; // @[Lookup.scala 11:37:@4328.4]
  wire [2:0] _T_397; // @[Lookup.scala 11:37:@4329.4]
  wire [2:0] _T_398; // @[Lookup.scala 11:37:@4330.4]
  wire [2:0] _T_399; // @[Lookup.scala 11:37:@4331.4]
  wire [2:0] _T_400; // @[Lookup.scala 11:37:@4332.4]
  wire [2:0] _T_401; // @[Lookup.scala 11:37:@4333.4]
  wire [2:0] _T_402; // @[Lookup.scala 11:37:@4334.4]
  wire [2:0] _T_403; // @[Lookup.scala 11:37:@4335.4]
  wire [2:0] _T_404; // @[Lookup.scala 11:37:@4336.4]
  wire [2:0] _T_405; // @[Lookup.scala 11:37:@4337.4]
  wire [2:0] _T_406; // @[Lookup.scala 11:37:@4338.4]
  wire  _T_415; // @[Lookup.scala 11:37:@4348.4]
  wire  _T_416; // @[Lookup.scala 11:37:@4349.4]
  wire  _T_417; // @[Lookup.scala 11:37:@4350.4]
  wire  _T_418; // @[Lookup.scala 11:37:@4351.4]
  wire  _T_419; // @[Lookup.scala 11:37:@4352.4]
  wire  _T_420; // @[Lookup.scala 11:37:@4353.4]
  wire  _T_421; // @[Lookup.scala 11:37:@4354.4]
  wire  _T_422; // @[Lookup.scala 11:37:@4355.4]
  wire  _T_423; // @[Lookup.scala 11:37:@4356.4]
  wire  _T_424; // @[Lookup.scala 11:37:@4357.4]
  wire  _T_425; // @[Lookup.scala 11:37:@4358.4]
  wire  _T_426; // @[Lookup.scala 11:37:@4359.4]
  wire  _T_427; // @[Lookup.scala 11:37:@4360.4]
  wire  _T_428; // @[Lookup.scala 11:37:@4361.4]
  wire  _T_429; // @[Lookup.scala 11:37:@4362.4]
  wire  _T_430; // @[Lookup.scala 11:37:@4363.4]
  wire  _T_431; // @[Lookup.scala 11:37:@4364.4]
  wire  _T_432; // @[Lookup.scala 11:37:@4365.4]
  wire  _T_433; // @[Lookup.scala 11:37:@4366.4]
  wire  _T_434; // @[Lookup.scala 11:37:@4367.4]
  wire  _T_435; // @[Lookup.scala 11:37:@4368.4]
  wire  _T_436; // @[Lookup.scala 11:37:@4369.4]
  wire  _T_437; // @[Lookup.scala 11:37:@4370.4]
  wire  _T_438; // @[Lookup.scala 11:37:@4371.4]
  wire  _T_439; // @[Lookup.scala 11:37:@4372.4]
  wire  _T_440; // @[Lookup.scala 11:37:@4373.4]
  wire  _T_441; // @[Lookup.scala 11:37:@4374.4]
  wire  _T_442; // @[Lookup.scala 11:37:@4375.4]
  wire  _T_443; // @[Lookup.scala 11:37:@4376.4]
  wire  _T_444; // @[Lookup.scala 11:37:@4377.4]
  wire  _T_445; // @[Lookup.scala 11:37:@4378.4]
  wire  _T_446; // @[Lookup.scala 11:37:@4379.4]
  wire  _T_447; // @[Lookup.scala 11:37:@4380.4]
  wire  _T_448; // @[Lookup.scala 11:37:@4381.4]
  wire  _T_449; // @[Lookup.scala 11:37:@4382.4]
  wire  _T_450; // @[Lookup.scala 11:37:@4383.4]
  wire  _T_451; // @[Lookup.scala 11:37:@4384.4]
  wire  _T_452; // @[Lookup.scala 11:37:@4385.4]
  wire  _T_453; // @[Lookup.scala 11:37:@4386.4]
  wire  _T_454; // @[Lookup.scala 11:37:@4387.4]
  wire  _T_455; // @[Lookup.scala 11:37:@4388.4]
  wire  _T_475; // @[Lookup.scala 11:37:@4409.4]
  wire  _T_476; // @[Lookup.scala 11:37:@4410.4]
  wire  _T_477; // @[Lookup.scala 11:37:@4411.4]
  wire  _T_478; // @[Lookup.scala 11:37:@4412.4]
  wire  _T_479; // @[Lookup.scala 11:37:@4413.4]
  wire  _T_480; // @[Lookup.scala 11:37:@4414.4]
  wire  _T_481; // @[Lookup.scala 11:37:@4415.4]
  wire  _T_482; // @[Lookup.scala 11:37:@4416.4]
  wire  _T_483; // @[Lookup.scala 11:37:@4417.4]
  wire  _T_484; // @[Lookup.scala 11:37:@4418.4]
  wire  _T_485; // @[Lookup.scala 11:37:@4419.4]
  wire  _T_486; // @[Lookup.scala 11:37:@4420.4]
  wire  _T_487; // @[Lookup.scala 11:37:@4421.4]
  wire  _T_488; // @[Lookup.scala 11:37:@4422.4]
  wire  _T_489; // @[Lookup.scala 11:37:@4423.4]
  wire  _T_490; // @[Lookup.scala 11:37:@4424.4]
  wire  _T_491; // @[Lookup.scala 11:37:@4425.4]
  wire  _T_492; // @[Lookup.scala 11:37:@4426.4]
  wire  _T_493; // @[Lookup.scala 11:37:@4427.4]
  wire  _T_494; // @[Lookup.scala 11:37:@4428.4]
  wire  _T_495; // @[Lookup.scala 11:37:@4429.4]
  wire  _T_496; // @[Lookup.scala 11:37:@4430.4]
  wire  _T_497; // @[Lookup.scala 11:37:@4431.4]
  wire  _T_498; // @[Lookup.scala 11:37:@4432.4]
  wire  _T_499; // @[Lookup.scala 11:37:@4433.4]
  wire  _T_500; // @[Lookup.scala 11:37:@4434.4]
  wire  _T_501; // @[Lookup.scala 11:37:@4435.4]
  wire  _T_502; // @[Lookup.scala 11:37:@4436.4]
  wire  _T_503; // @[Lookup.scala 11:37:@4437.4]
  wire  _T_504; // @[Lookup.scala 11:37:@4438.4]
  wire [3:0] _T_512; // @[Lookup.scala 11:37:@4447.4]
  wire [3:0] _T_513; // @[Lookup.scala 11:37:@4448.4]
  wire [3:0] _T_514; // @[Lookup.scala 11:37:@4449.4]
  wire [3:0] _T_515; // @[Lookup.scala 11:37:@4450.4]
  wire [3:0] _T_516; // @[Lookup.scala 11:37:@4451.4]
  wire [3:0] _T_517; // @[Lookup.scala 11:37:@4452.4]
  wire [3:0] _T_518; // @[Lookup.scala 11:37:@4453.4]
  wire [3:0] _T_519; // @[Lookup.scala 11:37:@4454.4]
  wire [3:0] _T_520; // @[Lookup.scala 11:37:@4455.4]
  wire [3:0] _T_521; // @[Lookup.scala 11:37:@4456.4]
  wire [3:0] _T_522; // @[Lookup.scala 11:37:@4457.4]
  wire [3:0] _T_523; // @[Lookup.scala 11:37:@4458.4]
  wire [3:0] _T_524; // @[Lookup.scala 11:37:@4459.4]
  wire [3:0] _T_525; // @[Lookup.scala 11:37:@4460.4]
  wire [3:0] _T_526; // @[Lookup.scala 11:37:@4461.4]
  wire [3:0] _T_527; // @[Lookup.scala 11:37:@4462.4]
  wire [3:0] _T_528; // @[Lookup.scala 11:37:@4463.4]
  wire [3:0] _T_529; // @[Lookup.scala 11:37:@4464.4]
  wire [3:0] _T_530; // @[Lookup.scala 11:37:@4465.4]
  wire [3:0] _T_531; // @[Lookup.scala 11:37:@4466.4]
  wire [3:0] _T_532; // @[Lookup.scala 11:37:@4467.4]
  wire [3:0] _T_533; // @[Lookup.scala 11:37:@4468.4]
  wire [3:0] _T_534; // @[Lookup.scala 11:37:@4469.4]
  wire [3:0] _T_535; // @[Lookup.scala 11:37:@4470.4]
  wire [3:0] _T_536; // @[Lookup.scala 11:37:@4471.4]
  wire [3:0] _T_537; // @[Lookup.scala 11:37:@4472.4]
  wire [3:0] _T_538; // @[Lookup.scala 11:37:@4473.4]
  wire [3:0] _T_539; // @[Lookup.scala 11:37:@4474.4]
  wire [3:0] _T_540; // @[Lookup.scala 11:37:@4475.4]
  wire [3:0] _T_541; // @[Lookup.scala 11:37:@4476.4]
  wire [3:0] _T_542; // @[Lookup.scala 11:37:@4477.4]
  wire [3:0] _T_543; // @[Lookup.scala 11:37:@4478.4]
  wire [3:0] _T_544; // @[Lookup.scala 11:37:@4479.4]
  wire [3:0] _T_545; // @[Lookup.scala 11:37:@4480.4]
  wire [3:0] _T_546; // @[Lookup.scala 11:37:@4481.4]
  wire [3:0] _T_547; // @[Lookup.scala 11:37:@4482.4]
  wire [3:0] _T_548; // @[Lookup.scala 11:37:@4483.4]
  wire [3:0] _T_549; // @[Lookup.scala 11:37:@4484.4]
  wire [3:0] _T_550; // @[Lookup.scala 11:37:@4485.4]
  wire [3:0] _T_551; // @[Lookup.scala 11:37:@4486.4]
  wire [3:0] _T_552; // @[Lookup.scala 11:37:@4487.4]
  wire [3:0] _T_553; // @[Lookup.scala 11:37:@4488.4]
  wire [1:0] _T_561; // @[Lookup.scala 11:37:@4497.4]
  wire [1:0] _T_562; // @[Lookup.scala 11:37:@4498.4]
  wire [1:0] _T_563; // @[Lookup.scala 11:37:@4499.4]
  wire [1:0] _T_564; // @[Lookup.scala 11:37:@4500.4]
  wire [1:0] _T_565; // @[Lookup.scala 11:37:@4501.4]
  wire [1:0] _T_566; // @[Lookup.scala 11:37:@4502.4]
  wire [1:0] _T_567; // @[Lookup.scala 11:37:@4503.4]
  wire [1:0] _T_568; // @[Lookup.scala 11:37:@4504.4]
  wire [1:0] _T_569; // @[Lookup.scala 11:37:@4505.4]
  wire [1:0] _T_570; // @[Lookup.scala 11:37:@4506.4]
  wire [1:0] _T_571; // @[Lookup.scala 11:37:@4507.4]
  wire [1:0] _T_572; // @[Lookup.scala 11:37:@4508.4]
  wire [1:0] _T_573; // @[Lookup.scala 11:37:@4509.4]
  wire [1:0] _T_574; // @[Lookup.scala 11:37:@4510.4]
  wire [1:0] _T_575; // @[Lookup.scala 11:37:@4511.4]
  wire [1:0] _T_576; // @[Lookup.scala 11:37:@4512.4]
  wire [1:0] _T_577; // @[Lookup.scala 11:37:@4513.4]
  wire [1:0] _T_578; // @[Lookup.scala 11:37:@4514.4]
  wire [1:0] _T_579; // @[Lookup.scala 11:37:@4515.4]
  wire [1:0] _T_580; // @[Lookup.scala 11:37:@4516.4]
  wire [1:0] _T_581; // @[Lookup.scala 11:37:@4517.4]
  wire [1:0] _T_582; // @[Lookup.scala 11:37:@4518.4]
  wire [1:0] _T_583; // @[Lookup.scala 11:37:@4519.4]
  wire [1:0] _T_584; // @[Lookup.scala 11:37:@4520.4]
  wire [1:0] _T_585; // @[Lookup.scala 11:37:@4521.4]
  wire [1:0] _T_586; // @[Lookup.scala 11:37:@4522.4]
  wire [1:0] _T_587; // @[Lookup.scala 11:37:@4523.4]
  wire [1:0] _T_588; // @[Lookup.scala 11:37:@4524.4]
  wire [1:0] _T_589; // @[Lookup.scala 11:37:@4525.4]
  wire [1:0] _T_590; // @[Lookup.scala 11:37:@4526.4]
  wire [1:0] _T_591; // @[Lookup.scala 11:37:@4527.4]
  wire [1:0] _T_592; // @[Lookup.scala 11:37:@4528.4]
  wire [1:0] _T_593; // @[Lookup.scala 11:37:@4529.4]
  wire [1:0] _T_594; // @[Lookup.scala 11:37:@4530.4]
  wire [1:0] _T_595; // @[Lookup.scala 11:37:@4531.4]
  wire [1:0] _T_596; // @[Lookup.scala 11:37:@4532.4]
  wire [1:0] _T_597; // @[Lookup.scala 11:37:@4533.4]
  wire [1:0] _T_598; // @[Lookup.scala 11:37:@4534.4]
  wire [1:0] _T_599; // @[Lookup.scala 11:37:@4535.4]
  wire [1:0] _T_600; // @[Lookup.scala 11:37:@4536.4]
  wire [1:0] _T_601; // @[Lookup.scala 11:37:@4537.4]
  wire [1:0] _T_602; // @[Lookup.scala 11:37:@4538.4]
  wire  _T_616; // @[Lookup.scala 11:37:@4553.4]
  wire  _T_617; // @[Lookup.scala 11:37:@4554.4]
  wire  _T_618; // @[Lookup.scala 11:37:@4555.4]
  wire  _T_619; // @[Lookup.scala 11:37:@4556.4]
  wire  _T_620; // @[Lookup.scala 11:37:@4557.4]
  wire  _T_621; // @[Lookup.scala 11:37:@4558.4]
  wire  _T_622; // @[Lookup.scala 11:37:@4559.4]
  wire  _T_623; // @[Lookup.scala 11:37:@4560.4]
  wire  _T_624; // @[Lookup.scala 11:37:@4561.4]
  wire  _T_625; // @[Lookup.scala 11:37:@4562.4]
  wire  _T_626; // @[Lookup.scala 11:37:@4563.4]
  wire  _T_627; // @[Lookup.scala 11:37:@4564.4]
  wire  _T_628; // @[Lookup.scala 11:37:@4565.4]
  wire  _T_629; // @[Lookup.scala 11:37:@4566.4]
  wire  _T_630; // @[Lookup.scala 11:37:@4567.4]
  wire  _T_631; // @[Lookup.scala 11:37:@4568.4]
  wire  _T_632; // @[Lookup.scala 11:37:@4569.4]
  wire  _T_633; // @[Lookup.scala 11:37:@4570.4]
  wire  _T_634; // @[Lookup.scala 11:37:@4571.4]
  wire  _T_635; // @[Lookup.scala 11:37:@4572.4]
  wire  _T_636; // @[Lookup.scala 11:37:@4573.4]
  wire  _T_637; // @[Lookup.scala 11:37:@4574.4]
  wire  _T_638; // @[Lookup.scala 11:37:@4575.4]
  wire  _T_639; // @[Lookup.scala 11:37:@4576.4]
  wire  _T_640; // @[Lookup.scala 11:37:@4577.4]
  wire  _T_641; // @[Lookup.scala 11:37:@4578.4]
  wire  _T_642; // @[Lookup.scala 11:37:@4579.4]
  wire  _T_643; // @[Lookup.scala 11:37:@4580.4]
  wire  _T_644; // @[Lookup.scala 11:37:@4581.4]
  wire  _T_645; // @[Lookup.scala 11:37:@4582.4]
  wire  _T_646; // @[Lookup.scala 11:37:@4583.4]
  wire  _T_647; // @[Lookup.scala 11:37:@4584.4]
  wire  _T_648; // @[Lookup.scala 11:37:@4585.4]
  wire  _T_649; // @[Lookup.scala 11:37:@4586.4]
  wire  _T_650; // @[Lookup.scala 11:37:@4587.4]
  wire  _T_651; // @[Lookup.scala 11:37:@4588.4]
  wire  _T_653; // @[Lookup.scala 11:37:@4591.4]
  wire  _T_654; // @[Lookup.scala 11:37:@4592.4]
  wire  _T_655; // @[Lookup.scala 11:37:@4593.4]
  wire  _T_656; // @[Lookup.scala 11:37:@4594.4]
  wire  _T_657; // @[Lookup.scala 11:37:@4595.4]
  wire  _T_658; // @[Lookup.scala 11:37:@4596.4]
  wire  _T_659; // @[Lookup.scala 11:37:@4597.4]
  wire  _T_660; // @[Lookup.scala 11:37:@4598.4]
  wire  _T_661; // @[Lookup.scala 11:37:@4599.4]
  wire  _T_662; // @[Lookup.scala 11:37:@4600.4]
  wire  _T_663; // @[Lookup.scala 11:37:@4601.4]
  wire  _T_664; // @[Lookup.scala 11:37:@4602.4]
  wire  _T_665; // @[Lookup.scala 11:37:@4603.4]
  wire  _T_666; // @[Lookup.scala 11:37:@4604.4]
  wire  _T_667; // @[Lookup.scala 11:37:@4605.4]
  wire  _T_668; // @[Lookup.scala 11:37:@4606.4]
  wire  _T_669; // @[Lookup.scala 11:37:@4607.4]
  wire  _T_670; // @[Lookup.scala 11:37:@4608.4]
  wire  _T_671; // @[Lookup.scala 11:37:@4609.4]
  wire  _T_672; // @[Lookup.scala 11:37:@4610.4]
  wire  _T_673; // @[Lookup.scala 11:37:@4611.4]
  wire  _T_674; // @[Lookup.scala 11:37:@4612.4]
  wire  _T_675; // @[Lookup.scala 11:37:@4613.4]
  wire  _T_676; // @[Lookup.scala 11:37:@4614.4]
  wire  _T_677; // @[Lookup.scala 11:37:@4615.4]
  wire  _T_678; // @[Lookup.scala 11:37:@4616.4]
  wire  _T_679; // @[Lookup.scala 11:37:@4617.4]
  wire  _T_680; // @[Lookup.scala 11:37:@4618.4]
  wire  _T_681; // @[Lookup.scala 11:37:@4619.4]
  wire  _T_682; // @[Lookup.scala 11:37:@4620.4]
  wire  _T_683; // @[Lookup.scala 11:37:@4621.4]
  wire  _T_684; // @[Lookup.scala 11:37:@4622.4]
  wire  _T_685; // @[Lookup.scala 11:37:@4623.4]
  wire  _T_686; // @[Lookup.scala 11:37:@4624.4]
  wire  _T_687; // @[Lookup.scala 11:37:@4625.4]
  wire  _T_688; // @[Lookup.scala 11:37:@4626.4]
  wire  _T_689; // @[Lookup.scala 11:37:@4627.4]
  wire  _T_690; // @[Lookup.scala 11:37:@4628.4]
  wire  _T_691; // @[Lookup.scala 11:37:@4629.4]
  wire  _T_692; // @[Lookup.scala 11:37:@4630.4]
  wire  _T_693; // @[Lookup.scala 11:37:@4631.4]
  wire  _T_694; // @[Lookup.scala 11:37:@4632.4]
  wire  _T_695; // @[Lookup.scala 11:37:@4633.4]
  wire  _T_696; // @[Lookup.scala 11:37:@4634.4]
  wire  _T_697; // @[Lookup.scala 11:37:@4635.4]
  wire  _T_698; // @[Lookup.scala 11:37:@4636.4]
  wire  _T_699; // @[Lookup.scala 11:37:@4637.4]
  wire  _T_700; // @[Lookup.scala 11:37:@4638.4]
  wire  _T_744; // @[Lookup.scala 11:37:@4683.4]
  wire  _T_745; // @[Lookup.scala 11:37:@4684.4]
  wire  _T_746; // @[Lookup.scala 11:37:@4685.4]
  wire  _T_747; // @[Lookup.scala 11:37:@4686.4]
  wire  _T_748; // @[Lookup.scala 11:37:@4687.4]
  wire  _T_749; // @[Lookup.scala 11:37:@4688.4]
  wire [2:0] _T_792; // @[Lookup.scala 11:37:@4732.4]
  wire [2:0] _T_793; // @[Lookup.scala 11:37:@4733.4]
  wire [2:0] _T_794; // @[Lookup.scala 11:37:@4734.4]
  wire [2:0] _T_795; // @[Lookup.scala 11:37:@4735.4]
  wire [2:0] _T_796; // @[Lookup.scala 11:37:@4736.4]
  wire [2:0] _T_797; // @[Lookup.scala 11:37:@4737.4]
  wire [2:0] _T_798; // @[Lookup.scala 11:37:@4738.4]
  wire [2:0] _T_802; // @[Lookup.scala 11:37:@4743.4]
  wire [2:0] _T_803; // @[Lookup.scala 11:37:@4744.4]
  wire [2:0] _T_804; // @[Lookup.scala 11:37:@4745.4]
  wire [2:0] _T_805; // @[Lookup.scala 11:37:@4746.4]
  wire [2:0] _T_806; // @[Lookup.scala 11:37:@4747.4]
  wire [2:0] _T_807; // @[Lookup.scala 11:37:@4748.4]
  wire [2:0] _T_808; // @[Lookup.scala 11:37:@4749.4]
  wire [2:0] _T_809; // @[Lookup.scala 11:37:@4750.4]
  wire [2:0] _T_810; // @[Lookup.scala 11:37:@4751.4]
  wire [2:0] _T_811; // @[Lookup.scala 11:37:@4752.4]
  wire [2:0] _T_812; // @[Lookup.scala 11:37:@4753.4]
  wire [2:0] _T_813; // @[Lookup.scala 11:37:@4754.4]
  wire [2:0] _T_814; // @[Lookup.scala 11:37:@4755.4]
  wire [2:0] _T_815; // @[Lookup.scala 11:37:@4756.4]
  wire [2:0] _T_816; // @[Lookup.scala 11:37:@4757.4]
  wire [2:0] _T_817; // @[Lookup.scala 11:37:@4758.4]
  wire [2:0] _T_818; // @[Lookup.scala 11:37:@4759.4]
  wire [2:0] _T_819; // @[Lookup.scala 11:37:@4760.4]
  wire [2:0] _T_820; // @[Lookup.scala 11:37:@4761.4]
  wire [2:0] _T_821; // @[Lookup.scala 11:37:@4762.4]
  wire [2:0] _T_822; // @[Lookup.scala 11:37:@4763.4]
  wire [2:0] _T_823; // @[Lookup.scala 11:37:@4764.4]
  wire [2:0] _T_824; // @[Lookup.scala 11:37:@4765.4]
  wire [2:0] _T_825; // @[Lookup.scala 11:37:@4766.4]
  wire [2:0] _T_826; // @[Lookup.scala 11:37:@4767.4]
  wire [2:0] _T_827; // @[Lookup.scala 11:37:@4768.4]
  wire [2:0] _T_828; // @[Lookup.scala 11:37:@4769.4]
  wire [2:0] _T_829; // @[Lookup.scala 11:37:@4770.4]
  wire [2:0] _T_830; // @[Lookup.scala 11:37:@4771.4]
  wire [2:0] _T_831; // @[Lookup.scala 11:37:@4772.4]
  wire [2:0] _T_832; // @[Lookup.scala 11:37:@4773.4]
  wire [2:0] _T_833; // @[Lookup.scala 11:37:@4774.4]
  wire [2:0] _T_834; // @[Lookup.scala 11:37:@4775.4]
  wire [2:0] _T_835; // @[Lookup.scala 11:37:@4776.4]
  wire [2:0] _T_836; // @[Lookup.scala 11:37:@4777.4]
  wire [2:0] _T_837; // @[Lookup.scala 11:37:@4778.4]
  wire [2:0] _T_838; // @[Lookup.scala 11:37:@4779.4]
  wire [2:0] _T_839; // @[Lookup.scala 11:37:@4780.4]
  wire [2:0] _T_840; // @[Lookup.scala 11:37:@4781.4]
  wire [2:0] _T_841; // @[Lookup.scala 11:37:@4782.4]
  wire [2:0] _T_842; // @[Lookup.scala 11:37:@4783.4]
  wire [2:0] _T_843; // @[Lookup.scala 11:37:@4784.4]
  wire [2:0] _T_844; // @[Lookup.scala 11:37:@4785.4]
  wire [2:0] _T_845; // @[Lookup.scala 11:37:@4786.4]
  wire [2:0] _T_846; // @[Lookup.scala 11:37:@4787.4]
  wire [2:0] _T_847; // @[Lookup.scala 11:37:@4788.4]
  wire  _T_850; // @[Lookup.scala 11:37:@4792.4]
  wire  _T_851; // @[Lookup.scala 11:37:@4793.4]
  wire  _T_852; // @[Lookup.scala 11:37:@4794.4]
  wire  _T_853; // @[Lookup.scala 11:37:@4795.4]
  wire  _T_854; // @[Lookup.scala 11:37:@4796.4]
  wire  _T_855; // @[Lookup.scala 11:37:@4797.4]
  wire  _T_856; // @[Lookup.scala 11:37:@4798.4]
  wire  _T_857; // @[Lookup.scala 11:37:@4799.4]
  wire  _T_858; // @[Lookup.scala 11:37:@4800.4]
  wire  _T_859; // @[Lookup.scala 11:37:@4801.4]
  wire  _T_860; // @[Lookup.scala 11:37:@4802.4]
  wire  _T_861; // @[Lookup.scala 11:37:@4803.4]
  wire  _T_862; // @[Lookup.scala 11:37:@4804.4]
  wire  _T_863; // @[Lookup.scala 11:37:@4805.4]
  wire  _T_864; // @[Lookup.scala 11:37:@4806.4]
  wire  _T_865; // @[Lookup.scala 11:37:@4807.4]
  wire  _T_866; // @[Lookup.scala 11:37:@4808.4]
  wire  _T_867; // @[Lookup.scala 11:37:@4809.4]
  wire  _T_868; // @[Lookup.scala 11:37:@4810.4]
  wire  _T_869; // @[Lookup.scala 11:37:@4811.4]
  wire  _T_870; // @[Lookup.scala 11:37:@4812.4]
  wire  _T_871; // @[Lookup.scala 11:37:@4813.4]
  wire  _T_872; // @[Lookup.scala 11:37:@4814.4]
  wire  _T_873; // @[Lookup.scala 11:37:@4815.4]
  wire  _T_874; // @[Lookup.scala 11:37:@4816.4]
  wire  _T_875; // @[Lookup.scala 11:37:@4817.4]
  wire  _T_876; // @[Lookup.scala 11:37:@4818.4]
  wire  _T_877; // @[Lookup.scala 11:37:@4819.4]
  wire  _T_878; // @[Lookup.scala 11:37:@4820.4]
  wire  _T_879; // @[Lookup.scala 11:37:@4821.4]
  wire  _T_880; // @[Lookup.scala 11:37:@4822.4]
  wire  _T_881; // @[Lookup.scala 11:37:@4823.4]
  wire  _T_882; // @[Lookup.scala 11:37:@4824.4]
  wire  _T_883; // @[Lookup.scala 11:37:@4825.4]
  wire  _T_884; // @[Lookup.scala 11:37:@4826.4]
  wire  _T_885; // @[Lookup.scala 11:37:@4827.4]
  wire  _T_886; // @[Lookup.scala 11:37:@4828.4]
  wire  _T_887; // @[Lookup.scala 11:37:@4829.4]
  wire  _T_888; // @[Lookup.scala 11:37:@4830.4]
  wire  _T_889; // @[Lookup.scala 11:37:@4831.4]
  wire  _T_890; // @[Lookup.scala 11:37:@4832.4]
  wire  _T_891; // @[Lookup.scala 11:37:@4833.4]
  wire  _T_892; // @[Lookup.scala 11:37:@4834.4]
  wire  _T_893; // @[Lookup.scala 11:37:@4835.4]
  wire  _T_894; // @[Lookup.scala 11:37:@4836.4]
  wire  _T_895; // @[Lookup.scala 11:37:@4837.4]
  wire  _T_896; // @[Lookup.scala 11:37:@4838.4]
  wire [4:0] _T_899; // @[InstDecoder.scala 130:31:@4855.4]
  wire [4:0] _T_901; // @[InstDecoder.scala 132:31:@4859.4]
  wire [4:0] func; // @[InstDecoder.scala 134:21:@4861.4]
  wire  _T_905; // @[InstDecoder.scala 136:38:@4864.4]
  wire  _T_907; // @[InstDecoder.scala 137:39:@4865.4]
  wire  _T_908; // @[InstDecoder.scala 141:32:@4866.4]
  wire  _T_910; // @[InstDecoder.scala 135:37:@4867.4]
  wire  _T_912; // @[InstDecoder.scala 135:53:@4868.4]
  wire  _T_913; // @[InstDecoder.scala 135:45:@4869.4]
  wire [4:0] _GEN_0; // @[InstDecoder.scala 142:24:@4873.4]
  wire  _T_917; // @[InstDecoder.scala 142:24:@4873.4]
  wire  _T_919; // @[InstDecoder.scala 135:37:@4874.4]
  wire  _T_921; // @[InstDecoder.scala 135:53:@4875.4]
  wire  _T_922; // @[InstDecoder.scala 135:45:@4876.4]
  wire  _T_923; // @[InstDecoder.scala 142:41:@4877.4]
  wire  _T_930; // @[InstDecoder.scala 143:6:@4881.4]
  wire  _T_931; // @[InstDecoder.scala 143:50:@4882.4]
  wire  _T_932; // @[InstDecoder.scala 143:29:@4883.4]
  wire [11:0] imm_itype; // @[InstDecoder.scala 146:27:@4886.4]
  wire [6:0] _T_934; // @[InstDecoder.scala 147:31:@4887.4]
  wire [11:0] imm_stype; // @[Cat.scala 30:58:@4889.4]
  wire  _T_936; // @[InstDecoder.scala 148:31:@4890.4]
  wire  _T_937; // @[InstDecoder.scala 148:44:@4891.4]
  wire [5:0] _T_938; // @[InstDecoder.scala 148:56:@4892.4]
  wire [3:0] _T_939; // @[InstDecoder.scala 148:73:@4893.4]
  wire [11:0] imm_sbtype; // @[Cat.scala 30:58:@4896.4]
  wire [19:0] imm_utype; // @[InstDecoder.scala 149:27:@4897.4]
  wire [7:0] _T_943; // @[InstDecoder.scala 150:44:@4899.4]
  wire  _T_944; // @[InstDecoder.scala 150:60:@4900.4]
  wire [9:0] _T_945; // @[InstDecoder.scala 150:73:@4901.4]
  wire [19:0] imm_ujtype; // @[Cat.scala 30:58:@4904.4]
  wire  _T_948; // @[InstDecoder.scala 153:43:@4905.4]
  wire [19:0] _T_952; // @[Bitwise.scala 72:12:@4907.4]
  wire  _T_954; // @[InstDecoder.scala 154:43:@4910.4]
  wire [19:0] _T_958; // @[Bitwise.scala 72:12:@4912.4]
  wire  _T_960; // @[InstDecoder.scala 155:44:@4915.4]
  wire [18:0] _T_964; // @[Bitwise.scala 72:12:@4917.4]
  wire [30:0] _T_966; // @[Cat.scala 30:58:@4918.4]
  wire  _T_974; // @[InstDecoder.scala 157:44:@4924.4]
  wire [10:0] _T_978; // @[Bitwise.scala 72:12:@4926.4]
  wire [30:0] _T_980; // @[Cat.scala 30:58:@4927.4]
  assign _T_13 = io_inst & 32'h707f; // @[Lookup.scala 9:38:@4040.4]
  assign _T_14 = 32'h2003 == _T_13; // @[Lookup.scala 9:38:@4041.4]
  assign _T_18 = 32'h3 == _T_13; // @[Lookup.scala 9:38:@4043.4]
  assign _T_22 = 32'h4003 == _T_13; // @[Lookup.scala 9:38:@4045.4]
  assign _T_26 = 32'h1003 == _T_13; // @[Lookup.scala 9:38:@4047.4]
  assign _T_30 = 32'h5003 == _T_13; // @[Lookup.scala 9:38:@4049.4]
  assign _T_34 = 32'h2023 == _T_13; // @[Lookup.scala 9:38:@4051.4]
  assign _T_38 = 32'h23 == _T_13; // @[Lookup.scala 9:38:@4053.4]
  assign _T_42 = 32'h1023 == _T_13; // @[Lookup.scala 9:38:@4055.4]
  assign _T_45 = io_inst & 32'h7f; // @[Lookup.scala 9:38:@4056.4]
  assign _T_46 = 32'h17 == _T_45; // @[Lookup.scala 9:38:@4057.4]
  assign _T_50 = 32'h37 == _T_45; // @[Lookup.scala 9:38:@4059.4]
  assign _T_54 = 32'h13 == _T_13; // @[Lookup.scala 9:38:@4061.4]
  assign _T_58 = 32'h7013 == _T_13; // @[Lookup.scala 9:38:@4063.4]
  assign _T_62 = 32'h6013 == _T_13; // @[Lookup.scala 9:38:@4065.4]
  assign _T_66 = 32'h4013 == _T_13; // @[Lookup.scala 9:38:@4067.4]
  assign _T_70 = 32'h2013 == _T_13; // @[Lookup.scala 9:38:@4069.4]
  assign _T_74 = 32'h3013 == _T_13; // @[Lookup.scala 9:38:@4071.4]
  assign _T_77 = io_inst & 32'hfc00707f; // @[Lookup.scala 9:38:@4072.4]
  assign _T_78 = 32'h1013 == _T_77; // @[Lookup.scala 9:38:@4073.4]
  assign _T_82 = 32'h40005013 == _T_77; // @[Lookup.scala 9:38:@4075.4]
  assign _T_86 = 32'h5013 == _T_77; // @[Lookup.scala 9:38:@4077.4]
  assign _T_89 = io_inst & 32'hfe00707f; // @[Lookup.scala 9:38:@4078.4]
  assign _T_90 = 32'h1033 == _T_89; // @[Lookup.scala 9:38:@4079.4]
  assign _T_94 = 32'h33 == _T_89; // @[Lookup.scala 9:38:@4081.4]
  assign _T_98 = 32'h40000033 == _T_89; // @[Lookup.scala 9:38:@4083.4]
  assign _T_102 = 32'h2033 == _T_89; // @[Lookup.scala 9:38:@4085.4]
  assign _T_106 = 32'h3033 == _T_89; // @[Lookup.scala 9:38:@4087.4]
  assign _T_110 = 32'h7033 == _T_89; // @[Lookup.scala 9:38:@4089.4]
  assign _T_114 = 32'h6033 == _T_89; // @[Lookup.scala 9:38:@4091.4]
  assign _T_118 = 32'h4033 == _T_89; // @[Lookup.scala 9:38:@4093.4]
  assign _T_122 = 32'h40005033 == _T_89; // @[Lookup.scala 9:38:@4095.4]
  assign _T_126 = 32'h5033 == _T_89; // @[Lookup.scala 9:38:@4097.4]
  assign _T_130 = 32'h6f == _T_45; // @[Lookup.scala 9:38:@4099.4]
  assign _T_134 = 32'h67 == _T_13; // @[Lookup.scala 9:38:@4101.4]
  assign _T_138 = 32'h63 == _T_13; // @[Lookup.scala 9:38:@4103.4]
  assign _T_142 = 32'h1063 == _T_13; // @[Lookup.scala 9:38:@4105.4]
  assign _T_146 = 32'h5063 == _T_13; // @[Lookup.scala 9:38:@4107.4]
  assign _T_150 = 32'h7063 == _T_13; // @[Lookup.scala 9:38:@4109.4]
  assign _T_154 = 32'h4063 == _T_13; // @[Lookup.scala 9:38:@4111.4]
  assign _T_158 = 32'h6063 == _T_13; // @[Lookup.scala 9:38:@4113.4]
  assign _T_162 = 32'h5073 == _T_13; // @[Lookup.scala 9:38:@4115.4]
  assign _T_166 = 32'h6073 == _T_13; // @[Lookup.scala 9:38:@4117.4]
  assign _T_170 = 32'h1073 == _T_13; // @[Lookup.scala 9:38:@4119.4]
  assign _T_174 = 32'h2073 == _T_13; // @[Lookup.scala 9:38:@4121.4]
  assign _T_178 = 32'h3073 == _T_13; // @[Lookup.scala 9:38:@4123.4]
  assign _T_182 = 32'h7073 == _T_13; // @[Lookup.scala 9:38:@4125.4]
  assign _T_186 = 32'h73 == io_inst; // @[Lookup.scala 9:38:@4127.4]
  assign _T_190 = 32'h30200073 == io_inst; // @[Lookup.scala 9:38:@4129.4]
  assign _T_194 = 32'h7b200073 == io_inst; // @[Lookup.scala 9:38:@4131.4]
  assign _T_198 = 32'h100073 == io_inst; // @[Lookup.scala 9:38:@4133.4]
  assign _T_202 = 32'h10500073 == io_inst; // @[Lookup.scala 9:38:@4135.4]
  assign _T_206 = 32'h100f == _T_13; // @[Lookup.scala 9:38:@4137.4]
  assign _T_210 = 32'hf == _T_13; // @[Lookup.scala 9:38:@4139.4]
  assign _T_212 = _T_206 ? 1'h1 : _T_210; // @[Lookup.scala 11:37:@4141.4]
  assign _T_213 = _T_202 ? 1'h1 : _T_212; // @[Lookup.scala 11:37:@4142.4]
  assign _T_214 = _T_198 ? 1'h1 : _T_213; // @[Lookup.scala 11:37:@4143.4]
  assign _T_215 = _T_194 ? 1'h1 : _T_214; // @[Lookup.scala 11:37:@4144.4]
  assign _T_216 = _T_190 ? 1'h1 : _T_215; // @[Lookup.scala 11:37:@4145.4]
  assign _T_217 = _T_186 ? 1'h1 : _T_216; // @[Lookup.scala 11:37:@4146.4]
  assign _T_218 = _T_182 ? 1'h1 : _T_217; // @[Lookup.scala 11:37:@4147.4]
  assign _T_219 = _T_178 ? 1'h1 : _T_218; // @[Lookup.scala 11:37:@4148.4]
  assign _T_220 = _T_174 ? 1'h1 : _T_219; // @[Lookup.scala 11:37:@4149.4]
  assign _T_221 = _T_170 ? 1'h1 : _T_220; // @[Lookup.scala 11:37:@4150.4]
  assign _T_222 = _T_166 ? 1'h1 : _T_221; // @[Lookup.scala 11:37:@4151.4]
  assign _T_223 = _T_162 ? 1'h1 : _T_222; // @[Lookup.scala 11:37:@4152.4]
  assign _T_224 = _T_158 ? 1'h1 : _T_223; // @[Lookup.scala 11:37:@4153.4]
  assign _T_225 = _T_154 ? 1'h1 : _T_224; // @[Lookup.scala 11:37:@4154.4]
  assign _T_226 = _T_150 ? 1'h1 : _T_225; // @[Lookup.scala 11:37:@4155.4]
  assign _T_227 = _T_146 ? 1'h1 : _T_226; // @[Lookup.scala 11:37:@4156.4]
  assign _T_228 = _T_142 ? 1'h1 : _T_227; // @[Lookup.scala 11:37:@4157.4]
  assign _T_229 = _T_138 ? 1'h1 : _T_228; // @[Lookup.scala 11:37:@4158.4]
  assign _T_230 = _T_134 ? 1'h1 : _T_229; // @[Lookup.scala 11:37:@4159.4]
  assign _T_231 = _T_130 ? 1'h1 : _T_230; // @[Lookup.scala 11:37:@4160.4]
  assign _T_232 = _T_126 ? 1'h1 : _T_231; // @[Lookup.scala 11:37:@4161.4]
  assign _T_233 = _T_122 ? 1'h1 : _T_232; // @[Lookup.scala 11:37:@4162.4]
  assign _T_234 = _T_118 ? 1'h1 : _T_233; // @[Lookup.scala 11:37:@4163.4]
  assign _T_235 = _T_114 ? 1'h1 : _T_234; // @[Lookup.scala 11:37:@4164.4]
  assign _T_236 = _T_110 ? 1'h1 : _T_235; // @[Lookup.scala 11:37:@4165.4]
  assign _T_237 = _T_106 ? 1'h1 : _T_236; // @[Lookup.scala 11:37:@4166.4]
  assign _T_238 = _T_102 ? 1'h1 : _T_237; // @[Lookup.scala 11:37:@4167.4]
  assign _T_239 = _T_98 ? 1'h1 : _T_238; // @[Lookup.scala 11:37:@4168.4]
  assign _T_240 = _T_94 ? 1'h1 : _T_239; // @[Lookup.scala 11:37:@4169.4]
  assign _T_241 = _T_90 ? 1'h1 : _T_240; // @[Lookup.scala 11:37:@4170.4]
  assign _T_242 = _T_86 ? 1'h1 : _T_241; // @[Lookup.scala 11:37:@4171.4]
  assign _T_243 = _T_82 ? 1'h1 : _T_242; // @[Lookup.scala 11:37:@4172.4]
  assign _T_244 = _T_78 ? 1'h1 : _T_243; // @[Lookup.scala 11:37:@4173.4]
  assign _T_245 = _T_74 ? 1'h1 : _T_244; // @[Lookup.scala 11:37:@4174.4]
  assign _T_246 = _T_70 ? 1'h1 : _T_245; // @[Lookup.scala 11:37:@4175.4]
  assign _T_247 = _T_66 ? 1'h1 : _T_246; // @[Lookup.scala 11:37:@4176.4]
  assign _T_248 = _T_62 ? 1'h1 : _T_247; // @[Lookup.scala 11:37:@4177.4]
  assign _T_249 = _T_58 ? 1'h1 : _T_248; // @[Lookup.scala 11:37:@4178.4]
  assign _T_250 = _T_54 ? 1'h1 : _T_249; // @[Lookup.scala 11:37:@4179.4]
  assign _T_251 = _T_50 ? 1'h1 : _T_250; // @[Lookup.scala 11:37:@4180.4]
  assign _T_252 = _T_46 ? 1'h1 : _T_251; // @[Lookup.scala 11:37:@4181.4]
  assign _T_253 = _T_42 ? 1'h1 : _T_252; // @[Lookup.scala 11:37:@4182.4]
  assign _T_254 = _T_38 ? 1'h1 : _T_253; // @[Lookup.scala 11:37:@4183.4]
  assign _T_255 = _T_34 ? 1'h1 : _T_254; // @[Lookup.scala 11:37:@4184.4]
  assign _T_256 = _T_30 ? 1'h1 : _T_255; // @[Lookup.scala 11:37:@4185.4]
  assign _T_257 = _T_26 ? 1'h1 : _T_256; // @[Lookup.scala 11:37:@4186.4]
  assign _T_258 = _T_22 ? 1'h1 : _T_257; // @[Lookup.scala 11:37:@4187.4]
  assign _T_259 = _T_18 ? 1'h1 : _T_258; // @[Lookup.scala 11:37:@4188.4]
  assign signals_0 = _T_14 ? 1'h1 : _T_259; // @[Lookup.scala 11:37:@4189.4]
  assign _T_273 = _T_158 ? 4'h6 : 4'h0; // @[Lookup.scala 11:37:@4203.4]
  assign _T_274 = _T_154 ? 4'h5 : _T_273; // @[Lookup.scala 11:37:@4204.4]
  assign _T_275 = _T_150 ? 4'h4 : _T_274; // @[Lookup.scala 11:37:@4205.4]
  assign _T_276 = _T_146 ? 4'h3 : _T_275; // @[Lookup.scala 11:37:@4206.4]
  assign _T_277 = _T_142 ? 4'h1 : _T_276; // @[Lookup.scala 11:37:@4207.4]
  assign _T_278 = _T_138 ? 4'h2 : _T_277; // @[Lookup.scala 11:37:@4208.4]
  assign _T_279 = _T_134 ? 4'h8 : _T_278; // @[Lookup.scala 11:37:@4209.4]
  assign _T_280 = _T_130 ? 4'h7 : _T_279; // @[Lookup.scala 11:37:@4210.4]
  assign _T_281 = _T_126 ? 4'h0 : _T_280; // @[Lookup.scala 11:37:@4211.4]
  assign _T_282 = _T_122 ? 4'h0 : _T_281; // @[Lookup.scala 11:37:@4212.4]
  assign _T_283 = _T_118 ? 4'h0 : _T_282; // @[Lookup.scala 11:37:@4213.4]
  assign _T_284 = _T_114 ? 4'h0 : _T_283; // @[Lookup.scala 11:37:@4214.4]
  assign _T_285 = _T_110 ? 4'h0 : _T_284; // @[Lookup.scala 11:37:@4215.4]
  assign _T_286 = _T_106 ? 4'h0 : _T_285; // @[Lookup.scala 11:37:@4216.4]
  assign _T_287 = _T_102 ? 4'h0 : _T_286; // @[Lookup.scala 11:37:@4217.4]
  assign _T_288 = _T_98 ? 4'h0 : _T_287; // @[Lookup.scala 11:37:@4218.4]
  assign _T_289 = _T_94 ? 4'h0 : _T_288; // @[Lookup.scala 11:37:@4219.4]
  assign _T_290 = _T_90 ? 4'h0 : _T_289; // @[Lookup.scala 11:37:@4220.4]
  assign _T_291 = _T_86 ? 4'h0 : _T_290; // @[Lookup.scala 11:37:@4221.4]
  assign _T_292 = _T_82 ? 4'h0 : _T_291; // @[Lookup.scala 11:37:@4222.4]
  assign _T_293 = _T_78 ? 4'h0 : _T_292; // @[Lookup.scala 11:37:@4223.4]
  assign _T_294 = _T_74 ? 4'h0 : _T_293; // @[Lookup.scala 11:37:@4224.4]
  assign _T_295 = _T_70 ? 4'h0 : _T_294; // @[Lookup.scala 11:37:@4225.4]
  assign _T_296 = _T_66 ? 4'h0 : _T_295; // @[Lookup.scala 11:37:@4226.4]
  assign _T_297 = _T_62 ? 4'h0 : _T_296; // @[Lookup.scala 11:37:@4227.4]
  assign _T_298 = _T_58 ? 4'h0 : _T_297; // @[Lookup.scala 11:37:@4228.4]
  assign _T_299 = _T_54 ? 4'h0 : _T_298; // @[Lookup.scala 11:37:@4229.4]
  assign _T_300 = _T_50 ? 4'h0 : _T_299; // @[Lookup.scala 11:37:@4230.4]
  assign _T_301 = _T_46 ? 4'h0 : _T_300; // @[Lookup.scala 11:37:@4231.4]
  assign _T_302 = _T_42 ? 4'h0 : _T_301; // @[Lookup.scala 11:37:@4232.4]
  assign _T_303 = _T_38 ? 4'h0 : _T_302; // @[Lookup.scala 11:37:@4233.4]
  assign _T_304 = _T_34 ? 4'h0 : _T_303; // @[Lookup.scala 11:37:@4234.4]
  assign _T_305 = _T_30 ? 4'h0 : _T_304; // @[Lookup.scala 11:37:@4235.4]
  assign _T_306 = _T_26 ? 4'h0 : _T_305; // @[Lookup.scala 11:37:@4236.4]
  assign _T_307 = _T_22 ? 4'h0 : _T_306; // @[Lookup.scala 11:37:@4237.4]
  assign _T_308 = _T_18 ? 4'h0 : _T_307; // @[Lookup.scala 11:37:@4238.4]
  assign _T_316 = _T_182 ? 2'h2 : 2'h0; // @[Lookup.scala 11:37:@4247.4]
  assign _T_317 = _T_178 ? 2'h0 : _T_316; // @[Lookup.scala 11:37:@4248.4]
  assign _T_318 = _T_174 ? 2'h0 : _T_317; // @[Lookup.scala 11:37:@4249.4]
  assign _T_319 = _T_170 ? 2'h0 : _T_318; // @[Lookup.scala 11:37:@4250.4]
  assign _T_320 = _T_166 ? 2'h2 : _T_319; // @[Lookup.scala 11:37:@4251.4]
  assign _T_321 = _T_162 ? 2'h2 : _T_320; // @[Lookup.scala 11:37:@4252.4]
  assign _T_322 = _T_158 ? 2'h0 : _T_321; // @[Lookup.scala 11:37:@4253.4]
  assign _T_323 = _T_154 ? 2'h0 : _T_322; // @[Lookup.scala 11:37:@4254.4]
  assign _T_324 = _T_150 ? 2'h0 : _T_323; // @[Lookup.scala 11:37:@4255.4]
  assign _T_325 = _T_146 ? 2'h0 : _T_324; // @[Lookup.scala 11:37:@4256.4]
  assign _T_326 = _T_142 ? 2'h0 : _T_325; // @[Lookup.scala 11:37:@4257.4]
  assign _T_327 = _T_138 ? 2'h0 : _T_326; // @[Lookup.scala 11:37:@4258.4]
  assign _T_328 = _T_134 ? 2'h0 : _T_327; // @[Lookup.scala 11:37:@4259.4]
  assign _T_329 = _T_130 ? 2'h0 : _T_328; // @[Lookup.scala 11:37:@4260.4]
  assign _T_330 = _T_126 ? 2'h0 : _T_329; // @[Lookup.scala 11:37:@4261.4]
  assign _T_331 = _T_122 ? 2'h0 : _T_330; // @[Lookup.scala 11:37:@4262.4]
  assign _T_332 = _T_118 ? 2'h0 : _T_331; // @[Lookup.scala 11:37:@4263.4]
  assign _T_333 = _T_114 ? 2'h0 : _T_332; // @[Lookup.scala 11:37:@4264.4]
  assign _T_334 = _T_110 ? 2'h0 : _T_333; // @[Lookup.scala 11:37:@4265.4]
  assign _T_335 = _T_106 ? 2'h0 : _T_334; // @[Lookup.scala 11:37:@4266.4]
  assign _T_336 = _T_102 ? 2'h0 : _T_335; // @[Lookup.scala 11:37:@4267.4]
  assign _T_337 = _T_98 ? 2'h0 : _T_336; // @[Lookup.scala 11:37:@4268.4]
  assign _T_338 = _T_94 ? 2'h0 : _T_337; // @[Lookup.scala 11:37:@4269.4]
  assign _T_339 = _T_90 ? 2'h0 : _T_338; // @[Lookup.scala 11:37:@4270.4]
  assign _T_340 = _T_86 ? 2'h0 : _T_339; // @[Lookup.scala 11:37:@4271.4]
  assign _T_341 = _T_82 ? 2'h0 : _T_340; // @[Lookup.scala 11:37:@4272.4]
  assign _T_342 = _T_78 ? 2'h0 : _T_341; // @[Lookup.scala 11:37:@4273.4]
  assign _T_343 = _T_74 ? 2'h0 : _T_342; // @[Lookup.scala 11:37:@4274.4]
  assign _T_344 = _T_70 ? 2'h0 : _T_343; // @[Lookup.scala 11:37:@4275.4]
  assign _T_345 = _T_66 ? 2'h0 : _T_344; // @[Lookup.scala 11:37:@4276.4]
  assign _T_346 = _T_62 ? 2'h0 : _T_345; // @[Lookup.scala 11:37:@4277.4]
  assign _T_347 = _T_58 ? 2'h0 : _T_346; // @[Lookup.scala 11:37:@4278.4]
  assign _T_348 = _T_54 ? 2'h0 : _T_347; // @[Lookup.scala 11:37:@4279.4]
  assign _T_349 = _T_50 ? 2'h0 : _T_348; // @[Lookup.scala 11:37:@4280.4]
  assign _T_350 = _T_46 ? 2'h1 : _T_349; // @[Lookup.scala 11:37:@4281.4]
  assign _T_351 = _T_42 ? 2'h0 : _T_350; // @[Lookup.scala 11:37:@4282.4]
  assign _T_352 = _T_38 ? 2'h0 : _T_351; // @[Lookup.scala 11:37:@4283.4]
  assign _T_353 = _T_34 ? 2'h0 : _T_352; // @[Lookup.scala 11:37:@4284.4]
  assign _T_354 = _T_30 ? 2'h0 : _T_353; // @[Lookup.scala 11:37:@4285.4]
  assign _T_355 = _T_26 ? 2'h0 : _T_354; // @[Lookup.scala 11:37:@4286.4]
  assign _T_356 = _T_22 ? 2'h0 : _T_355; // @[Lookup.scala 11:37:@4287.4]
  assign _T_357 = _T_18 ? 2'h0 : _T_356; // @[Lookup.scala 11:37:@4288.4]
  assign _T_371 = _T_158 ? 3'h3 : 3'h0; // @[Lookup.scala 11:37:@4303.4]
  assign _T_372 = _T_154 ? 3'h3 : _T_371; // @[Lookup.scala 11:37:@4304.4]
  assign _T_373 = _T_150 ? 3'h3 : _T_372; // @[Lookup.scala 11:37:@4305.4]
  assign _T_374 = _T_146 ? 3'h3 : _T_373; // @[Lookup.scala 11:37:@4306.4]
  assign _T_375 = _T_142 ? 3'h3 : _T_374; // @[Lookup.scala 11:37:@4307.4]
  assign _T_376 = _T_138 ? 3'h3 : _T_375; // @[Lookup.scala 11:37:@4308.4]
  assign _T_377 = _T_134 ? 3'h1 : _T_376; // @[Lookup.scala 11:37:@4309.4]
  assign _T_378 = _T_130 ? 3'h5 : _T_377; // @[Lookup.scala 11:37:@4310.4]
  assign _T_379 = _T_126 ? 3'h0 : _T_378; // @[Lookup.scala 11:37:@4311.4]
  assign _T_380 = _T_122 ? 3'h0 : _T_379; // @[Lookup.scala 11:37:@4312.4]
  assign _T_381 = _T_118 ? 3'h0 : _T_380; // @[Lookup.scala 11:37:@4313.4]
  assign _T_382 = _T_114 ? 3'h0 : _T_381; // @[Lookup.scala 11:37:@4314.4]
  assign _T_383 = _T_110 ? 3'h0 : _T_382; // @[Lookup.scala 11:37:@4315.4]
  assign _T_384 = _T_106 ? 3'h0 : _T_383; // @[Lookup.scala 11:37:@4316.4]
  assign _T_385 = _T_102 ? 3'h0 : _T_384; // @[Lookup.scala 11:37:@4317.4]
  assign _T_386 = _T_98 ? 3'h0 : _T_385; // @[Lookup.scala 11:37:@4318.4]
  assign _T_387 = _T_94 ? 3'h0 : _T_386; // @[Lookup.scala 11:37:@4319.4]
  assign _T_388 = _T_90 ? 3'h0 : _T_387; // @[Lookup.scala 11:37:@4320.4]
  assign _T_389 = _T_86 ? 3'h1 : _T_388; // @[Lookup.scala 11:37:@4321.4]
  assign _T_390 = _T_82 ? 3'h1 : _T_389; // @[Lookup.scala 11:37:@4322.4]
  assign _T_391 = _T_78 ? 3'h1 : _T_390; // @[Lookup.scala 11:37:@4323.4]
  assign _T_392 = _T_74 ? 3'h1 : _T_391; // @[Lookup.scala 11:37:@4324.4]
  assign _T_393 = _T_70 ? 3'h1 : _T_392; // @[Lookup.scala 11:37:@4325.4]
  assign _T_394 = _T_66 ? 3'h1 : _T_393; // @[Lookup.scala 11:37:@4326.4]
  assign _T_395 = _T_62 ? 3'h1 : _T_394; // @[Lookup.scala 11:37:@4327.4]
  assign _T_396 = _T_58 ? 3'h1 : _T_395; // @[Lookup.scala 11:37:@4328.4]
  assign _T_397 = _T_54 ? 3'h1 : _T_396; // @[Lookup.scala 11:37:@4329.4]
  assign _T_398 = _T_50 ? 3'h4 : _T_397; // @[Lookup.scala 11:37:@4330.4]
  assign _T_399 = _T_46 ? 3'h4 : _T_398; // @[Lookup.scala 11:37:@4331.4]
  assign _T_400 = _T_42 ? 3'h2 : _T_399; // @[Lookup.scala 11:37:@4332.4]
  assign _T_401 = _T_38 ? 3'h2 : _T_400; // @[Lookup.scala 11:37:@4333.4]
  assign _T_402 = _T_34 ? 3'h2 : _T_401; // @[Lookup.scala 11:37:@4334.4]
  assign _T_403 = _T_30 ? 3'h1 : _T_402; // @[Lookup.scala 11:37:@4335.4]
  assign _T_404 = _T_26 ? 3'h1 : _T_403; // @[Lookup.scala 11:37:@4336.4]
  assign _T_405 = _T_22 ? 3'h1 : _T_404; // @[Lookup.scala 11:37:@4337.4]
  assign _T_406 = _T_18 ? 3'h1 : _T_405; // @[Lookup.scala 11:37:@4338.4]
  assign _T_415 = _T_178 ? 1'h1 : _T_182; // @[Lookup.scala 11:37:@4348.4]
  assign _T_416 = _T_174 ? 1'h1 : _T_415; // @[Lookup.scala 11:37:@4349.4]
  assign _T_417 = _T_170 ? 1'h1 : _T_416; // @[Lookup.scala 11:37:@4350.4]
  assign _T_418 = _T_166 ? 1'h1 : _T_417; // @[Lookup.scala 11:37:@4351.4]
  assign _T_419 = _T_162 ? 1'h1 : _T_418; // @[Lookup.scala 11:37:@4352.4]
  assign _T_420 = _T_158 ? 1'h1 : _T_419; // @[Lookup.scala 11:37:@4353.4]
  assign _T_421 = _T_154 ? 1'h1 : _T_420; // @[Lookup.scala 11:37:@4354.4]
  assign _T_422 = _T_150 ? 1'h1 : _T_421; // @[Lookup.scala 11:37:@4355.4]
  assign _T_423 = _T_146 ? 1'h1 : _T_422; // @[Lookup.scala 11:37:@4356.4]
  assign _T_424 = _T_142 ? 1'h1 : _T_423; // @[Lookup.scala 11:37:@4357.4]
  assign _T_425 = _T_138 ? 1'h1 : _T_424; // @[Lookup.scala 11:37:@4358.4]
  assign _T_426 = _T_134 ? 1'h1 : _T_425; // @[Lookup.scala 11:37:@4359.4]
  assign _T_427 = _T_130 ? 1'h0 : _T_426; // @[Lookup.scala 11:37:@4360.4]
  assign _T_428 = _T_126 ? 1'h1 : _T_427; // @[Lookup.scala 11:37:@4361.4]
  assign _T_429 = _T_122 ? 1'h1 : _T_428; // @[Lookup.scala 11:37:@4362.4]
  assign _T_430 = _T_118 ? 1'h1 : _T_429; // @[Lookup.scala 11:37:@4363.4]
  assign _T_431 = _T_114 ? 1'h1 : _T_430; // @[Lookup.scala 11:37:@4364.4]
  assign _T_432 = _T_110 ? 1'h1 : _T_431; // @[Lookup.scala 11:37:@4365.4]
  assign _T_433 = _T_106 ? 1'h1 : _T_432; // @[Lookup.scala 11:37:@4366.4]
  assign _T_434 = _T_102 ? 1'h1 : _T_433; // @[Lookup.scala 11:37:@4367.4]
  assign _T_435 = _T_98 ? 1'h1 : _T_434; // @[Lookup.scala 11:37:@4368.4]
  assign _T_436 = _T_94 ? 1'h1 : _T_435; // @[Lookup.scala 11:37:@4369.4]
  assign _T_437 = _T_90 ? 1'h1 : _T_436; // @[Lookup.scala 11:37:@4370.4]
  assign _T_438 = _T_86 ? 1'h1 : _T_437; // @[Lookup.scala 11:37:@4371.4]
  assign _T_439 = _T_82 ? 1'h1 : _T_438; // @[Lookup.scala 11:37:@4372.4]
  assign _T_440 = _T_78 ? 1'h1 : _T_439; // @[Lookup.scala 11:37:@4373.4]
  assign _T_441 = _T_74 ? 1'h1 : _T_440; // @[Lookup.scala 11:37:@4374.4]
  assign _T_442 = _T_70 ? 1'h1 : _T_441; // @[Lookup.scala 11:37:@4375.4]
  assign _T_443 = _T_66 ? 1'h1 : _T_442; // @[Lookup.scala 11:37:@4376.4]
  assign _T_444 = _T_62 ? 1'h1 : _T_443; // @[Lookup.scala 11:37:@4377.4]
  assign _T_445 = _T_58 ? 1'h1 : _T_444; // @[Lookup.scala 11:37:@4378.4]
  assign _T_446 = _T_54 ? 1'h1 : _T_445; // @[Lookup.scala 11:37:@4379.4]
  assign _T_447 = _T_50 ? 1'h0 : _T_446; // @[Lookup.scala 11:37:@4380.4]
  assign _T_448 = _T_46 ? 1'h0 : _T_447; // @[Lookup.scala 11:37:@4381.4]
  assign _T_449 = _T_42 ? 1'h1 : _T_448; // @[Lookup.scala 11:37:@4382.4]
  assign _T_450 = _T_38 ? 1'h1 : _T_449; // @[Lookup.scala 11:37:@4383.4]
  assign _T_451 = _T_34 ? 1'h1 : _T_450; // @[Lookup.scala 11:37:@4384.4]
  assign _T_452 = _T_30 ? 1'h1 : _T_451; // @[Lookup.scala 11:37:@4385.4]
  assign _T_453 = _T_26 ? 1'h1 : _T_452; // @[Lookup.scala 11:37:@4386.4]
  assign _T_454 = _T_22 ? 1'h1 : _T_453; // @[Lookup.scala 11:37:@4387.4]
  assign _T_455 = _T_18 ? 1'h1 : _T_454; // @[Lookup.scala 11:37:@4388.4]
  assign _T_475 = _T_134 ? 1'h0 : _T_425; // @[Lookup.scala 11:37:@4409.4]
  assign _T_476 = _T_130 ? 1'h0 : _T_475; // @[Lookup.scala 11:37:@4410.4]
  assign _T_477 = _T_126 ? 1'h1 : _T_476; // @[Lookup.scala 11:37:@4411.4]
  assign _T_478 = _T_122 ? 1'h1 : _T_477; // @[Lookup.scala 11:37:@4412.4]
  assign _T_479 = _T_118 ? 1'h1 : _T_478; // @[Lookup.scala 11:37:@4413.4]
  assign _T_480 = _T_114 ? 1'h1 : _T_479; // @[Lookup.scala 11:37:@4414.4]
  assign _T_481 = _T_110 ? 1'h1 : _T_480; // @[Lookup.scala 11:37:@4415.4]
  assign _T_482 = _T_106 ? 1'h1 : _T_481; // @[Lookup.scala 11:37:@4416.4]
  assign _T_483 = _T_102 ? 1'h1 : _T_482; // @[Lookup.scala 11:37:@4417.4]
  assign _T_484 = _T_98 ? 1'h1 : _T_483; // @[Lookup.scala 11:37:@4418.4]
  assign _T_485 = _T_94 ? 1'h1 : _T_484; // @[Lookup.scala 11:37:@4419.4]
  assign _T_486 = _T_90 ? 1'h1 : _T_485; // @[Lookup.scala 11:37:@4420.4]
  assign _T_487 = _T_86 ? 1'h0 : _T_486; // @[Lookup.scala 11:37:@4421.4]
  assign _T_488 = _T_82 ? 1'h0 : _T_487; // @[Lookup.scala 11:37:@4422.4]
  assign _T_489 = _T_78 ? 1'h0 : _T_488; // @[Lookup.scala 11:37:@4423.4]
  assign _T_490 = _T_74 ? 1'h0 : _T_489; // @[Lookup.scala 11:37:@4424.4]
  assign _T_491 = _T_70 ? 1'h0 : _T_490; // @[Lookup.scala 11:37:@4425.4]
  assign _T_492 = _T_66 ? 1'h0 : _T_491; // @[Lookup.scala 11:37:@4426.4]
  assign _T_493 = _T_62 ? 1'h0 : _T_492; // @[Lookup.scala 11:37:@4427.4]
  assign _T_494 = _T_58 ? 1'h0 : _T_493; // @[Lookup.scala 11:37:@4428.4]
  assign _T_495 = _T_54 ? 1'h0 : _T_494; // @[Lookup.scala 11:37:@4429.4]
  assign _T_496 = _T_50 ? 1'h0 : _T_495; // @[Lookup.scala 11:37:@4430.4]
  assign _T_497 = _T_46 ? 1'h0 : _T_496; // @[Lookup.scala 11:37:@4431.4]
  assign _T_498 = _T_42 ? 1'h1 : _T_497; // @[Lookup.scala 11:37:@4432.4]
  assign _T_499 = _T_38 ? 1'h1 : _T_498; // @[Lookup.scala 11:37:@4433.4]
  assign _T_500 = _T_34 ? 1'h1 : _T_499; // @[Lookup.scala 11:37:@4434.4]
  assign _T_501 = _T_30 ? 1'h0 : _T_500; // @[Lookup.scala 11:37:@4435.4]
  assign _T_502 = _T_26 ? 1'h0 : _T_501; // @[Lookup.scala 11:37:@4436.4]
  assign _T_503 = _T_22 ? 1'h0 : _T_502; // @[Lookup.scala 11:37:@4437.4]
  assign _T_504 = _T_18 ? 1'h0 : _T_503; // @[Lookup.scala 11:37:@4438.4]
  assign _T_512 = _T_182 ? 4'ha : 4'h0; // @[Lookup.scala 11:37:@4447.4]
  assign _T_513 = _T_178 ? 4'ha : _T_512; // @[Lookup.scala 11:37:@4448.4]
  assign _T_514 = _T_174 ? 4'ha : _T_513; // @[Lookup.scala 11:37:@4449.4]
  assign _T_515 = _T_170 ? 4'ha : _T_514; // @[Lookup.scala 11:37:@4450.4]
  assign _T_516 = _T_166 ? 4'ha : _T_515; // @[Lookup.scala 11:37:@4451.4]
  assign _T_517 = _T_162 ? 4'ha : _T_516; // @[Lookup.scala 11:37:@4452.4]
  assign _T_518 = _T_158 ? 4'h0 : _T_517; // @[Lookup.scala 11:37:@4453.4]
  assign _T_519 = _T_154 ? 4'h0 : _T_518; // @[Lookup.scala 11:37:@4454.4]
  assign _T_520 = _T_150 ? 4'h0 : _T_519; // @[Lookup.scala 11:37:@4455.4]
  assign _T_521 = _T_146 ? 4'h0 : _T_520; // @[Lookup.scala 11:37:@4456.4]
  assign _T_522 = _T_142 ? 4'h0 : _T_521; // @[Lookup.scala 11:37:@4457.4]
  assign _T_523 = _T_138 ? 4'h0 : _T_522; // @[Lookup.scala 11:37:@4458.4]
  assign _T_524 = _T_134 ? 4'h0 : _T_523; // @[Lookup.scala 11:37:@4459.4]
  assign _T_525 = _T_130 ? 4'h0 : _T_524; // @[Lookup.scala 11:37:@4460.4]
  assign _T_526 = _T_126 ? 4'h3 : _T_525; // @[Lookup.scala 11:37:@4461.4]
  assign _T_527 = _T_122 ? 4'h4 : _T_526; // @[Lookup.scala 11:37:@4462.4]
  assign _T_528 = _T_118 ? 4'h7 : _T_527; // @[Lookup.scala 11:37:@4463.4]
  assign _T_529 = _T_114 ? 4'h6 : _T_528; // @[Lookup.scala 11:37:@4464.4]
  assign _T_530 = _T_110 ? 4'h5 : _T_529; // @[Lookup.scala 11:37:@4465.4]
  assign _T_531 = _T_106 ? 4'h9 : _T_530; // @[Lookup.scala 11:37:@4466.4]
  assign _T_532 = _T_102 ? 4'h8 : _T_531; // @[Lookup.scala 11:37:@4467.4]
  assign _T_533 = _T_98 ? 4'h1 : _T_532; // @[Lookup.scala 11:37:@4468.4]
  assign _T_534 = _T_94 ? 4'h0 : _T_533; // @[Lookup.scala 11:37:@4469.4]
  assign _T_535 = _T_90 ? 4'h2 : _T_534; // @[Lookup.scala 11:37:@4470.4]
  assign _T_536 = _T_86 ? 4'h3 : _T_535; // @[Lookup.scala 11:37:@4471.4]
  assign _T_537 = _T_82 ? 4'h4 : _T_536; // @[Lookup.scala 11:37:@4472.4]
  assign _T_538 = _T_78 ? 4'h2 : _T_537; // @[Lookup.scala 11:37:@4473.4]
  assign _T_539 = _T_74 ? 4'h9 : _T_538; // @[Lookup.scala 11:37:@4474.4]
  assign _T_540 = _T_70 ? 4'h8 : _T_539; // @[Lookup.scala 11:37:@4475.4]
  assign _T_541 = _T_66 ? 4'h7 : _T_540; // @[Lookup.scala 11:37:@4476.4]
  assign _T_542 = _T_62 ? 4'h6 : _T_541; // @[Lookup.scala 11:37:@4477.4]
  assign _T_543 = _T_58 ? 4'h5 : _T_542; // @[Lookup.scala 11:37:@4478.4]
  assign _T_544 = _T_54 ? 4'h0 : _T_543; // @[Lookup.scala 11:37:@4479.4]
  assign _T_545 = _T_50 ? 4'hb : _T_544; // @[Lookup.scala 11:37:@4480.4]
  assign _T_546 = _T_46 ? 4'h0 : _T_545; // @[Lookup.scala 11:37:@4481.4]
  assign _T_547 = _T_42 ? 4'h0 : _T_546; // @[Lookup.scala 11:37:@4482.4]
  assign _T_548 = _T_38 ? 4'h0 : _T_547; // @[Lookup.scala 11:37:@4483.4]
  assign _T_549 = _T_34 ? 4'h0 : _T_548; // @[Lookup.scala 11:37:@4484.4]
  assign _T_550 = _T_30 ? 4'h0 : _T_549; // @[Lookup.scala 11:37:@4485.4]
  assign _T_551 = _T_26 ? 4'h0 : _T_550; // @[Lookup.scala 11:37:@4486.4]
  assign _T_552 = _T_22 ? 4'h0 : _T_551; // @[Lookup.scala 11:37:@4487.4]
  assign _T_553 = _T_18 ? 4'h0 : _T_552; // @[Lookup.scala 11:37:@4488.4]
  assign _T_561 = _T_182 ? 2'h3 : 2'h0; // @[Lookup.scala 11:37:@4497.4]
  assign _T_562 = _T_178 ? 2'h3 : _T_561; // @[Lookup.scala 11:37:@4498.4]
  assign _T_563 = _T_174 ? 2'h3 : _T_562; // @[Lookup.scala 11:37:@4499.4]
  assign _T_564 = _T_170 ? 2'h3 : _T_563; // @[Lookup.scala 11:37:@4500.4]
  assign _T_565 = _T_166 ? 2'h3 : _T_564; // @[Lookup.scala 11:37:@4501.4]
  assign _T_566 = _T_162 ? 2'h3 : _T_565; // @[Lookup.scala 11:37:@4502.4]
  assign _T_567 = _T_158 ? 2'h0 : _T_566; // @[Lookup.scala 11:37:@4503.4]
  assign _T_568 = _T_154 ? 2'h0 : _T_567; // @[Lookup.scala 11:37:@4504.4]
  assign _T_569 = _T_150 ? 2'h0 : _T_568; // @[Lookup.scala 11:37:@4505.4]
  assign _T_570 = _T_146 ? 2'h0 : _T_569; // @[Lookup.scala 11:37:@4506.4]
  assign _T_571 = _T_142 ? 2'h0 : _T_570; // @[Lookup.scala 11:37:@4507.4]
  assign _T_572 = _T_138 ? 2'h0 : _T_571; // @[Lookup.scala 11:37:@4508.4]
  assign _T_573 = _T_134 ? 2'h2 : _T_572; // @[Lookup.scala 11:37:@4509.4]
  assign _T_574 = _T_130 ? 2'h2 : _T_573; // @[Lookup.scala 11:37:@4510.4]
  assign _T_575 = _T_126 ? 2'h0 : _T_574; // @[Lookup.scala 11:37:@4511.4]
  assign _T_576 = _T_122 ? 2'h0 : _T_575; // @[Lookup.scala 11:37:@4512.4]
  assign _T_577 = _T_118 ? 2'h0 : _T_576; // @[Lookup.scala 11:37:@4513.4]
  assign _T_578 = _T_114 ? 2'h0 : _T_577; // @[Lookup.scala 11:37:@4514.4]
  assign _T_579 = _T_110 ? 2'h0 : _T_578; // @[Lookup.scala 11:37:@4515.4]
  assign _T_580 = _T_106 ? 2'h0 : _T_579; // @[Lookup.scala 11:37:@4516.4]
  assign _T_581 = _T_102 ? 2'h0 : _T_580; // @[Lookup.scala 11:37:@4517.4]
  assign _T_582 = _T_98 ? 2'h0 : _T_581; // @[Lookup.scala 11:37:@4518.4]
  assign _T_583 = _T_94 ? 2'h0 : _T_582; // @[Lookup.scala 11:37:@4519.4]
  assign _T_584 = _T_90 ? 2'h0 : _T_583; // @[Lookup.scala 11:37:@4520.4]
  assign _T_585 = _T_86 ? 2'h0 : _T_584; // @[Lookup.scala 11:37:@4521.4]
  assign _T_586 = _T_82 ? 2'h0 : _T_585; // @[Lookup.scala 11:37:@4522.4]
  assign _T_587 = _T_78 ? 2'h0 : _T_586; // @[Lookup.scala 11:37:@4523.4]
  assign _T_588 = _T_74 ? 2'h0 : _T_587; // @[Lookup.scala 11:37:@4524.4]
  assign _T_589 = _T_70 ? 2'h0 : _T_588; // @[Lookup.scala 11:37:@4525.4]
  assign _T_590 = _T_66 ? 2'h0 : _T_589; // @[Lookup.scala 11:37:@4526.4]
  assign _T_591 = _T_62 ? 2'h0 : _T_590; // @[Lookup.scala 11:37:@4527.4]
  assign _T_592 = _T_58 ? 2'h0 : _T_591; // @[Lookup.scala 11:37:@4528.4]
  assign _T_593 = _T_54 ? 2'h0 : _T_592; // @[Lookup.scala 11:37:@4529.4]
  assign _T_594 = _T_50 ? 2'h0 : _T_593; // @[Lookup.scala 11:37:@4530.4]
  assign _T_595 = _T_46 ? 2'h0 : _T_594; // @[Lookup.scala 11:37:@4531.4]
  assign _T_596 = _T_42 ? 2'h0 : _T_595; // @[Lookup.scala 11:37:@4532.4]
  assign _T_597 = _T_38 ? 2'h0 : _T_596; // @[Lookup.scala 11:37:@4533.4]
  assign _T_598 = _T_34 ? 2'h0 : _T_597; // @[Lookup.scala 11:37:@4534.4]
  assign _T_599 = _T_30 ? 2'h1 : _T_598; // @[Lookup.scala 11:37:@4535.4]
  assign _T_600 = _T_26 ? 2'h1 : _T_599; // @[Lookup.scala 11:37:@4536.4]
  assign _T_601 = _T_22 ? 2'h1 : _T_600; // @[Lookup.scala 11:37:@4537.4]
  assign _T_602 = _T_18 ? 2'h1 : _T_601; // @[Lookup.scala 11:37:@4538.4]
  assign _T_616 = _T_158 ? 1'h0 : _T_419; // @[Lookup.scala 11:37:@4553.4]
  assign _T_617 = _T_154 ? 1'h0 : _T_616; // @[Lookup.scala 11:37:@4554.4]
  assign _T_618 = _T_150 ? 1'h0 : _T_617; // @[Lookup.scala 11:37:@4555.4]
  assign _T_619 = _T_146 ? 1'h0 : _T_618; // @[Lookup.scala 11:37:@4556.4]
  assign _T_620 = _T_142 ? 1'h0 : _T_619; // @[Lookup.scala 11:37:@4557.4]
  assign _T_621 = _T_138 ? 1'h0 : _T_620; // @[Lookup.scala 11:37:@4558.4]
  assign _T_622 = _T_134 ? 1'h1 : _T_621; // @[Lookup.scala 11:37:@4559.4]
  assign _T_623 = _T_130 ? 1'h1 : _T_622; // @[Lookup.scala 11:37:@4560.4]
  assign _T_624 = _T_126 ? 1'h1 : _T_623; // @[Lookup.scala 11:37:@4561.4]
  assign _T_625 = _T_122 ? 1'h1 : _T_624; // @[Lookup.scala 11:37:@4562.4]
  assign _T_626 = _T_118 ? 1'h1 : _T_625; // @[Lookup.scala 11:37:@4563.4]
  assign _T_627 = _T_114 ? 1'h1 : _T_626; // @[Lookup.scala 11:37:@4564.4]
  assign _T_628 = _T_110 ? 1'h1 : _T_627; // @[Lookup.scala 11:37:@4565.4]
  assign _T_629 = _T_106 ? 1'h1 : _T_628; // @[Lookup.scala 11:37:@4566.4]
  assign _T_630 = _T_102 ? 1'h1 : _T_629; // @[Lookup.scala 11:37:@4567.4]
  assign _T_631 = _T_98 ? 1'h1 : _T_630; // @[Lookup.scala 11:37:@4568.4]
  assign _T_632 = _T_94 ? 1'h1 : _T_631; // @[Lookup.scala 11:37:@4569.4]
  assign _T_633 = _T_90 ? 1'h1 : _T_632; // @[Lookup.scala 11:37:@4570.4]
  assign _T_634 = _T_86 ? 1'h1 : _T_633; // @[Lookup.scala 11:37:@4571.4]
  assign _T_635 = _T_82 ? 1'h1 : _T_634; // @[Lookup.scala 11:37:@4572.4]
  assign _T_636 = _T_78 ? 1'h1 : _T_635; // @[Lookup.scala 11:37:@4573.4]
  assign _T_637 = _T_74 ? 1'h1 : _T_636; // @[Lookup.scala 11:37:@4574.4]
  assign _T_638 = _T_70 ? 1'h1 : _T_637; // @[Lookup.scala 11:37:@4575.4]
  assign _T_639 = _T_66 ? 1'h1 : _T_638; // @[Lookup.scala 11:37:@4576.4]
  assign _T_640 = _T_62 ? 1'h1 : _T_639; // @[Lookup.scala 11:37:@4577.4]
  assign _T_641 = _T_58 ? 1'h1 : _T_640; // @[Lookup.scala 11:37:@4578.4]
  assign _T_642 = _T_54 ? 1'h1 : _T_641; // @[Lookup.scala 11:37:@4579.4]
  assign _T_643 = _T_50 ? 1'h1 : _T_642; // @[Lookup.scala 11:37:@4580.4]
  assign _T_644 = _T_46 ? 1'h1 : _T_643; // @[Lookup.scala 11:37:@4581.4]
  assign _T_645 = _T_42 ? 1'h0 : _T_644; // @[Lookup.scala 11:37:@4582.4]
  assign _T_646 = _T_38 ? 1'h0 : _T_645; // @[Lookup.scala 11:37:@4583.4]
  assign _T_647 = _T_34 ? 1'h0 : _T_646; // @[Lookup.scala 11:37:@4584.4]
  assign _T_648 = _T_30 ? 1'h1 : _T_647; // @[Lookup.scala 11:37:@4585.4]
  assign _T_649 = _T_26 ? 1'h1 : _T_648; // @[Lookup.scala 11:37:@4586.4]
  assign _T_650 = _T_22 ? 1'h1 : _T_649; // @[Lookup.scala 11:37:@4587.4]
  assign _T_651 = _T_18 ? 1'h1 : _T_650; // @[Lookup.scala 11:37:@4588.4]
  assign _T_653 = _T_206 ? 1'h0 : _T_210; // @[Lookup.scala 11:37:@4591.4]
  assign _T_654 = _T_202 ? 1'h0 : _T_653; // @[Lookup.scala 11:37:@4592.4]
  assign _T_655 = _T_198 ? 1'h0 : _T_654; // @[Lookup.scala 11:37:@4593.4]
  assign _T_656 = _T_194 ? 1'h0 : _T_655; // @[Lookup.scala 11:37:@4594.4]
  assign _T_657 = _T_190 ? 1'h0 : _T_656; // @[Lookup.scala 11:37:@4595.4]
  assign _T_658 = _T_186 ? 1'h0 : _T_657; // @[Lookup.scala 11:37:@4596.4]
  assign _T_659 = _T_182 ? 1'h0 : _T_658; // @[Lookup.scala 11:37:@4597.4]
  assign _T_660 = _T_178 ? 1'h0 : _T_659; // @[Lookup.scala 11:37:@4598.4]
  assign _T_661 = _T_174 ? 1'h0 : _T_660; // @[Lookup.scala 11:37:@4599.4]
  assign _T_662 = _T_170 ? 1'h0 : _T_661; // @[Lookup.scala 11:37:@4600.4]
  assign _T_663 = _T_166 ? 1'h0 : _T_662; // @[Lookup.scala 11:37:@4601.4]
  assign _T_664 = _T_162 ? 1'h0 : _T_663; // @[Lookup.scala 11:37:@4602.4]
  assign _T_665 = _T_158 ? 1'h0 : _T_664; // @[Lookup.scala 11:37:@4603.4]
  assign _T_666 = _T_154 ? 1'h0 : _T_665; // @[Lookup.scala 11:37:@4604.4]
  assign _T_667 = _T_150 ? 1'h0 : _T_666; // @[Lookup.scala 11:37:@4605.4]
  assign _T_668 = _T_146 ? 1'h0 : _T_667; // @[Lookup.scala 11:37:@4606.4]
  assign _T_669 = _T_142 ? 1'h0 : _T_668; // @[Lookup.scala 11:37:@4607.4]
  assign _T_670 = _T_138 ? 1'h0 : _T_669; // @[Lookup.scala 11:37:@4608.4]
  assign _T_671 = _T_134 ? 1'h0 : _T_670; // @[Lookup.scala 11:37:@4609.4]
  assign _T_672 = _T_130 ? 1'h0 : _T_671; // @[Lookup.scala 11:37:@4610.4]
  assign _T_673 = _T_126 ? 1'h0 : _T_672; // @[Lookup.scala 11:37:@4611.4]
  assign _T_674 = _T_122 ? 1'h0 : _T_673; // @[Lookup.scala 11:37:@4612.4]
  assign _T_675 = _T_118 ? 1'h0 : _T_674; // @[Lookup.scala 11:37:@4613.4]
  assign _T_676 = _T_114 ? 1'h0 : _T_675; // @[Lookup.scala 11:37:@4614.4]
  assign _T_677 = _T_110 ? 1'h0 : _T_676; // @[Lookup.scala 11:37:@4615.4]
  assign _T_678 = _T_106 ? 1'h0 : _T_677; // @[Lookup.scala 11:37:@4616.4]
  assign _T_679 = _T_102 ? 1'h0 : _T_678; // @[Lookup.scala 11:37:@4617.4]
  assign _T_680 = _T_98 ? 1'h0 : _T_679; // @[Lookup.scala 11:37:@4618.4]
  assign _T_681 = _T_94 ? 1'h0 : _T_680; // @[Lookup.scala 11:37:@4619.4]
  assign _T_682 = _T_90 ? 1'h0 : _T_681; // @[Lookup.scala 11:37:@4620.4]
  assign _T_683 = _T_86 ? 1'h0 : _T_682; // @[Lookup.scala 11:37:@4621.4]
  assign _T_684 = _T_82 ? 1'h0 : _T_683; // @[Lookup.scala 11:37:@4622.4]
  assign _T_685 = _T_78 ? 1'h0 : _T_684; // @[Lookup.scala 11:37:@4623.4]
  assign _T_686 = _T_74 ? 1'h0 : _T_685; // @[Lookup.scala 11:37:@4624.4]
  assign _T_687 = _T_70 ? 1'h0 : _T_686; // @[Lookup.scala 11:37:@4625.4]
  assign _T_688 = _T_66 ? 1'h0 : _T_687; // @[Lookup.scala 11:37:@4626.4]
  assign _T_689 = _T_62 ? 1'h0 : _T_688; // @[Lookup.scala 11:37:@4627.4]
  assign _T_690 = _T_58 ? 1'h0 : _T_689; // @[Lookup.scala 11:37:@4628.4]
  assign _T_691 = _T_54 ? 1'h0 : _T_690; // @[Lookup.scala 11:37:@4629.4]
  assign _T_692 = _T_50 ? 1'h0 : _T_691; // @[Lookup.scala 11:37:@4630.4]
  assign _T_693 = _T_46 ? 1'h0 : _T_692; // @[Lookup.scala 11:37:@4631.4]
  assign _T_694 = _T_42 ? 1'h1 : _T_693; // @[Lookup.scala 11:37:@4632.4]
  assign _T_695 = _T_38 ? 1'h1 : _T_694; // @[Lookup.scala 11:37:@4633.4]
  assign _T_696 = _T_34 ? 1'h1 : _T_695; // @[Lookup.scala 11:37:@4634.4]
  assign _T_697 = _T_30 ? 1'h1 : _T_696; // @[Lookup.scala 11:37:@4635.4]
  assign _T_698 = _T_26 ? 1'h1 : _T_697; // @[Lookup.scala 11:37:@4636.4]
  assign _T_699 = _T_22 ? 1'h1 : _T_698; // @[Lookup.scala 11:37:@4637.4]
  assign _T_700 = _T_18 ? 1'h1 : _T_699; // @[Lookup.scala 11:37:@4638.4]
  assign _T_744 = _T_38 ? 1'h1 : _T_42; // @[Lookup.scala 11:37:@4683.4]
  assign _T_745 = _T_34 ? 1'h1 : _T_744; // @[Lookup.scala 11:37:@4684.4]
  assign _T_746 = _T_30 ? 1'h0 : _T_745; // @[Lookup.scala 11:37:@4685.4]
  assign _T_747 = _T_26 ? 1'h0 : _T_746; // @[Lookup.scala 11:37:@4686.4]
  assign _T_748 = _T_22 ? 1'h0 : _T_747; // @[Lookup.scala 11:37:@4687.4]
  assign _T_749 = _T_18 ? 1'h0 : _T_748; // @[Lookup.scala 11:37:@4688.4]
  assign _T_792 = _T_42 ? 3'h2 : 3'h0; // @[Lookup.scala 11:37:@4732.4]
  assign _T_793 = _T_38 ? 3'h1 : _T_792; // @[Lookup.scala 11:37:@4733.4]
  assign _T_794 = _T_34 ? 3'h3 : _T_793; // @[Lookup.scala 11:37:@4734.4]
  assign _T_795 = _T_30 ? 3'h6 : _T_794; // @[Lookup.scala 11:37:@4735.4]
  assign _T_796 = _T_26 ? 3'h2 : _T_795; // @[Lookup.scala 11:37:@4736.4]
  assign _T_797 = _T_22 ? 3'h5 : _T_796; // @[Lookup.scala 11:37:@4737.4]
  assign _T_798 = _T_18 ? 3'h1 : _T_797; // @[Lookup.scala 11:37:@4738.4]
  assign _T_802 = _T_198 ? 3'h4 : 3'h0; // @[Lookup.scala 11:37:@4743.4]
  assign _T_803 = _T_194 ? 3'h4 : _T_802; // @[Lookup.scala 11:37:@4744.4]
  assign _T_804 = _T_190 ? 3'h4 : _T_803; // @[Lookup.scala 11:37:@4745.4]
  assign _T_805 = _T_186 ? 3'h4 : _T_804; // @[Lookup.scala 11:37:@4746.4]
  assign _T_806 = _T_182 ? 3'h3 : _T_805; // @[Lookup.scala 11:37:@4747.4]
  assign _T_807 = _T_178 ? 3'h3 : _T_806; // @[Lookup.scala 11:37:@4748.4]
  assign _T_808 = _T_174 ? 3'h2 : _T_807; // @[Lookup.scala 11:37:@4749.4]
  assign _T_809 = _T_170 ? 3'h1 : _T_808; // @[Lookup.scala 11:37:@4750.4]
  assign _T_810 = _T_166 ? 3'h2 : _T_809; // @[Lookup.scala 11:37:@4751.4]
  assign _T_811 = _T_162 ? 3'h1 : _T_810; // @[Lookup.scala 11:37:@4752.4]
  assign _T_812 = _T_158 ? 3'h0 : _T_811; // @[Lookup.scala 11:37:@4753.4]
  assign _T_813 = _T_154 ? 3'h0 : _T_812; // @[Lookup.scala 11:37:@4754.4]
  assign _T_814 = _T_150 ? 3'h0 : _T_813; // @[Lookup.scala 11:37:@4755.4]
  assign _T_815 = _T_146 ? 3'h0 : _T_814; // @[Lookup.scala 11:37:@4756.4]
  assign _T_816 = _T_142 ? 3'h0 : _T_815; // @[Lookup.scala 11:37:@4757.4]
  assign _T_817 = _T_138 ? 3'h0 : _T_816; // @[Lookup.scala 11:37:@4758.4]
  assign _T_818 = _T_134 ? 3'h0 : _T_817; // @[Lookup.scala 11:37:@4759.4]
  assign _T_819 = _T_130 ? 3'h0 : _T_818; // @[Lookup.scala 11:37:@4760.4]
  assign _T_820 = _T_126 ? 3'h0 : _T_819; // @[Lookup.scala 11:37:@4761.4]
  assign _T_821 = _T_122 ? 3'h0 : _T_820; // @[Lookup.scala 11:37:@4762.4]
  assign _T_822 = _T_118 ? 3'h0 : _T_821; // @[Lookup.scala 11:37:@4763.4]
  assign _T_823 = _T_114 ? 3'h0 : _T_822; // @[Lookup.scala 11:37:@4764.4]
  assign _T_824 = _T_110 ? 3'h0 : _T_823; // @[Lookup.scala 11:37:@4765.4]
  assign _T_825 = _T_106 ? 3'h0 : _T_824; // @[Lookup.scala 11:37:@4766.4]
  assign _T_826 = _T_102 ? 3'h0 : _T_825; // @[Lookup.scala 11:37:@4767.4]
  assign _T_827 = _T_98 ? 3'h0 : _T_826; // @[Lookup.scala 11:37:@4768.4]
  assign _T_828 = _T_94 ? 3'h0 : _T_827; // @[Lookup.scala 11:37:@4769.4]
  assign _T_829 = _T_90 ? 3'h0 : _T_828; // @[Lookup.scala 11:37:@4770.4]
  assign _T_830 = _T_86 ? 3'h0 : _T_829; // @[Lookup.scala 11:37:@4771.4]
  assign _T_831 = _T_82 ? 3'h0 : _T_830; // @[Lookup.scala 11:37:@4772.4]
  assign _T_832 = _T_78 ? 3'h0 : _T_831; // @[Lookup.scala 11:37:@4773.4]
  assign _T_833 = _T_74 ? 3'h0 : _T_832; // @[Lookup.scala 11:37:@4774.4]
  assign _T_834 = _T_70 ? 3'h0 : _T_833; // @[Lookup.scala 11:37:@4775.4]
  assign _T_835 = _T_66 ? 3'h0 : _T_834; // @[Lookup.scala 11:37:@4776.4]
  assign _T_836 = _T_62 ? 3'h0 : _T_835; // @[Lookup.scala 11:37:@4777.4]
  assign _T_837 = _T_58 ? 3'h0 : _T_836; // @[Lookup.scala 11:37:@4778.4]
  assign _T_838 = _T_54 ? 3'h0 : _T_837; // @[Lookup.scala 11:37:@4779.4]
  assign _T_839 = _T_50 ? 3'h0 : _T_838; // @[Lookup.scala 11:37:@4780.4]
  assign _T_840 = _T_46 ? 3'h0 : _T_839; // @[Lookup.scala 11:37:@4781.4]
  assign _T_841 = _T_42 ? 3'h0 : _T_840; // @[Lookup.scala 11:37:@4782.4]
  assign _T_842 = _T_38 ? 3'h0 : _T_841; // @[Lookup.scala 11:37:@4783.4]
  assign _T_843 = _T_34 ? 3'h0 : _T_842; // @[Lookup.scala 11:37:@4784.4]
  assign _T_844 = _T_30 ? 3'h0 : _T_843; // @[Lookup.scala 11:37:@4785.4]
  assign _T_845 = _T_26 ? 3'h0 : _T_844; // @[Lookup.scala 11:37:@4786.4]
  assign _T_846 = _T_22 ? 3'h0 : _T_845; // @[Lookup.scala 11:37:@4787.4]
  assign _T_847 = _T_18 ? 3'h0 : _T_846; // @[Lookup.scala 11:37:@4788.4]
  assign _T_850 = _T_202 ? 1'h0 : _T_206; // @[Lookup.scala 11:37:@4792.4]
  assign _T_851 = _T_198 ? 1'h0 : _T_850; // @[Lookup.scala 11:37:@4793.4]
  assign _T_852 = _T_194 ? 1'h0 : _T_851; // @[Lookup.scala 11:37:@4794.4]
  assign _T_853 = _T_190 ? 1'h0 : _T_852; // @[Lookup.scala 11:37:@4795.4]
  assign _T_854 = _T_186 ? 1'h0 : _T_853; // @[Lookup.scala 11:37:@4796.4]
  assign _T_855 = _T_182 ? 1'h0 : _T_854; // @[Lookup.scala 11:37:@4797.4]
  assign _T_856 = _T_178 ? 1'h0 : _T_855; // @[Lookup.scala 11:37:@4798.4]
  assign _T_857 = _T_174 ? 1'h0 : _T_856; // @[Lookup.scala 11:37:@4799.4]
  assign _T_858 = _T_170 ? 1'h0 : _T_857; // @[Lookup.scala 11:37:@4800.4]
  assign _T_859 = _T_166 ? 1'h0 : _T_858; // @[Lookup.scala 11:37:@4801.4]
  assign _T_860 = _T_162 ? 1'h0 : _T_859; // @[Lookup.scala 11:37:@4802.4]
  assign _T_861 = _T_158 ? 1'h0 : _T_860; // @[Lookup.scala 11:37:@4803.4]
  assign _T_862 = _T_154 ? 1'h0 : _T_861; // @[Lookup.scala 11:37:@4804.4]
  assign _T_863 = _T_150 ? 1'h0 : _T_862; // @[Lookup.scala 11:37:@4805.4]
  assign _T_864 = _T_146 ? 1'h0 : _T_863; // @[Lookup.scala 11:37:@4806.4]
  assign _T_865 = _T_142 ? 1'h0 : _T_864; // @[Lookup.scala 11:37:@4807.4]
  assign _T_866 = _T_138 ? 1'h0 : _T_865; // @[Lookup.scala 11:37:@4808.4]
  assign _T_867 = _T_134 ? 1'h0 : _T_866; // @[Lookup.scala 11:37:@4809.4]
  assign _T_868 = _T_130 ? 1'h0 : _T_867; // @[Lookup.scala 11:37:@4810.4]
  assign _T_869 = _T_126 ? 1'h0 : _T_868; // @[Lookup.scala 11:37:@4811.4]
  assign _T_870 = _T_122 ? 1'h0 : _T_869; // @[Lookup.scala 11:37:@4812.4]
  assign _T_871 = _T_118 ? 1'h0 : _T_870; // @[Lookup.scala 11:37:@4813.4]
  assign _T_872 = _T_114 ? 1'h0 : _T_871; // @[Lookup.scala 11:37:@4814.4]
  assign _T_873 = _T_110 ? 1'h0 : _T_872; // @[Lookup.scala 11:37:@4815.4]
  assign _T_874 = _T_106 ? 1'h0 : _T_873; // @[Lookup.scala 11:37:@4816.4]
  assign _T_875 = _T_102 ? 1'h0 : _T_874; // @[Lookup.scala 11:37:@4817.4]
  assign _T_876 = _T_98 ? 1'h0 : _T_875; // @[Lookup.scala 11:37:@4818.4]
  assign _T_877 = _T_94 ? 1'h0 : _T_876; // @[Lookup.scala 11:37:@4819.4]
  assign _T_878 = _T_90 ? 1'h0 : _T_877; // @[Lookup.scala 11:37:@4820.4]
  assign _T_879 = _T_86 ? 1'h0 : _T_878; // @[Lookup.scala 11:37:@4821.4]
  assign _T_880 = _T_82 ? 1'h0 : _T_879; // @[Lookup.scala 11:37:@4822.4]
  assign _T_881 = _T_78 ? 1'h0 : _T_880; // @[Lookup.scala 11:37:@4823.4]
  assign _T_882 = _T_74 ? 1'h0 : _T_881; // @[Lookup.scala 11:37:@4824.4]
  assign _T_883 = _T_70 ? 1'h0 : _T_882; // @[Lookup.scala 11:37:@4825.4]
  assign _T_884 = _T_66 ? 1'h0 : _T_883; // @[Lookup.scala 11:37:@4826.4]
  assign _T_885 = _T_62 ? 1'h0 : _T_884; // @[Lookup.scala 11:37:@4827.4]
  assign _T_886 = _T_58 ? 1'h0 : _T_885; // @[Lookup.scala 11:37:@4828.4]
  assign _T_887 = _T_54 ? 1'h0 : _T_886; // @[Lookup.scala 11:37:@4829.4]
  assign _T_888 = _T_50 ? 1'h0 : _T_887; // @[Lookup.scala 11:37:@4830.4]
  assign _T_889 = _T_46 ? 1'h0 : _T_888; // @[Lookup.scala 11:37:@4831.4]
  assign _T_890 = _T_42 ? 1'h0 : _T_889; // @[Lookup.scala 11:37:@4832.4]
  assign _T_891 = _T_38 ? 1'h0 : _T_890; // @[Lookup.scala 11:37:@4833.4]
  assign _T_892 = _T_34 ? 1'h0 : _T_891; // @[Lookup.scala 11:37:@4834.4]
  assign _T_893 = _T_30 ? 1'h0 : _T_892; // @[Lookup.scala 11:37:@4835.4]
  assign _T_894 = _T_26 ? 1'h0 : _T_893; // @[Lookup.scala 11:37:@4836.4]
  assign _T_895 = _T_22 ? 1'h0 : _T_894; // @[Lookup.scala 11:37:@4837.4]
  assign _T_896 = _T_18 ? 1'h0 : _T_895; // @[Lookup.scala 11:37:@4838.4]
  assign _T_899 = io_inst[19:15]; // @[InstDecoder.scala 130:31:@4855.4]
  assign _T_901 = io_inst[11:7]; // @[InstDecoder.scala 132:31:@4859.4]
  assign func = io_inst[6:2]; // @[InstDecoder.scala 134:21:@4861.4]
  assign _T_905 = func == 5'h1b; // @[InstDecoder.scala 136:38:@4864.4]
  assign _T_907 = func == 5'h19; // @[InstDecoder.scala 137:39:@4865.4]
  assign _T_908 = _T_905 | _T_907; // @[InstDecoder.scala 141:32:@4866.4]
  assign _T_910 = io_cinfo_wbaddr == 5'h1; // @[InstDecoder.scala 135:37:@4867.4]
  assign _T_912 = io_cinfo_wbaddr == 5'h5; // @[InstDecoder.scala 135:53:@4868.4]
  assign _T_913 = _T_910 | _T_912; // @[InstDecoder.scala 135:45:@4869.4]
  assign _GEN_0 = {{4'd0}, _T_907}; // @[InstDecoder.scala 142:24:@4873.4]
  assign _T_917 = func == _GEN_0; // @[InstDecoder.scala 142:24:@4873.4]
  assign _T_919 = io_cinfo_rs1_addr == 5'h1; // @[InstDecoder.scala 135:37:@4874.4]
  assign _T_921 = io_cinfo_rs1_addr == 5'h5; // @[InstDecoder.scala 135:53:@4875.4]
  assign _T_922 = _T_919 | _T_921; // @[InstDecoder.scala 135:45:@4876.4]
  assign _T_923 = _T_917 & _T_922; // @[InstDecoder.scala 142:41:@4877.4]
  assign _T_930 = _T_913 == 1'h0; // @[InstDecoder.scala 143:6:@4881.4]
  assign _T_931 = io_cinfo_rs1_addr != io_cinfo_wbaddr; // @[InstDecoder.scala 143:50:@4882.4]
  assign _T_932 = _T_930 | _T_931; // @[InstDecoder.scala 143:29:@4883.4]
  assign imm_itype = io_inst[31:20]; // @[InstDecoder.scala 146:27:@4886.4]
  assign _T_934 = io_inst[31:25]; // @[InstDecoder.scala 147:31:@4887.4]
  assign imm_stype = {_T_934,_T_901}; // @[Cat.scala 30:58:@4889.4]
  assign _T_936 = io_inst[31]; // @[InstDecoder.scala 148:31:@4890.4]
  assign _T_937 = io_inst[7]; // @[InstDecoder.scala 148:44:@4891.4]
  assign _T_938 = io_inst[30:25]; // @[InstDecoder.scala 148:56:@4892.4]
  assign _T_939 = io_inst[11:8]; // @[InstDecoder.scala 148:73:@4893.4]
  assign imm_sbtype = {_T_936,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@4896.4]
  assign imm_utype = io_inst[31:12]; // @[InstDecoder.scala 149:27:@4897.4]
  assign _T_943 = io_inst[19:12]; // @[InstDecoder.scala 150:44:@4899.4]
  assign _T_944 = io_inst[20]; // @[InstDecoder.scala 150:60:@4900.4]
  assign _T_945 = io_inst[30:21]; // @[InstDecoder.scala 150:73:@4901.4]
  assign imm_ujtype = {_T_936,_T_943,_T_944,_T_945}; // @[Cat.scala 30:58:@4904.4]
  assign _T_948 = imm_itype[11]; // @[InstDecoder.scala 153:43:@4905.4]
  assign _T_952 = _T_948 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@4907.4]
  assign _T_954 = imm_stype[11]; // @[InstDecoder.scala 154:43:@4910.4]
  assign _T_958 = _T_954 ? 20'hfffff : 20'h0; // @[Bitwise.scala 72:12:@4912.4]
  assign _T_960 = imm_sbtype[11]; // @[InstDecoder.scala 155:44:@4915.4]
  assign _T_964 = _T_960 ? 19'h7ffff : 19'h0; // @[Bitwise.scala 72:12:@4917.4]
  assign _T_966 = {_T_964,_T_936,_T_937,_T_938,_T_939}; // @[Cat.scala 30:58:@4918.4]
  assign _T_974 = imm_ujtype[19]; // @[InstDecoder.scala 157:44:@4924.4]
  assign _T_978 = _T_974 ? 11'h7ff : 11'h0; // @[Bitwise.scala 72:12:@4926.4]
  assign _T_980 = {_T_978,_T_936,_T_943,_T_944,_T_945}; // @[Cat.scala 30:58:@4927.4]
  assign io_cinfo_br_type = _T_14 ? 4'h0 : _T_308; // @[InstDecoder.scala 115:20:@4840.4]
  assign io_cinfo_op1_sel = _T_14 ? 2'h0 : _T_357; // @[InstDecoder.scala 116:20:@4841.4]
  assign io_cinfo_op2_sel = _T_14 ? 3'h1 : _T_406; // @[InstDecoder.scala 117:20:@4842.4]
  assign io_cinfo_rs1_oen = _T_14 ? 1'h1 : _T_455; // @[InstDecoder.scala 118:20:@4843.4]
  assign io_cinfo_rs2_oen = _T_14 ? 1'h0 : _T_504; // @[InstDecoder.scala 119:20:@4844.4]
  assign io_cinfo_alu_fun = _T_14 ? 4'h0 : _T_553; // @[InstDecoder.scala 120:20:@4845.4]
  assign io_cinfo_wb_sel = _T_14 ? 2'h1 : _T_602; // @[InstDecoder.scala 121:20:@4846.4]
  assign io_cinfo_rf_wen = _T_14 ? 1'h1 : _T_651; // @[InstDecoder.scala 122:20:@4847.4]
  assign io_cinfo_mem_en = _T_14 ? 1'h1 : _T_700; // @[InstDecoder.scala 123:20:@4848.4]
  assign io_cinfo_mem_fcn = _T_14 ? 1'h0 : _T_749; // @[InstDecoder.scala 124:20:@4849.4]
  assign io_cinfo_mem_typ = _T_14 ? 3'h3 : _T_798; // @[InstDecoder.scala 125:20:@4850.4]
  assign io_cinfo_csr_cmd = _T_14 ? 3'h0 : _T_847; // @[InstDecoder.scala 126:20:@4851.4]
  assign io_cinfo_illegal = signals_0 == 1'h0; // @[InstDecoder.scala 127:20:@4853.4]
  assign io_cinfo_fencei = _T_14 ? 1'h0 : _T_896; // @[InstDecoder.scala 128:20:@4854.4]
  assign io_cinfo_is_branch = func == 5'h18; // @[InstDecoder.scala 139:22:@4863.4]
  assign io_cinfo_push = _T_908 & _T_913; // @[InstDecoder.scala 141:17:@4871.4]
  assign io_cinfo_pop = _T_923 & _T_932; // @[InstDecoder.scala 142:16:@4885.4]
  assign io_cinfo_rs1_addr = io_inst[19:15]; // @[InstDecoder.scala 130:21:@4856.4]
  assign io_cinfo_rs2_addr = io_inst[24:20]; // @[InstDecoder.scala 131:21:@4858.4]
  assign io_cinfo_wbaddr = io_inst[11:7]; // @[InstDecoder.scala 132:21:@4860.4]
  assign io_dinfo_imm_i = {_T_952,imm_itype}; // @[InstDecoder.scala 153:19:@4909.4]
  assign io_dinfo_imm_s = {_T_958,imm_stype}; // @[InstDecoder.scala 154:19:@4914.4]
  assign io_dinfo_imm_sb = {_T_966,1'h0}; // @[InstDecoder.scala 155:19:@4920.4]
  assign io_dinfo_imm_u = {imm_utype,12'h0}; // @[InstDecoder.scala 156:19:@4923.4]
  assign io_dinfo_imm_uj = {_T_980,1'h0}; // @[InstDecoder.scala 157:19:@4929.4]
  assign io_dinfo_imm_z = {27'h0,_T_899}; // @[InstDecoder.scala 158:19:@4933.4]
endmodule
module Regfile( // @[:@4935.2]
  input         clock, // @[:@4936.4]
  input  [4:0]  io_rs1_addr, // @[:@4938.4]
  output [31:0] io_rs1_data, // @[:@4938.4]
  input  [4:0]  io_rs2_addr, // @[:@4938.4]
  output [31:0] io_rs2_data, // @[:@4938.4]
  input  [4:0]  io_waddr, // @[:@4938.4]
  input  [31:0] io_wdata, // @[:@4938.4]
  input         io_wen // @[:@4938.4]
);
  reg [31:0] regfile [0:31]; // @[Regfile.scala 24:21:@4940.4]
  reg [31:0] _RAND_0;
  wire [31:0] regfile__T_27_data; // @[Regfile.scala 24:21:@4940.4]
  wire [4:0] regfile__T_27_addr; // @[Regfile.scala 24:21:@4940.4]
  wire [31:0] regfile__T_32_data; // @[Regfile.scala 24:21:@4940.4]
  wire [4:0] regfile__T_32_addr; // @[Regfile.scala 24:21:@4940.4]
  wire [31:0] regfile__T_24_data; // @[Regfile.scala 24:21:@4940.4]
  wire [4:0] regfile__T_24_addr; // @[Regfile.scala 24:21:@4940.4]
  wire  regfile__T_24_mask; // @[Regfile.scala 24:21:@4940.4]
  wire  regfile__T_24_en; // @[Regfile.scala 24:21:@4940.4]
  wire  _T_22; // @[Regfile.scala 26:30:@4941.4]
  wire  _T_26; // @[Regfile.scala 30:35:@4947.4]
  wire  _T_31; // @[Regfile.scala 31:35:@4951.4]
  assign regfile__T_27_addr = io_rs1_addr;
  assign regfile__T_27_data = regfile[regfile__T_27_addr]; // @[Regfile.scala 24:21:@4940.4]
  assign regfile__T_32_addr = io_rs2_addr;
  assign regfile__T_32_data = regfile[regfile__T_32_addr]; // @[Regfile.scala 24:21:@4940.4]
  assign regfile__T_24_data = io_wdata;
  assign regfile__T_24_addr = io_waddr;
  assign regfile__T_24_mask = 1'h1;
  assign regfile__T_24_en = io_wen & _T_22;
  assign _T_22 = io_waddr != 5'h0; // @[Regfile.scala 26:30:@4941.4]
  assign _T_26 = io_rs1_addr != 5'h0; // @[Regfile.scala 30:35:@4947.4]
  assign _T_31 = io_rs2_addr != 5'h0; // @[Regfile.scala 31:35:@4951.4]
  assign io_rs1_data = _T_26 ? regfile__T_27_data : 32'h0; // @[Regfile.scala 30:16:@4950.4]
  assign io_rs2_data = _T_31 ? regfile__T_32_data : 32'h0; // @[Regfile.scala 31:16:@4954.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  _RAND_0 = {1{`RANDOM}};
  `ifdef RANDOMIZE_MEM_INIT
  for (initvar = 0; initvar < 32; initvar = initvar+1)
    regfile[initvar] = _RAND_0[31:0];
  `endif // RANDOMIZE_MEM_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if(regfile__T_24_en & regfile__T_24_mask) begin
      regfile[regfile__T_24_addr] <= regfile__T_24_data; // @[Regfile.scala 24:21:@4940.4]
    end
  end
endmodule
module ALU( // @[:@4956.2]
  input  [31:0] io_op1, // @[:@4959.4]
  input  [31:0] io_op2, // @[:@4959.4]
  input  [31:0] io_pc, // @[:@4959.4]
  input  [3:0]  io_ctrl_fun, // @[:@4959.4]
  input  [3:0]  io_ctrl_br_type, // @[:@4959.4]
  input  [1:0]  io_ctrl_wb_sel, // @[:@4959.4]
  output [1:0]  io_ctrl_pc_sel, // @[:@4959.4]
  input  [31:0] io_rs2_data, // @[:@4959.4]
  output [31:0] io_result, // @[:@4959.4]
  output [31:0] io_target_brjmp, // @[:@4959.4]
  output [31:0] io_target_jpreg, // @[:@4959.4]
  output [31:0] io_target_conti // @[:@4959.4]
);
  wire [4:0] alu_shamt; // @[ALU.scala 32:32:@4961.4]
  wire [32:0] _T_25; // @[ALU.scala 33:34:@4962.4]
  wire [31:0] add_result; // @[ALU.scala 33:34:@4963.4]
  wire  _T_29; // @[ALU.scala 38:18:@4966.4]
  wire  _T_30; // @[ALU.scala 39:18:@4967.4]
  wire [32:0] _T_31; // @[ALU.scala 39:44:@4968.4]
  wire [32:0] _T_32; // @[ALU.scala 39:44:@4969.4]
  wire [31:0] _T_33; // @[ALU.scala 39:44:@4970.4]
  wire  _T_34; // @[ALU.scala 40:18:@4971.4]
  wire [31:0] _T_35; // @[ALU.scala 40:44:@4972.4]
  wire  _T_36; // @[ALU.scala 41:18:@4973.4]
  wire [31:0] _T_37; // @[ALU.scala 41:44:@4974.4]
  wire  _T_38; // @[ALU.scala 42:18:@4975.4]
  wire [31:0] _T_39; // @[ALU.scala 42:44:@4976.4]
  wire  _T_40; // @[ALU.scala 43:18:@4977.4]
  wire [31:0] _T_41; // @[ALU.scala 43:44:@4978.4]
  wire [31:0] _T_42; // @[ALU.scala 43:60:@4979.4]
  wire  _T_43; // @[ALU.scala 43:51:@4980.4]
  wire  _T_44; // @[ALU.scala 44:18:@4981.4]
  wire  _T_45; // @[ALU.scala 44:44:@4982.4]
  wire  _T_46; // @[ALU.scala 45:18:@4983.4]
  wire [62:0] _GEN_0; // @[ALU.scala 45:44:@4984.4]
  wire [62:0] _T_47; // @[ALU.scala 45:44:@4984.4]
  wire [31:0] _T_48; // @[ALU.scala 45:57:@4985.4]
  wire  _T_49; // @[ALU.scala 46:18:@4986.4]
  wire [31:0] _T_51; // @[ALU.scala 46:51:@4988.4]
  wire [31:0] _T_52; // @[ALU.scala 46:65:@4989.4]
  wire  _T_53; // @[ALU.scala 47:18:@4990.4]
  wire [31:0] _T_54; // @[ALU.scala 47:44:@4991.4]
  wire  _T_55; // @[ALU.scala 48:18:@4992.4]
  wire  _T_56; // @[ALU.scala 49:18:@4993.4]
  wire [31:0] _T_57; // @[Mux.scala 61:16:@4994.4]
  wire [31:0] _T_58; // @[Mux.scala 61:16:@4995.4]
  wire [31:0] _T_59; // @[Mux.scala 61:16:@4996.4]
  wire [31:0] _T_60; // @[Mux.scala 61:16:@4997.4]
  wire [31:0] _T_61; // @[Mux.scala 61:16:@4998.4]
  wire [31:0] _T_62; // @[Mux.scala 61:16:@4999.4]
  wire [31:0] _T_63; // @[Mux.scala 61:16:@5000.4]
  wire [31:0] _T_64; // @[Mux.scala 61:16:@5001.4]
  wire [31:0] _T_65; // @[Mux.scala 61:16:@5002.4]
  wire [31:0] _T_66; // @[Mux.scala 61:16:@5003.4]
  wire [31:0] _T_67; // @[Mux.scala 61:16:@5004.4]
  wire [31:0] result; // @[Mux.scala 61:16:@5005.4]
  wire [32:0] _T_69; // @[ALU.scala 52:31:@5007.4]
  wire [30:0] _T_71; // @[ALU.scala 53:39:@5010.4]
  wire [32:0] _T_75; // @[ALU.scala 54:31:@5013.4]
  wire  _T_77; // @[ALU.scala 55:40:@5016.4]
  wire  br_eq; // @[ALU.scala 57:29:@5019.4]
  wire [31:0] _T_80; // @[ALU.scala 58:50:@5021.4]
  wire  br_lt; // @[ALU.scala 58:36:@5022.4]
  wire  br_ltu; // @[ALU.scala 59:36:@5023.4]
  wire  _T_81; // @[ALU.scala 63:25:@5024.4]
  wire  _T_82; // @[ALU.scala 64:25:@5025.4]
  wire  _T_84; // @[ALU.scala 64:41:@5026.4]
  wire [1:0] _T_85; // @[ALU.scala 64:40:@5027.4]
  wire  _T_86; // @[ALU.scala 65:25:@5028.4]
  wire [1:0] _T_87; // @[ALU.scala 65:40:@5029.4]
  wire  _T_88; // @[ALU.scala 66:25:@5030.4]
  wire  _T_90; // @[ALU.scala 66:41:@5031.4]
  wire [1:0] _T_91; // @[ALU.scala 66:40:@5032.4]
  wire  _T_92; // @[ALU.scala 67:25:@5033.4]
  wire  _T_94; // @[ALU.scala 67:41:@5034.4]
  wire [1:0] _T_95; // @[ALU.scala 67:40:@5035.4]
  wire  _T_96; // @[ALU.scala 68:25:@5036.4]
  wire [1:0] _T_97; // @[ALU.scala 68:40:@5037.4]
  wire  _T_98; // @[ALU.scala 69:25:@5038.4]
  wire [1:0] _T_99; // @[ALU.scala 69:40:@5039.4]
  wire  _T_100; // @[ALU.scala 70:25:@5040.4]
  wire  _T_101; // @[ALU.scala 71:25:@5041.4]
  wire [1:0] _T_102; // @[ALU.scala 71:8:@5042.4]
  wire [1:0] _T_103; // @[ALU.scala 70:8:@5043.4]
  wire [1:0] _T_104; // @[ALU.scala 69:8:@5044.4]
  wire [1:0] _T_105; // @[ALU.scala 68:8:@5045.4]
  wire [1:0] _T_106; // @[ALU.scala 67:8:@5046.4]
  wire [1:0] _T_107; // @[ALU.scala 66:8:@5047.4]
  wire [1:0] _T_108; // @[ALU.scala 65:8:@5048.4]
  wire [1:0] _T_109; // @[ALU.scala 64:8:@5049.4]
  assign alu_shamt = io_op2[4:0]; // @[ALU.scala 32:32:@4961.4]
  assign _T_25 = io_op1 + io_op2; // @[ALU.scala 33:34:@4962.4]
  assign add_result = io_op1 + io_op2; // @[ALU.scala 33:34:@4963.4]
  assign _T_29 = io_ctrl_fun == 4'h0; // @[ALU.scala 38:18:@4966.4]
  assign _T_30 = io_ctrl_fun == 4'h1; // @[ALU.scala 39:18:@4967.4]
  assign _T_31 = io_op1 - io_op2; // @[ALU.scala 39:44:@4968.4]
  assign _T_32 = $unsigned(_T_31); // @[ALU.scala 39:44:@4969.4]
  assign _T_33 = _T_32[31:0]; // @[ALU.scala 39:44:@4970.4]
  assign _T_34 = io_ctrl_fun == 4'h5; // @[ALU.scala 40:18:@4971.4]
  assign _T_35 = io_op1 & io_op2; // @[ALU.scala 40:44:@4972.4]
  assign _T_36 = io_ctrl_fun == 4'h6; // @[ALU.scala 41:18:@4973.4]
  assign _T_37 = io_op1 | io_op2; // @[ALU.scala 41:44:@4974.4]
  assign _T_38 = io_ctrl_fun == 4'h7; // @[ALU.scala 42:18:@4975.4]
  assign _T_39 = io_op1 ^ io_op2; // @[ALU.scala 42:44:@4976.4]
  assign _T_40 = io_ctrl_fun == 4'h8; // @[ALU.scala 43:18:@4977.4]
  assign _T_41 = $signed(io_op1); // @[ALU.scala 43:44:@4978.4]
  assign _T_42 = $signed(io_op2); // @[ALU.scala 43:60:@4979.4]
  assign _T_43 = $signed(_T_41) < $signed(_T_42); // @[ALU.scala 43:51:@4980.4]
  assign _T_44 = io_ctrl_fun == 4'h9; // @[ALU.scala 44:18:@4981.4]
  assign _T_45 = io_op1 < io_op2; // @[ALU.scala 44:44:@4982.4]
  assign _T_46 = io_ctrl_fun == 4'h2; // @[ALU.scala 45:18:@4983.4]
  assign _GEN_0 = {{31'd0}, io_op1}; // @[ALU.scala 45:44:@4984.4]
  assign _T_47 = _GEN_0 << alu_shamt; // @[ALU.scala 45:44:@4984.4]
  assign _T_48 = _T_47[31:0]; // @[ALU.scala 45:57:@4985.4]
  assign _T_49 = io_ctrl_fun == 4'h4; // @[ALU.scala 46:18:@4986.4]
  assign _T_51 = $signed(_T_41) >>> alu_shamt; // @[ALU.scala 46:51:@4988.4]
  assign _T_52 = $unsigned(_T_51); // @[ALU.scala 46:65:@4989.4]
  assign _T_53 = io_ctrl_fun == 4'h3; // @[ALU.scala 47:18:@4990.4]
  assign _T_54 = io_op1 >> alu_shamt; // @[ALU.scala 47:44:@4991.4]
  assign _T_55 = io_ctrl_fun == 4'ha; // @[ALU.scala 48:18:@4992.4]
  assign _T_56 = io_ctrl_fun == 4'hb; // @[ALU.scala 49:18:@4993.4]
  assign _T_57 = _T_56 ? io_op2 : 32'h0; // @[Mux.scala 61:16:@4994.4]
  assign _T_58 = _T_55 ? io_op1 : _T_57; // @[Mux.scala 61:16:@4995.4]
  assign _T_59 = _T_53 ? _T_54 : _T_58; // @[Mux.scala 61:16:@4996.4]
  assign _T_60 = _T_49 ? _T_52 : _T_59; // @[Mux.scala 61:16:@4997.4]
  assign _T_61 = _T_46 ? _T_48 : _T_60; // @[Mux.scala 61:16:@4998.4]
  assign _T_62 = _T_44 ? {{31'd0}, _T_45} : _T_61; // @[Mux.scala 61:16:@4999.4]
  assign _T_63 = _T_40 ? {{31'd0}, _T_43} : _T_62; // @[Mux.scala 61:16:@5000.4]
  assign _T_64 = _T_38 ? _T_39 : _T_63; // @[Mux.scala 61:16:@5001.4]
  assign _T_65 = _T_36 ? _T_37 : _T_64; // @[Mux.scala 61:16:@5002.4]
  assign _T_66 = _T_34 ? _T_35 : _T_65; // @[Mux.scala 61:16:@5003.4]
  assign _T_67 = _T_30 ? _T_33 : _T_66; // @[Mux.scala 61:16:@5004.4]
  assign result = _T_29 ? add_result : _T_67; // @[Mux.scala 61:16:@5005.4]
  assign _T_69 = io_pc + io_op2; // @[ALU.scala 52:31:@5007.4]
  assign _T_71 = add_result[31:1]; // @[ALU.scala 53:39:@5010.4]
  assign _T_75 = io_pc + 32'h4; // @[ALU.scala 54:31:@5013.4]
  assign _T_77 = io_ctrl_wb_sel == 2'h2; // @[ALU.scala 55:40:@5016.4]
  assign br_eq = io_op1 == io_rs2_data; // @[ALU.scala 57:29:@5019.4]
  assign _T_80 = $signed(io_rs2_data); // @[ALU.scala 58:50:@5021.4]
  assign br_lt = $signed(_T_41) < $signed(_T_80); // @[ALU.scala 58:36:@5022.4]
  assign br_ltu = io_op1 < io_rs2_data; // @[ALU.scala 59:36:@5023.4]
  assign _T_81 = io_ctrl_br_type == 4'h0; // @[ALU.scala 63:25:@5024.4]
  assign _T_82 = io_ctrl_br_type == 4'h1; // @[ALU.scala 64:25:@5025.4]
  assign _T_84 = br_eq == 1'h0; // @[ALU.scala 64:41:@5026.4]
  assign _T_85 = _T_84 ? 2'h1 : 2'h0; // @[ALU.scala 64:40:@5027.4]
  assign _T_86 = io_ctrl_br_type == 4'h2; // @[ALU.scala 65:25:@5028.4]
  assign _T_87 = br_eq ? 2'h1 : 2'h0; // @[ALU.scala 65:40:@5029.4]
  assign _T_88 = io_ctrl_br_type == 4'h3; // @[ALU.scala 66:25:@5030.4]
  assign _T_90 = br_lt == 1'h0; // @[ALU.scala 66:41:@5031.4]
  assign _T_91 = _T_90 ? 2'h1 : 2'h0; // @[ALU.scala 66:40:@5032.4]
  assign _T_92 = io_ctrl_br_type == 4'h4; // @[ALU.scala 67:25:@5033.4]
  assign _T_94 = br_ltu == 1'h0; // @[ALU.scala 67:41:@5034.4]
  assign _T_95 = _T_94 ? 2'h1 : 2'h0; // @[ALU.scala 67:40:@5035.4]
  assign _T_96 = io_ctrl_br_type == 4'h5; // @[ALU.scala 68:25:@5036.4]
  assign _T_97 = br_lt ? 2'h1 : 2'h0; // @[ALU.scala 68:40:@5037.4]
  assign _T_98 = io_ctrl_br_type == 4'h6; // @[ALU.scala 69:25:@5038.4]
  assign _T_99 = br_ltu ? 2'h1 : 2'h0; // @[ALU.scala 69:40:@5039.4]
  assign _T_100 = io_ctrl_br_type == 4'h7; // @[ALU.scala 70:25:@5040.4]
  assign _T_101 = io_ctrl_br_type == 4'h8; // @[ALU.scala 71:25:@5041.4]
  assign _T_102 = _T_101 ? 2'h2 : 2'h0; // @[ALU.scala 71:8:@5042.4]
  assign _T_103 = _T_100 ? 2'h1 : _T_102; // @[ALU.scala 70:8:@5043.4]
  assign _T_104 = _T_98 ? _T_99 : _T_103; // @[ALU.scala 69:8:@5044.4]
  assign _T_105 = _T_96 ? _T_97 : _T_104; // @[ALU.scala 68:8:@5045.4]
  assign _T_106 = _T_92 ? _T_95 : _T_105; // @[ALU.scala 67:8:@5046.4]
  assign _T_107 = _T_88 ? _T_91 : _T_106; // @[ALU.scala 66:8:@5047.4]
  assign _T_108 = _T_86 ? _T_87 : _T_107; // @[ALU.scala 65:8:@5048.4]
  assign _T_109 = _T_82 ? _T_85 : _T_108; // @[ALU.scala 64:8:@5049.4]
  assign io_ctrl_pc_sel = _T_81 ? 2'h0 : _T_109; // @[ALU.scala 62:18:@5051.4]
  assign io_result = _T_77 ? io_target_conti : result; // @[ALU.scala 55:18:@5018.4]
  assign io_target_brjmp = io_pc + io_op2; // @[ALU.scala 52:22:@5009.4]
  assign io_target_jpreg = {_T_71,1'h0}; // @[ALU.scala 53:22:@5012.4]
  assign io_target_conti = io_pc + 32'h4; // @[ALU.scala 54:22:@5015.4]
endmodule
module BackEnd( // @[:@5053.2]
  input         clock, // @[:@5054.4]
  input         reset, // @[:@5055.4]
  output        io_mem_req_valid, // @[:@5056.4]
  output [31:0] io_mem_req_bits_addr, // @[:@5056.4]
  output [31:0] io_mem_req_bits_data, // @[:@5056.4]
  output        io_mem_req_bits_fcn, // @[:@5056.4]
  output [2:0]  io_mem_req_bits_typ, // @[:@5056.4]
  input         io_mem_resp_valid, // @[:@5056.4]
  input  [31:0] io_mem_resp_bits_data, // @[:@5056.4]
  output [31:0] io_cyc, // @[:@5056.4]
  output        io_front_xcpt_valid, // @[:@5056.4]
  output [31:0] io_front_xcpt_bits, // @[:@5056.4]
  output        io_front_kill, // @[:@5056.4]
  output        io_front_fence, // @[:@5056.4]
  output        io_front_forward, // @[:@5056.4]
  output        io_front_ras_pop, // @[:@5056.4]
  output        io_front_ras_push_valid, // @[:@5056.4]
  output [31:0] io_front_ras_push_bits, // @[:@5056.4]
  output [31:0] io_front_fb_pc, // @[:@5056.4]
  output [1:0]  io_front_fb_type, // @[:@5056.4]
  output        io_front_feedBack_valid, // @[:@5056.4]
  output        io_front_feedBack_bits_redirect, // @[:@5056.4]
  output [31:0] io_front_feedBack_bits_tgt, // @[:@5056.4]
  input         io_front_inst_valid, // @[:@5056.4]
  input  [31:0] io_front_inst_bits, // @[:@5056.4]
  input  [31:0] io_front_pc, // @[:@5056.4]
  input  [31:0] io_front_pred // @[:@5056.4]
);
  wire  csr_clock; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_reset; // @[BackEnd.scala 86:19:@5058.4]
  wire [2:0] csr_io_rw_cmd; // @[BackEnd.scala 86:19:@5058.4]
  wire [11:0] csr_io_rw_addr; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_rw_rdata; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_rw_wdata; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_eret; // @[BackEnd.scala 86:19:@5058.4]
  wire [1:0] csr_io_status_prv; // @[BackEnd.scala 86:19:@5058.4]
  wire [13:0] csr_io_status_unimp5; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_status_mprv; // @[BackEnd.scala 86:19:@5058.4]
  wire [1:0] csr_io_status_unimp4; // @[BackEnd.scala 86:19:@5058.4]
  wire [1:0] csr_io_status_mpp; // @[BackEnd.scala 86:19:@5058.4]
  wire [2:0] csr_io_status_unimp3; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_status_mpie; // @[BackEnd.scala 86:19:@5058.4]
  wire [2:0] csr_io_status_unimp2; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_status_mie; // @[BackEnd.scala 86:19:@5058.4]
  wire [2:0] csr_io_status_unimp1; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_xcpt; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_cause; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_tval; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_evec; // @[BackEnd.scala 86:19:@5058.4]
  wire  csr_io_illegal; // @[BackEnd.scala 86:19:@5058.4]
  wire [1:0] csr_io_retire; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_pc; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] csr_io_time; // @[BackEnd.scala 86:19:@5058.4]
  wire [31:0] InstDecoder_io_inst; // @[BackEnd.scala 91:25:@5064.4]
  wire [3:0] InstDecoder_io_cinfo_br_type; // @[BackEnd.scala 91:25:@5064.4]
  wire [1:0] InstDecoder_io_cinfo_op1_sel; // @[BackEnd.scala 91:25:@5064.4]
  wire [2:0] InstDecoder_io_cinfo_op2_sel; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 91:25:@5064.4]
  wire [3:0] InstDecoder_io_cinfo_alu_fun; // @[BackEnd.scala 91:25:@5064.4]
  wire [1:0] InstDecoder_io_cinfo_wb_sel; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_rf_wen; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_mem_en; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_mem_fcn; // @[BackEnd.scala 91:25:@5064.4]
  wire [2:0] InstDecoder_io_cinfo_mem_typ; // @[BackEnd.scala 91:25:@5064.4]
  wire [2:0] InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_illegal; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_fencei; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_is_branch; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_push; // @[BackEnd.scala 91:25:@5064.4]
  wire  InstDecoder_io_cinfo_pop; // @[BackEnd.scala 91:25:@5064.4]
  wire [4:0] InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 91:25:@5064.4]
  wire [4:0] InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 91:25:@5064.4]
  wire [4:0] InstDecoder_io_cinfo_wbaddr; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_i; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_s; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_sb; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_u; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_uj; // @[BackEnd.scala 91:25:@5064.4]
  wire [31:0] InstDecoder_io_dinfo_imm_z; // @[BackEnd.scala 91:25:@5064.4]
  wire  regfile_clock; // @[BackEnd.scala 122:23:@5095.4]
  wire [4:0] regfile_io_rs1_addr; // @[BackEnd.scala 122:23:@5095.4]
  wire [31:0] regfile_io_rs1_data; // @[BackEnd.scala 122:23:@5095.4]
  wire [4:0] regfile_io_rs2_addr; // @[BackEnd.scala 122:23:@5095.4]
  wire [31:0] regfile_io_rs2_data; // @[BackEnd.scala 122:23:@5095.4]
  wire [4:0] regfile_io_waddr; // @[BackEnd.scala 122:23:@5095.4]
  wire [31:0] regfile_io_wdata; // @[BackEnd.scala 122:23:@5095.4]
  wire  regfile_io_wen; // @[BackEnd.scala 122:23:@5095.4]
  wire [31:0] ALU_io_op1; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_op2; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_pc; // @[BackEnd.scala 193:19:@5203.4]
  wire [3:0] ALU_io_ctrl_fun; // @[BackEnd.scala 193:19:@5203.4]
  wire [3:0] ALU_io_ctrl_br_type; // @[BackEnd.scala 193:19:@5203.4]
  wire [1:0] ALU_io_ctrl_wb_sel; // @[BackEnd.scala 193:19:@5203.4]
  wire [1:0] ALU_io_ctrl_pc_sel; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_rs2_data; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_result; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_target_brjmp; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_target_jpreg; // @[BackEnd.scala 193:19:@5203.4]
  wire [31:0] ALU_io_target_conti; // @[BackEnd.scala 193:19:@5203.4]
  reg  exe_rf_wen; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_0;
  reg [4:0] exe_wbaddr; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_1;
  reg  exe_mem_en; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_2;
  reg [2:0] exe_csr_cmd; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_3;
  reg  exe_illegal; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_4;
  reg [31:0] exe_pc; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_5;
  reg [31:0] exe_inst; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_6;
  reg [31:0] exe_rs2_data; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_7;
  reg [1:0] exe_wb_sel; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_8;
  reg  exe_mem_fcn; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_9;
  reg [2:0] exe_mem_typ; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_10;
  reg  exe_fencei; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_11;
  reg [3:0] exe_br_type; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_12;
  reg  exe_branch; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_13;
  reg  exe_push; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_14;
  reg  exe_pop; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_15;
  reg [31:0] exe_pred; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_16;
  reg [31:0] exe_op1_data; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_17;
  reg [31:0] exe_op2_data; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_18;
  reg [3:0] exe_alu_fun; // @[BackEnd.scala 94:22:@5069.4]
  reg [31:0] _RAND_19;
  reg  exe_valid; // @[BackEnd.scala 95:26:@5070.4]
  reg [31:0] _RAND_20;
  reg  mem_rf_wen; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_21;
  reg [4:0] mem_wbaddr; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_22;
  reg  mem_mem_en; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_23;
  reg [2:0] mem_csr_cmd; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_24;
  reg  mem_illegal; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_25;
  reg [31:0] mem_pc; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_26;
  reg [31:0] mem_inst; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_27;
  reg [1:0] mem_wb_sel; // @[BackEnd.scala 97:22:@5072.4]
  reg [31:0] _RAND_28;
  reg  mem_valid; // @[BackEnd.scala 98:26:@5073.4]
  reg [31:0] _RAND_29;
  reg  wb_rf_wen; // @[BackEnd.scala 100:22:@5075.4]
  reg [31:0] _RAND_30;
  reg [4:0] wb_wbaddr; // @[BackEnd.scala 100:22:@5075.4]
  reg [31:0] _RAND_31;
  reg  wb_valid; // @[BackEnd.scala 101:26:@5076.4]
  reg [31:0] _RAND_32;
  reg [31:0] wb_wbdata; // @[BackEnd.scala 106:23:@5080.4]
  reg [31:0] _RAND_33;
  wire  dec_wire_rs1_oen; // @[BackEnd.scala 110:33:@5083.4]
  wire  dec_wire_rs2_oen; // @[BackEnd.scala 111:33:@5085.4]
  wire  dec_wire_fencei; // @[BackEnd.scala 112:33:@5087.4]
  wire  exe_wire_fencei; // @[BackEnd.scala 191:34:@5201.4]
  wire  _T_177; // @[BackEnd.scala 131:18:@5104.4]
  wire  _T_232; // @[BackEnd.scala 183:34:@5183.4]
  wire  _T_234; // @[BackEnd.scala 183:61:@5184.4]
  wire  exe_wire_rf_wen; // @[BackEnd.scala 183:47:@5185.4]
  wire  _T_178; // @[BackEnd.scala 131:42:@5105.4]
  wire  _T_179; // @[BackEnd.scala 132:18:@5106.4]
  wire  _T_329; // @[BackEnd.scala 267:35:@5329.4]
  wire  _T_331; // @[BackEnd.scala 267:62:@5330.4]
  wire  mem_wire_rf_wen; // @[BackEnd.scala 267:48:@5331.4]
  wire  _T_180; // @[BackEnd.scala 132:42:@5107.4]
  wire  _T_181; // @[BackEnd.scala 133:18:@5108.4]
  wire  _T_366; // @[BackEnd.scala 315:33:@5473.4]
  wire  _T_368; // @[BackEnd.scala 315:58:@5474.4]
  wire  wb_wire_rf_wen; // @[BackEnd.scala 315:45:@5475.4]
  wire  _T_182; // @[BackEnd.scala 133:42:@5109.4]
  wire [31:0] rf_rs1_data; // @[BackEnd.scala 123:25:@5098.4 BackEnd.scala 127:15:@5102.4]
  wire [31:0] _T_183; // @[Mux.scala 61:16:@5110.4]
  wire  _T_360; // @[BackEnd.scala 302:17:@5458.4]
  wire  _T_361; // @[BackEnd.scala 303:17:@5459.4]
  reg [31:0] mem_exe_out; // @[BackEnd.scala 239:25:@5290.4]
  reg [31:0] _RAND_34;
  wire [31:0] _T_362; // @[Mux.scala 61:16:@5460.4]
  wire [31:0] mem_wbdata; // @[Mux.scala 61:16:@5461.4]
  wire [31:0] _T_184; // @[Mux.scala 61:16:@5111.4]
  wire [31:0] exe_wbdata; // @[BackEnd.scala 104:24:@5078.4 BackEnd.scala 201:20:@5213.4]
  wire [31:0] dec_rs1_data; // @[Mux.scala 61:16:@5112.4]
  wire  _T_186; // @[BackEnd.scala 137:18:@5114.4]
  wire  _T_187; // @[BackEnd.scala 137:42:@5115.4]
  wire  _T_188; // @[BackEnd.scala 138:18:@5116.4]
  wire  _T_189; // @[BackEnd.scala 138:42:@5117.4]
  wire  _T_190; // @[BackEnd.scala 139:18:@5118.4]
  wire  _T_191; // @[BackEnd.scala 139:42:@5119.4]
  wire [31:0] rf_rs2_data; // @[BackEnd.scala 124:25:@5099.4 BackEnd.scala 128:15:@5103.4]
  wire [31:0] _T_192; // @[Mux.scala 61:16:@5120.4]
  wire [31:0] _T_193; // @[Mux.scala 61:16:@5121.4]
  wire [31:0] dec_rs2_data; // @[Mux.scala 61:16:@5122.4]
  wire  _T_195; // @[BackEnd.scala 143:24:@5124.4]
  wire  _T_196; // @[BackEnd.scala 144:24:@5125.4]
  wire [31:0] _T_197; // @[Mux.scala 61:16:@5126.4]
  wire [31:0] dec_op1_data; // @[Mux.scala 61:16:@5127.4]
  wire  _T_199; // @[BackEnd.scala 147:24:@5129.4]
  wire  _T_200; // @[BackEnd.scala 148:24:@5130.4]
  wire  _T_201; // @[BackEnd.scala 149:24:@5131.4]
  wire  _T_202; // @[BackEnd.scala 150:24:@5132.4]
  wire  _T_203; // @[BackEnd.scala 151:24:@5133.4]
  wire [31:0] _T_204; // @[Mux.scala 61:16:@5134.4]
  wire [31:0] _T_205; // @[Mux.scala 61:16:@5135.4]
  wire [31:0] _T_206; // @[Mux.scala 61:16:@5136.4]
  wire [31:0] _T_207; // @[Mux.scala 61:16:@5137.4]
  wire [31:0] dec_op2_data; // @[Mux.scala 61:16:@5138.4]
  wire  exe_wire_mem_en; // @[BackEnd.scala 184:34:@5187.4]
  wire  _T_430; // @[BackEnd.scala 325:60:@5541.4]
  wire  exe_load_inst; // @[BackEnd.scala 325:45:@5542.4]
  wire  _T_432; // @[BackEnd.scala 328:20:@5544.4]
  wire  _T_434; // @[BackEnd.scala 328:79:@5545.4]
  wire  _T_435; // @[BackEnd.scala 328:57:@5546.4]
  wire  _T_436; // @[BackEnd.scala 328:87:@5547.4]
  wire  _T_438; // @[BackEnd.scala 329:20:@5549.4]
  wire  _T_440; // @[BackEnd.scala 329:79:@5550.4]
  wire  _T_441; // @[BackEnd.scala 329:57:@5551.4]
  wire  _T_442; // @[BackEnd.scala 329:87:@5552.4]
  wire  _T_443; // @[BackEnd.scala 328:108:@5553.4]
  wire [2:0] exe_wire_csr_cmd; // @[BackEnd.scala 185:26:@5189.4]
  wire  _T_444; // @[BackEnd.scala 330:22:@5554.4]
  wire  stall_0; // @[BackEnd.scala 329:108:@5555.4]
  wire  mem_wire_mem_en; // @[BackEnd.scala 268:35:@5333.4]
  wire  _T_450; // @[BackEnd.scala 333:42:@5560.4]
  wire  _T_451; // @[BackEnd.scala 333:39:@5561.4]
  reg  mem_ma_load; // @[BackEnd.scala 241:25:@5292.4]
  reg [31:0] _RAND_35;
  wire  mem_wire_ma_load; // @[BackEnd.scala 271:36:@5339.4]
  reg  mem_ma_store; // @[BackEnd.scala 242:25:@5293.4]
  reg [31:0] _RAND_36;
  wire  mem_wire_ma_store; // @[BackEnd.scala 272:37:@5341.4]
  wire  mem_wire_ma_valid; // @[BackEnd.scala 273:41:@5343.4]
  wire  _T_453; // @[BackEnd.scala 333:64:@5562.4]
  wire  stall_2; // @[BackEnd.scala 333:61:@5563.4]
  wire  _T_213; // @[BackEnd.scala 153:51:@5142.4]
  wire  _T_214; // @[BackEnd.scala 153:48:@5143.4]
  wire  _T_215; // @[BackEnd.scala 153:70:@5144.4]
  wire  _T_223; // @[BackEnd.scala 157:34:@5153.8]
  wire  _T_224; // @[BackEnd.scala 157:31:@5154.8]
  wire  _T_225; // @[BackEnd.scala 161:44:@5158.8]
  wire  _T_226; // @[BackEnd.scala 161:75:@5159.8]
  wire  _T_227; // @[BackEnd.scala 161:54:@5160.8]
  wire  _T_229; // @[BackEnd.scala 162:26:@5161.8]
  wire  _T_230; // @[BackEnd.scala 161:86:@5162.8]
  wire [2:0] _T_231; // @[BackEnd.scala 161:24:@5163.8]
  wire  _GEN_0; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_1; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_2; // @[BackEnd.scala 156:54:@5152.6]
  wire [2:0] _GEN_3; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_4; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_5; // @[BackEnd.scala 156:54:@5152.6]
  wire [3:0] _GEN_6; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_7; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_8; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_9; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_10; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_11; // @[BackEnd.scala 156:54:@5152.6]
  wire [3:0] _GEN_12; // @[BackEnd.scala 156:54:@5152.6]
  wire [1:0] _GEN_13; // @[BackEnd.scala 156:54:@5152.6]
  wire [4:0] _GEN_14; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_15; // @[BackEnd.scala 156:54:@5152.6]
  wire [2:0] _GEN_16; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_17; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_18; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_19; // @[BackEnd.scala 156:54:@5152.6]
  wire [31:0] _GEN_20; // @[BackEnd.scala 156:54:@5152.6]
  wire  _GEN_21; // @[BackEnd.scala 153:94:@5145.4]
  wire [3:0] exe_wire_br_type; // @[BackEnd.scala 186:26:@5191.4]
  wire  exe_wire_branch; // @[BackEnd.scala 187:33:@5193.4]
  wire  exe_wire_push; // @[BackEnd.scala 188:33:@5195.4]
  wire  exe_wire_pop; // @[BackEnd.scala 189:33:@5197.4]
  reg  _T_248; // @[BackEnd.scala 72:27:@5215.4]
  reg [31:0] _RAND_37;
  wire  _GEN_42; // @[BackEnd.scala 74:20:@5220.6]
  wire  _GEN_43; // @[BackEnd.scala 73:20:@5216.4]
  reg  _T_256; // @[BackEnd.scala 72:27:@5226.4]
  reg [31:0] _RAND_38;
  wire  _GEN_44; // @[BackEnd.scala 74:20:@5231.6]
  wire  _GEN_45; // @[BackEnd.scala 73:20:@5227.4]
  wire  _T_260; // @[BackEnd.scala 208:25:@5237.4]
  wire  _T_261; // @[BackEnd.scala 209:25:@5238.4]
  wire [31:0] _T_262; // @[BackEnd.scala 209:8:@5239.4]
  wire [31:0] next_pc; // @[BackEnd.scala 208:8:@5240.4]
  wire [1:0] _T_266; // @[BackEnd.scala 215:10:@5242.4]
  wire  _T_268; // @[BackEnd.scala 217:53:@5245.4]
  reg  _T_273; // @[BackEnd.scala 72:27:@5247.4]
  reg [31:0] _RAND_39;
  wire  _GEN_46; // @[BackEnd.scala 74:20:@5252.6]
  wire  _GEN_47; // @[BackEnd.scala 73:20:@5248.4]
  wire  _T_281; // @[BackEnd.scala 221:42:@5263.4]
  wire  mispredict; // @[BackEnd.scala 221:55:@5264.4]
  wire [1:0] _T_283; // @[BackEnd.scala 224:45:@5266.4]
  wire  _T_286; // @[BackEnd.scala 225:22:@5267.4]
  wire [1:0] _T_288; // @[BackEnd.scala 226:22:@5268.4]
  wire  _T_290; // @[BackEnd.scala 226:28:@5269.4]
  wire  _T_291; // @[Mux.scala 46:19:@5270.4]
  wire  _T_292; // @[Mux.scala 46:16:@5271.4]
  wire  _T_293; // @[Mux.scala 46:19:@5272.4]
  wire  exe_wire_ma_valid; // @[Mux.scala 46:16:@5273.4]
  wire  exe_wire_ma_load; // @[BackEnd.scala 228:46:@5276.4]
  wire  exe_wire_ma_store; // @[BackEnd.scala 229:46:@5279.4]
  wire  _T_300; // @[BackEnd.scala 232:46:@5281.4]
  wire  _T_301; // @[BackEnd.scala 232:43:@5282.4]
  wire  _T_303; // @[BackEnd.scala 232:68:@5283.4]
  reg [31:0] mem_jpnpc; // @[BackEnd.scala 240:25:@5291.4]
  reg [31:0] _RAND_40;
  wire  _T_312; // @[BackEnd.scala 243:47:@5296.4]
  wire [31:0] _T_320; // @[Bitwise.scala 72:12:@5320.8]
  wire [31:0] _T_321; // @[BackEnd.scala 262:70:@5321.8]
  wire [31:0] _T_326; // @[Bitwise.scala 72:12:@5324.8]
  wire [31:0] _T_327; // @[BackEnd.scala 263:74:@5325.8]
  wire [31:0] _T_328; // @[BackEnd.scala 262:90:@5326.8]
  wire  _GEN_48; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_49; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_50; // @[BackEnd.scala 245:34:@5302.6]
  wire [2:0] _GEN_51; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_52; // @[BackEnd.scala 245:34:@5302.6]
  wire [31:0] _GEN_53; // @[BackEnd.scala 245:34:@5302.6]
  wire [31:0] _GEN_54; // @[BackEnd.scala 245:34:@5302.6]
  wire [1:0] _GEN_55; // @[BackEnd.scala 245:34:@5302.6]
  wire [4:0] _GEN_56; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_60; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_61; // @[BackEnd.scala 245:34:@5302.6]
  wire [31:0] _GEN_62; // @[BackEnd.scala 245:34:@5302.6]
  wire [31:0] _GEN_63; // @[BackEnd.scala 245:34:@5302.6]
  wire  _GEN_64; // @[BackEnd.scala 243:71:@5297.4]
  wire  mem_wire_illegal; // @[BackEnd.scala 270:36:@5337.4]
  wire [1:0] _T_340; // @[BackEnd.scala 281:32:@5439.4]
  wire  _T_342; // @[BackEnd.scala 281:38:@5440.4]
  wire  ma_jump; // @[BackEnd.scala 281:42:@5441.4]
  wire  _T_344; // @[BackEnd.scala 283:57:@5443.4]
  wire [1:0] _T_351; // @[Mux.scala 61:16:@5446.4]
  wire [2:0] _T_352; // @[Mux.scala 61:16:@5447.4]
  wire [2:0] _T_353; // @[Mux.scala 61:16:@5448.4]
  wire [2:0] _T_354; // @[Mux.scala 61:16:@5449.4]
  wire [31:0] _T_356; // @[Mux.scala 61:16:@5451.4]
  wire [31:0] _T_357; // @[Mux.scala 61:16:@5452.4]
  wire  _GEN_80; // @[BackEnd.scala 305:50:@5464.4]
  reg  _T_459; // @[BackEnd.scala 72:27:@5566.4]
  reg [31:0] _RAND_41;
  wire  _GEN_84; // @[BackEnd.scala 74:20:@5571.6]
  wire  _GEN_85; // @[BackEnd.scala 73:20:@5567.4]
  wire [2:0] _T_464; // @[BackEnd.scala 336:32:@5577.4]
  wire  _T_466; // @[BackEnd.scala 336:39:@5578.4]
  wire [7:0] _T_472; // @[BackEnd.scala 345:10:@5581.4]
  wire [7:0] _T_473; // @[BackEnd.scala 344:10:@5582.4]
  wire  _T_481; // @[BackEnd.scala 348:27:@5585.4]
  wire  _T_484; // @[BackEnd.scala 349:27:@5586.4]
  wire [7:0] _T_487; // @[BackEnd.scala 349:10:@5587.4]
  wire [7:0] _T_488; // @[BackEnd.scala 348:10:@5588.4]
  wire [7:0] _T_489; // @[BackEnd.scala 347:10:@5589.4]
  wire [7:0] _T_490; // @[BackEnd.scala 346:10:@5590.4]
  wire [7:0] _T_493; // @[BackEnd.scala 350:10:@5591.4]
  wire  _T_495; // @[BackEnd.scala 351:34:@5592.4]
  wire  _T_496; // @[BackEnd.scala 351:31:@5593.4]
  wire [31:0] _T_497; // @[BackEnd.scala 351:10:@5594.4]
  wire  _T_500; // @[BackEnd.scala 339:9:@5596.4]
  wire  _T_504; // @[BackEnd.scala 368:24:@5608.6]
  CSRFile csr ( // @[BackEnd.scala 86:19:@5058.4]
    .clock(csr_clock),
    .reset(csr_reset),
    .io_rw_cmd(csr_io_rw_cmd),
    .io_rw_addr(csr_io_rw_addr),
    .io_rw_rdata(csr_io_rw_rdata),
    .io_rw_wdata(csr_io_rw_wdata),
    .io_eret(csr_io_eret),
    .io_status_prv(csr_io_status_prv),
    .io_status_unimp5(csr_io_status_unimp5),
    .io_status_mprv(csr_io_status_mprv),
    .io_status_unimp4(csr_io_status_unimp4),
    .io_status_mpp(csr_io_status_mpp),
    .io_status_unimp3(csr_io_status_unimp3),
    .io_status_mpie(csr_io_status_mpie),
    .io_status_unimp2(csr_io_status_unimp2),
    .io_status_mie(csr_io_status_mie),
    .io_status_unimp1(csr_io_status_unimp1),
    .io_xcpt(csr_io_xcpt),
    .io_cause(csr_io_cause),
    .io_tval(csr_io_tval),
    .io_evec(csr_io_evec),
    .io_illegal(csr_io_illegal),
    .io_retire(csr_io_retire),
    .io_pc(csr_io_pc),
    .io_time(csr_io_time)
  );
  InstDecoder InstDecoder ( // @[BackEnd.scala 91:25:@5064.4]
    .io_inst(InstDecoder_io_inst),
    .io_cinfo_br_type(InstDecoder_io_cinfo_br_type),
    .io_cinfo_op1_sel(InstDecoder_io_cinfo_op1_sel),
    .io_cinfo_op2_sel(InstDecoder_io_cinfo_op2_sel),
    .io_cinfo_rs1_oen(InstDecoder_io_cinfo_rs1_oen),
    .io_cinfo_rs2_oen(InstDecoder_io_cinfo_rs2_oen),
    .io_cinfo_alu_fun(InstDecoder_io_cinfo_alu_fun),
    .io_cinfo_wb_sel(InstDecoder_io_cinfo_wb_sel),
    .io_cinfo_rf_wen(InstDecoder_io_cinfo_rf_wen),
    .io_cinfo_mem_en(InstDecoder_io_cinfo_mem_en),
    .io_cinfo_mem_fcn(InstDecoder_io_cinfo_mem_fcn),
    .io_cinfo_mem_typ(InstDecoder_io_cinfo_mem_typ),
    .io_cinfo_csr_cmd(InstDecoder_io_cinfo_csr_cmd),
    .io_cinfo_illegal(InstDecoder_io_cinfo_illegal),
    .io_cinfo_fencei(InstDecoder_io_cinfo_fencei),
    .io_cinfo_is_branch(InstDecoder_io_cinfo_is_branch),
    .io_cinfo_push(InstDecoder_io_cinfo_push),
    .io_cinfo_pop(InstDecoder_io_cinfo_pop),
    .io_cinfo_rs1_addr(InstDecoder_io_cinfo_rs1_addr),
    .io_cinfo_rs2_addr(InstDecoder_io_cinfo_rs2_addr),
    .io_cinfo_wbaddr(InstDecoder_io_cinfo_wbaddr),
    .io_dinfo_imm_i(InstDecoder_io_dinfo_imm_i),
    .io_dinfo_imm_s(InstDecoder_io_dinfo_imm_s),
    .io_dinfo_imm_sb(InstDecoder_io_dinfo_imm_sb),
    .io_dinfo_imm_u(InstDecoder_io_dinfo_imm_u),
    .io_dinfo_imm_uj(InstDecoder_io_dinfo_imm_uj),
    .io_dinfo_imm_z(InstDecoder_io_dinfo_imm_z)
  );
  Regfile regfile ( // @[BackEnd.scala 122:23:@5095.4]
    .clock(regfile_clock),
    .io_rs1_addr(regfile_io_rs1_addr),
    .io_rs1_data(regfile_io_rs1_data),
    .io_rs2_addr(regfile_io_rs2_addr),
    .io_rs2_data(regfile_io_rs2_data),
    .io_waddr(regfile_io_waddr),
    .io_wdata(regfile_io_wdata),
    .io_wen(regfile_io_wen)
  );
  ALU ALU ( // @[BackEnd.scala 193:19:@5203.4]
    .io_op1(ALU_io_op1),
    .io_op2(ALU_io_op2),
    .io_pc(ALU_io_pc),
    .io_ctrl_fun(ALU_io_ctrl_fun),
    .io_ctrl_br_type(ALU_io_ctrl_br_type),
    .io_ctrl_wb_sel(ALU_io_ctrl_wb_sel),
    .io_ctrl_pc_sel(ALU_io_ctrl_pc_sel),
    .io_rs2_data(ALU_io_rs2_data),
    .io_result(ALU_io_result),
    .io_target_brjmp(ALU_io_target_brjmp),
    .io_target_jpreg(ALU_io_target_jpreg),
    .io_target_conti(ALU_io_target_conti)
  );
  assign dec_wire_rs1_oen = io_front_inst_valid & InstDecoder_io_cinfo_rs1_oen; // @[BackEnd.scala 110:33:@5083.4]
  assign dec_wire_rs2_oen = io_front_inst_valid & InstDecoder_io_cinfo_rs2_oen; // @[BackEnd.scala 111:33:@5085.4]
  assign dec_wire_fencei = io_front_inst_valid & InstDecoder_io_cinfo_fencei; // @[BackEnd.scala 112:33:@5087.4]
  assign exe_wire_fencei = exe_fencei & exe_valid; // @[BackEnd.scala 191:34:@5201.4]
  assign _T_177 = exe_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 131:18:@5104.4]
  assign _T_232 = exe_rf_wen & exe_valid; // @[BackEnd.scala 183:34:@5183.4]
  assign _T_234 = exe_wbaddr != 5'h0; // @[BackEnd.scala 183:61:@5184.4]
  assign exe_wire_rf_wen = _T_232 & _T_234; // @[BackEnd.scala 183:47:@5185.4]
  assign _T_178 = _T_177 & exe_wire_rf_wen; // @[BackEnd.scala 131:42:@5105.4]
  assign _T_179 = mem_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 132:18:@5106.4]
  assign _T_329 = mem_rf_wen & mem_valid; // @[BackEnd.scala 267:35:@5329.4]
  assign _T_331 = mem_wbaddr != 5'h0; // @[BackEnd.scala 267:62:@5330.4]
  assign mem_wire_rf_wen = _T_329 & _T_331; // @[BackEnd.scala 267:48:@5331.4]
  assign _T_180 = _T_179 & mem_wire_rf_wen; // @[BackEnd.scala 132:42:@5107.4]
  assign _T_181 = wb_wbaddr == InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 133:18:@5108.4]
  assign _T_366 = wb_rf_wen & wb_valid; // @[BackEnd.scala 315:33:@5473.4]
  assign _T_368 = wb_wbaddr != 5'h0; // @[BackEnd.scala 315:58:@5474.4]
  assign wb_wire_rf_wen = _T_366 & _T_368; // @[BackEnd.scala 315:45:@5475.4]
  assign _T_182 = _T_181 & wb_wire_rf_wen; // @[BackEnd.scala 133:42:@5109.4]
  assign rf_rs1_data = regfile_io_rs1_data; // @[BackEnd.scala 123:25:@5098.4 BackEnd.scala 127:15:@5102.4]
  assign _T_183 = _T_182 ? wb_wbdata : rf_rs1_data; // @[Mux.scala 61:16:@5110.4]
  assign _T_360 = mem_wb_sel == 2'h1; // @[BackEnd.scala 302:17:@5458.4]
  assign _T_361 = mem_wb_sel == 2'h3; // @[BackEnd.scala 303:17:@5459.4]
  assign _T_362 = _T_361 ? csr_io_rw_rdata : mem_exe_out; // @[Mux.scala 61:16:@5460.4]
  assign mem_wbdata = _T_360 ? io_mem_resp_bits_data : _T_362; // @[Mux.scala 61:16:@5461.4]
  assign _T_184 = _T_180 ? mem_wbdata : _T_183; // @[Mux.scala 61:16:@5111.4]
  assign exe_wbdata = ALU_io_result; // @[BackEnd.scala 104:24:@5078.4 BackEnd.scala 201:20:@5213.4]
  assign dec_rs1_data = _T_178 ? exe_wbdata : _T_184; // @[Mux.scala 61:16:@5112.4]
  assign _T_186 = exe_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 137:18:@5114.4]
  assign _T_187 = _T_186 & exe_wire_rf_wen; // @[BackEnd.scala 137:42:@5115.4]
  assign _T_188 = mem_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 138:18:@5116.4]
  assign _T_189 = _T_188 & mem_wire_rf_wen; // @[BackEnd.scala 138:42:@5117.4]
  assign _T_190 = wb_wbaddr == InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 139:18:@5118.4]
  assign _T_191 = _T_190 & wb_wire_rf_wen; // @[BackEnd.scala 139:42:@5119.4]
  assign rf_rs2_data = regfile_io_rs2_data; // @[BackEnd.scala 124:25:@5099.4 BackEnd.scala 128:15:@5103.4]
  assign _T_192 = _T_191 ? wb_wbdata : rf_rs2_data; // @[Mux.scala 61:16:@5120.4]
  assign _T_193 = _T_189 ? mem_wbdata : _T_192; // @[Mux.scala 61:16:@5121.4]
  assign dec_rs2_data = _T_187 ? exe_wbdata : _T_193; // @[Mux.scala 61:16:@5122.4]
  assign _T_195 = InstDecoder_io_cinfo_op1_sel == 2'h2; // @[BackEnd.scala 143:24:@5124.4]
  assign _T_196 = InstDecoder_io_cinfo_op1_sel == 2'h1; // @[BackEnd.scala 144:24:@5125.4]
  assign _T_197 = _T_196 ? io_front_pc : dec_rs1_data; // @[Mux.scala 61:16:@5126.4]
  assign dec_op1_data = _T_195 ? InstDecoder_io_dinfo_imm_z : _T_197; // @[Mux.scala 61:16:@5127.4]
  assign _T_199 = InstDecoder_io_cinfo_op2_sel == 3'h1; // @[BackEnd.scala 147:24:@5129.4]
  assign _T_200 = InstDecoder_io_cinfo_op2_sel == 3'h2; // @[BackEnd.scala 148:24:@5130.4]
  assign _T_201 = InstDecoder_io_cinfo_op2_sel == 3'h3; // @[BackEnd.scala 149:24:@5131.4]
  assign _T_202 = InstDecoder_io_cinfo_op2_sel == 3'h4; // @[BackEnd.scala 150:24:@5132.4]
  assign _T_203 = InstDecoder_io_cinfo_op2_sel == 3'h5; // @[BackEnd.scala 151:24:@5133.4]
  assign _T_204 = _T_203 ? InstDecoder_io_dinfo_imm_uj : dec_rs2_data; // @[Mux.scala 61:16:@5134.4]
  assign _T_205 = _T_202 ? InstDecoder_io_dinfo_imm_u : _T_204; // @[Mux.scala 61:16:@5135.4]
  assign _T_206 = _T_201 ? InstDecoder_io_dinfo_imm_sb : _T_205; // @[Mux.scala 61:16:@5136.4]
  assign _T_207 = _T_200 ? InstDecoder_io_dinfo_imm_s : _T_206; // @[Mux.scala 61:16:@5137.4]
  assign dec_op2_data = _T_199 ? InstDecoder_io_dinfo_imm_i : _T_207; // @[Mux.scala 61:16:@5138.4]
  assign exe_wire_mem_en = exe_mem_en & exe_valid; // @[BackEnd.scala 184:34:@5187.4]
  assign _T_430 = exe_mem_fcn == 1'h0; // @[BackEnd.scala 325:60:@5541.4]
  assign exe_load_inst = exe_wire_mem_en & _T_430; // @[BackEnd.scala 325:45:@5542.4]
  assign _T_432 = exe_load_inst & _T_177; // @[BackEnd.scala 328:20:@5544.4]
  assign _T_434 = InstDecoder_io_cinfo_rs1_addr != 5'h0; // @[BackEnd.scala 328:79:@5545.4]
  assign _T_435 = _T_432 & _T_434; // @[BackEnd.scala 328:57:@5546.4]
  assign _T_436 = _T_435 & dec_wire_rs1_oen; // @[BackEnd.scala 328:87:@5547.4]
  assign _T_438 = exe_load_inst & _T_186; // @[BackEnd.scala 329:20:@5549.4]
  assign _T_440 = InstDecoder_io_cinfo_rs2_addr != 5'h0; // @[BackEnd.scala 329:79:@5550.4]
  assign _T_441 = _T_438 & _T_440; // @[BackEnd.scala 329:57:@5551.4]
  assign _T_442 = _T_441 & dec_wire_rs2_oen; // @[BackEnd.scala 329:87:@5552.4]
  assign _T_443 = _T_436 | _T_442; // @[BackEnd.scala 328:108:@5553.4]
  assign exe_wire_csr_cmd = exe_valid ? exe_csr_cmd : 3'h0; // @[BackEnd.scala 185:26:@5189.4]
  assign _T_444 = exe_wire_csr_cmd != 3'h0; // @[BackEnd.scala 330:22:@5554.4]
  assign stall_0 = _T_443 | _T_444; // @[BackEnd.scala 329:108:@5555.4]
  assign mem_wire_mem_en = mem_mem_en & mem_valid; // @[BackEnd.scala 268:35:@5333.4]
  assign _T_450 = io_mem_resp_valid == 1'h0; // @[BackEnd.scala 333:42:@5560.4]
  assign _T_451 = mem_wire_mem_en & _T_450; // @[BackEnd.scala 333:39:@5561.4]
  assign mem_wire_ma_load = mem_ma_load & mem_valid; // @[BackEnd.scala 271:36:@5339.4]
  assign mem_wire_ma_store = mem_ma_store & mem_valid; // @[BackEnd.scala 272:37:@5341.4]
  assign mem_wire_ma_valid = mem_wire_ma_load | mem_wire_ma_store; // @[BackEnd.scala 273:41:@5343.4]
  assign _T_453 = mem_wire_ma_valid == 1'h0; // @[BackEnd.scala 333:64:@5562.4]
  assign stall_2 = _T_451 & _T_453; // @[BackEnd.scala 333:61:@5563.4]
  assign _T_213 = stall_2 == 1'h0; // @[BackEnd.scala 153:51:@5142.4]
  assign _T_214 = stall_0 & _T_213; // @[BackEnd.scala 153:48:@5143.4]
  assign _T_215 = _T_214 | io_front_xcpt_valid; // @[BackEnd.scala 153:70:@5144.4]
  assign _T_223 = io_front_kill == 1'h0; // @[BackEnd.scala 157:34:@5153.8]
  assign _T_224 = io_front_inst_valid & _T_223; // @[BackEnd.scala 157:31:@5154.8]
  assign _T_225 = InstDecoder_io_cinfo_csr_cmd == 3'h2; // @[BackEnd.scala 161:44:@5158.8]
  assign _T_226 = InstDecoder_io_cinfo_csr_cmd == 3'h3; // @[BackEnd.scala 161:75:@5159.8]
  assign _T_227 = _T_225 | _T_226; // @[BackEnd.scala 161:54:@5160.8]
  assign _T_229 = InstDecoder_io_cinfo_rs1_addr == 5'h0; // @[BackEnd.scala 162:26:@5161.8]
  assign _T_230 = _T_227 & _T_229; // @[BackEnd.scala 161:86:@5162.8]
  assign _T_231 = _T_230 ? 3'h5 : InstDecoder_io_cinfo_csr_cmd; // @[BackEnd.scala 161:24:@5163.8]
  assign _GEN_0 = _T_213 ? _T_224 : exe_valid; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_1 = _T_213 ? InstDecoder_io_cinfo_rf_wen : exe_rf_wen; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_2 = _T_213 ? InstDecoder_io_cinfo_mem_en : exe_mem_en; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_3 = _T_213 ? _T_231 : exe_csr_cmd; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_4 = _T_213 ? InstDecoder_io_cinfo_illegal : exe_illegal; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_5 = _T_213 ? InstDecoder_io_cinfo_fencei : exe_fencei; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_6 = _T_213 ? InstDecoder_io_cinfo_br_type : exe_br_type; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_7 = _T_213 ? io_front_pc : exe_pc; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_8 = _T_213 ? dec_op1_data : exe_op1_data; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_9 = _T_213 ? dec_op2_data : exe_op2_data; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_10 = _T_213 ? dec_rs2_data : exe_rs2_data; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_11 = _T_213 ? InstDecoder_io_inst : exe_inst; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_12 = _T_213 ? InstDecoder_io_cinfo_alu_fun : exe_alu_fun; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_13 = _T_213 ? InstDecoder_io_cinfo_wb_sel : exe_wb_sel; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_14 = _T_213 ? InstDecoder_io_cinfo_wbaddr : exe_wbaddr; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_15 = _T_213 ? InstDecoder_io_cinfo_mem_fcn : exe_mem_fcn; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_16 = _T_213 ? InstDecoder_io_cinfo_mem_typ : exe_mem_typ; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_17 = _T_213 ? InstDecoder_io_cinfo_is_branch : exe_branch; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_18 = _T_213 ? InstDecoder_io_cinfo_push : exe_push; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_19 = _T_213 ? InstDecoder_io_cinfo_pop : exe_pop; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_20 = _T_213 ? io_front_pred : exe_pred; // @[BackEnd.scala 156:54:@5152.6]
  assign _GEN_21 = _T_215 ? 1'h0 : _GEN_0; // @[BackEnd.scala 153:94:@5145.4]
  assign exe_wire_br_type = exe_valid ? exe_br_type : 4'h0; // @[BackEnd.scala 186:26:@5191.4]
  assign exe_wire_branch = exe_valid & exe_branch; // @[BackEnd.scala 187:33:@5193.4]
  assign exe_wire_push = exe_valid & exe_push; // @[BackEnd.scala 188:33:@5195.4]
  assign exe_wire_pop = exe_valid & exe_pop; // @[BackEnd.scala 189:33:@5197.4]
  assign _GEN_42 = exe_wire_pop ? 1'h0 : _T_248; // @[BackEnd.scala 74:20:@5220.6]
  assign _GEN_43 = _T_213 ? 1'h1 : _GEN_42; // @[BackEnd.scala 73:20:@5216.4]
  assign _GEN_44 = exe_wire_push ? 1'h0 : _T_256; // @[BackEnd.scala 74:20:@5231.6]
  assign _GEN_45 = _T_213 ? 1'h1 : _GEN_44; // @[BackEnd.scala 73:20:@5227.4]
  assign _T_260 = ALU_io_ctrl_pc_sel == 2'h1; // @[BackEnd.scala 208:25:@5237.4]
  assign _T_261 = ALU_io_ctrl_pc_sel == 2'h2; // @[BackEnd.scala 209:25:@5238.4]
  assign _T_262 = _T_261 ? ALU_io_target_jpreg : ALU_io_target_conti; // @[BackEnd.scala 209:8:@5239.4]
  assign next_pc = _T_260 ? ALU_io_target_brjmp : _T_262; // @[BackEnd.scala 208:8:@5240.4]
  assign _T_266 = exe_wire_pop ? 2'h1 : 2'h3; // @[BackEnd.scala 215:10:@5242.4]
  assign _T_268 = exe_wire_br_type != 4'h0; // @[BackEnd.scala 217:53:@5245.4]
  assign _GEN_46 = _T_268 ? 1'h0 : _T_273; // @[BackEnd.scala 74:20:@5252.6]
  assign _GEN_47 = _T_213 ? 1'h1 : _GEN_46; // @[BackEnd.scala 73:20:@5248.4]
  assign _T_281 = next_pc != exe_pred; // @[BackEnd.scala 221:42:@5263.4]
  assign mispredict = _T_281 & exe_valid; // @[BackEnd.scala 221:55:@5264.4]
  assign _T_283 = exe_mem_typ[1:0]; // @[BackEnd.scala 224:45:@5266.4]
  assign _T_286 = ALU_io_result[0]; // @[BackEnd.scala 225:22:@5267.4]
  assign _T_288 = ALU_io_result[1:0]; // @[BackEnd.scala 226:22:@5268.4]
  assign _T_290 = _T_288 != 2'h0; // @[BackEnd.scala 226:28:@5269.4]
  assign _T_291 = 2'h3 == _T_283; // @[Mux.scala 46:19:@5270.4]
  assign _T_292 = _T_291 ? _T_290 : 1'h0; // @[Mux.scala 46:16:@5271.4]
  assign _T_293 = 2'h2 == _T_283; // @[Mux.scala 46:19:@5272.4]
  assign exe_wire_ma_valid = _T_293 ? _T_286 : _T_292; // @[Mux.scala 46:16:@5273.4]
  assign exe_wire_ma_load = _T_430 & exe_wire_ma_valid; // @[BackEnd.scala 228:46:@5276.4]
  assign exe_wire_ma_store = exe_mem_fcn & exe_wire_ma_valid; // @[BackEnd.scala 229:46:@5279.4]
  assign _T_300 = exe_wire_ma_valid == 1'h0; // @[BackEnd.scala 232:46:@5281.4]
  assign _T_301 = exe_wire_mem_en & _T_300; // @[BackEnd.scala 232:43:@5282.4]
  assign _T_303 = io_front_xcpt_valid == 1'h0; // @[BackEnd.scala 232:68:@5283.4]
  assign _T_312 = stall_2 | io_front_xcpt_valid; // @[BackEnd.scala 243:47:@5296.4]
  assign _T_320 = _T_260 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@5320.8]
  assign _T_321 = _T_320 & ALU_io_target_brjmp; // @[BackEnd.scala 262:70:@5321.8]
  assign _T_326 = _T_261 ? 32'hffffffff : 32'h0; // @[Bitwise.scala 72:12:@5324.8]
  assign _T_327 = _T_326 & ALU_io_target_jpreg; // @[BackEnd.scala 263:74:@5325.8]
  assign _T_328 = _T_321 | _T_327; // @[BackEnd.scala 262:90:@5326.8]
  assign _GEN_48 = _T_213 ? exe_valid : mem_valid; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_49 = _T_213 ? exe_rf_wen : mem_rf_wen; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_50 = _T_213 ? exe_mem_en : mem_mem_en; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_51 = _T_213 ? exe_csr_cmd : mem_csr_cmd; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_52 = _T_213 ? exe_illegal : mem_illegal; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_53 = _T_213 ? exe_pc : mem_pc; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_54 = _T_213 ? exe_inst : mem_inst; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_55 = _T_213 ? exe_wb_sel : mem_wb_sel; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_56 = _T_213 ? exe_wbaddr : mem_wbaddr; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_60 = _T_213 ? exe_wire_ma_load : mem_ma_load; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_61 = _T_213 ? exe_wire_ma_store : mem_ma_store; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_62 = _T_213 ? exe_wbdata : mem_exe_out; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_63 = _T_213 ? _T_328 : mem_jpnpc; // @[BackEnd.scala 245:34:@5302.6]
  assign _GEN_64 = _T_312 ? 1'h0 : _GEN_48; // @[BackEnd.scala 243:71:@5297.4]
  assign mem_wire_illegal = mem_illegal & mem_valid; // @[BackEnd.scala 270:36:@5337.4]
  assign _T_340 = mem_jpnpc[1:0]; // @[BackEnd.scala 281:32:@5439.4]
  assign _T_342 = _T_340 != 2'h0; // @[BackEnd.scala 281:38:@5440.4]
  assign ma_jump = _T_342 & mem_valid; // @[BackEnd.scala 281:42:@5441.4]
  assign _T_344 = mem_wire_ma_valid | ma_jump; // @[BackEnd.scala 283:57:@5443.4]
  assign _T_351 = mem_wire_illegal ? 2'h2 : 2'h0; // @[Mux.scala 61:16:@5446.4]
  assign _T_352 = mem_wire_ma_store ? 3'h6 : {{1'd0}, _T_351}; // @[Mux.scala 61:16:@5447.4]
  assign _T_353 = mem_wire_ma_load ? 3'h4 : _T_352; // @[Mux.scala 61:16:@5448.4]
  assign _T_354 = ma_jump ? 3'h0 : _T_353; // @[Mux.scala 61:16:@5449.4]
  assign _T_356 = mem_wire_illegal ? mem_inst : 32'h0; // @[Mux.scala 61:16:@5451.4]
  assign _T_357 = mem_wire_ma_valid ? mem_exe_out : _T_356; // @[Mux.scala 61:16:@5452.4]
  assign _GEN_80 = _T_312 ? 1'h0 : mem_valid; // @[BackEnd.scala 305:50:@5464.4]
  assign _GEN_84 = mispredict ? 1'h0 : _T_459; // @[BackEnd.scala 74:20:@5571.6]
  assign _GEN_85 = _T_213 ? 1'h1 : _GEN_84; // @[BackEnd.scala 73:20:@5567.4]
  assign _T_464 = {stall_2,1'h0,stall_0}; // @[BackEnd.scala 336:32:@5577.4]
  assign _T_466 = _T_464 != 3'h0; // @[BackEnd.scala 336:39:@5578.4]
  assign _T_472 = stall_0 ? 8'h53 : 8'h20; // @[BackEnd.scala 345:10:@5581.4]
  assign _T_473 = stall_2 ? 8'h46 : _T_472; // @[BackEnd.scala 344:10:@5582.4]
  assign _T_481 = ALU_io_ctrl_pc_sel == 2'h3; // @[BackEnd.scala 348:27:@5585.4]
  assign _T_484 = ALU_io_ctrl_pc_sel == 2'h0; // @[BackEnd.scala 349:27:@5586.4]
  assign _T_487 = _T_484 ? 8'h20 : 8'h3f; // @[BackEnd.scala 349:10:@5587.4]
  assign _T_488 = _T_481 ? 8'h45 : _T_487; // @[BackEnd.scala 348:10:@5588.4]
  assign _T_489 = _T_261 ? 8'h4a : _T_488; // @[BackEnd.scala 347:10:@5589.4]
  assign _T_490 = _T_260 ? 8'h42 : _T_489; // @[BackEnd.scala 346:10:@5590.4]
  assign _T_493 = csr_io_illegal ? 8'h58 : 8'h20; // @[BackEnd.scala 350:10:@5591.4]
  assign _T_495 = exe_valid == 1'h0; // @[BackEnd.scala 351:34:@5592.4]
  assign _T_496 = io_front_xcpt_valid | _T_495; // @[BackEnd.scala 351:31:@5593.4]
  assign _T_497 = _T_496 ? 32'h4033 : exe_inst; // @[BackEnd.scala 351:10:@5594.4]
  assign _T_500 = reset == 1'h0; // @[BackEnd.scala 339:9:@5596.4]
  assign _T_504 = ALU_io_target_conti != exe_pred; // @[BackEnd.scala 368:24:@5608.6]
  assign io_mem_req_valid = _T_301 & _T_303; // @[BackEnd.scala 232:24:@5285.4]
  assign io_mem_req_bits_addr = ALU_io_result; // @[BackEnd.scala 233:24:@5286.4]
  assign io_mem_req_bits_data = exe_rs2_data; // @[BackEnd.scala 236:24:@5289.4]
  assign io_mem_req_bits_fcn = exe_mem_fcn; // @[BackEnd.scala 234:24:@5287.4]
  assign io_mem_req_bits_typ = exe_mem_typ; // @[BackEnd.scala 235:24:@5288.4]
  assign io_cyc = csr_io_time; // @[BackEnd.scala 87:10:@5062.4]
  assign io_front_xcpt_valid = csr_io_xcpt | csr_io_eret; // @[BackEnd.scala 295:23:@5456.4]
  assign io_front_xcpt_bits = csr_io_evec; // @[BackEnd.scala 296:23:@5457.4]
  assign io_front_kill = mispredict & _T_459; // @[BackEnd.scala 335:17:@5575.4]
  assign io_front_fence = dec_wire_fencei | exe_wire_fencei; // @[BackEnd.scala 113:20:@5090.4]
  assign io_front_forward = _T_466 == 1'h0; // @[BackEnd.scala 336:21:@5580.4]
  assign io_front_ras_pop = exe_wire_pop & _T_248; // @[BackEnd.scala 203:27:@5224.4]
  assign io_front_ras_push_valid = exe_wire_push & _T_256; // @[BackEnd.scala 204:27:@5235.4]
  assign io_front_ras_push_bits = ALU_io_target_conti; // @[BackEnd.scala 205:27:@5236.4]
  assign io_front_fb_pc = exe_pc; // @[BackEnd.scala 212:18:@5241.4]
  assign io_front_fb_type = exe_wire_branch ? 2'h2 : _T_266; // @[BackEnd.scala 213:20:@5244.4]
  assign io_front_feedBack_valid = _T_268 & _T_273; // @[BackEnd.scala 217:27:@5256.4]
  assign io_front_feedBack_bits_redirect = _T_260 | _T_261; // @[BackEnd.scala 219:35:@5261.4]
  assign io_front_feedBack_bits_tgt = _T_260 ? ALU_io_target_brjmp : _T_262; // @[BackEnd.scala 218:30:@5257.4]
  assign csr_clock = clock; // @[:@5059.4]
  assign csr_reset = reset; // @[:@5060.4]
  assign csr_io_rw_cmd = mem_valid ? mem_csr_cmd : 3'h0; // @[BackEnd.scala 278:19:@5437.4]
  assign csr_io_rw_addr = mem_inst[31:20]; // @[BackEnd.scala 276:19:@5435.4]
  assign csr_io_rw_wdata = mem_exe_out; // @[BackEnd.scala 277:19:@5436.4]
  assign csr_io_xcpt = _T_344 | mem_wire_illegal; // @[BackEnd.scala 283:16:@5445.4]
  assign csr_io_cause = {{29'd0}, _T_354}; // @[BackEnd.scala 284:16:@5450.4]
  assign csr_io_tval = ma_jump ? mem_jpnpc : _T_357; // @[BackEnd.scala 290:16:@5454.4]
  assign csr_io_illegal = 1'h0;
  assign csr_io_retire = {{1'd0}, wb_valid}; // @[BackEnd.scala 320:20:@5480.4]
  assign csr_io_pc = mem_pc; // @[BackEnd.scala 279:19:@5438.4]
  assign InstDecoder_io_inst = io_front_inst_bits; // @[BackEnd.scala 108:20:@5081.4]
  assign regfile_clock = clock; // @[:@5096.4]
  assign regfile_io_rs1_addr = InstDecoder_io_cinfo_rs1_addr; // @[BackEnd.scala 125:23:@5100.4]
  assign regfile_io_rs2_addr = InstDecoder_io_cinfo_rs2_addr; // @[BackEnd.scala 126:23:@5101.4]
  assign regfile_io_waddr = wb_wbaddr; // @[BackEnd.scala 316:20:@5477.4]
  assign regfile_io_wdata = wb_wbdata; // @[BackEnd.scala 317:20:@5478.4]
  assign regfile_io_wen = _T_366 & _T_368; // @[BackEnd.scala 318:20:@5479.4]
  assign ALU_io_op1 = exe_op1_data; // @[BackEnd.scala 194:20:@5206.4]
  assign ALU_io_op2 = exe_op2_data; // @[BackEnd.scala 195:20:@5207.4]
  assign ALU_io_pc = exe_pc; // @[BackEnd.scala 197:20:@5209.4]
  assign ALU_io_ctrl_fun = exe_alu_fun; // @[BackEnd.scala 198:20:@5210.4]
  assign ALU_io_ctrl_br_type = exe_valid ? exe_br_type : 4'h0; // @[BackEnd.scala 199:20:@5211.4]
  assign ALU_io_ctrl_wb_sel = exe_wb_sel; // @[BackEnd.scala 200:20:@5212.4]
  assign ALU_io_rs2_data = exe_rs2_data; // @[BackEnd.scala 196:20:@5208.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifndef RANDOM
`define RANDOM $random
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifdef INIT_RANDOM
      `INIT_RANDOM
    `endif
    `ifndef VERILATOR
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{`RANDOM}};
  exe_rf_wen = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{`RANDOM}};
  exe_wbaddr = _RAND_1[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{`RANDOM}};
  exe_mem_en = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{`RANDOM}};
  exe_csr_cmd = _RAND_3[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{`RANDOM}};
  exe_illegal = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{`RANDOM}};
  exe_pc = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{`RANDOM}};
  exe_inst = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{`RANDOM}};
  exe_rs2_data = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{`RANDOM}};
  exe_wb_sel = _RAND_8[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{`RANDOM}};
  exe_mem_fcn = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{`RANDOM}};
  exe_mem_typ = _RAND_10[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{`RANDOM}};
  exe_fencei = _RAND_11[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{`RANDOM}};
  exe_br_type = _RAND_12[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{`RANDOM}};
  exe_branch = _RAND_13[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{`RANDOM}};
  exe_push = _RAND_14[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{`RANDOM}};
  exe_pop = _RAND_15[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{`RANDOM}};
  exe_pred = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{`RANDOM}};
  exe_op1_data = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{`RANDOM}};
  exe_op2_data = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{`RANDOM}};
  exe_alu_fun = _RAND_19[3:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{`RANDOM}};
  exe_valid = _RAND_20[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{`RANDOM}};
  mem_rf_wen = _RAND_21[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{`RANDOM}};
  mem_wbaddr = _RAND_22[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{`RANDOM}};
  mem_mem_en = _RAND_23[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{`RANDOM}};
  mem_csr_cmd = _RAND_24[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{`RANDOM}};
  mem_illegal = _RAND_25[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{`RANDOM}};
  mem_pc = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{`RANDOM}};
  mem_inst = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{`RANDOM}};
  mem_wb_sel = _RAND_28[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{`RANDOM}};
  mem_valid = _RAND_29[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{`RANDOM}};
  wb_rf_wen = _RAND_30[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{`RANDOM}};
  wb_wbaddr = _RAND_31[4:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{`RANDOM}};
  wb_valid = _RAND_32[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{`RANDOM}};
  wb_wbdata = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{`RANDOM}};
  mem_exe_out = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{`RANDOM}};
  mem_ma_load = _RAND_35[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{`RANDOM}};
  mem_ma_store = _RAND_36[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{`RANDOM}};
  _T_248 = _RAND_37[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{`RANDOM}};
  _T_256 = _RAND_38[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{`RANDOM}};
  _T_273 = _RAND_39[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{`RANDOM}};
  mem_jpnpc = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{`RANDOM}};
  _T_459 = _RAND_41[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_rf_wen <= InstDecoder_io_cinfo_rf_wen;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_wbaddr <= InstDecoder_io_cinfo_wbaddr;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_mem_en <= InstDecoder_io_cinfo_mem_en;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        if (_T_230) begin
          exe_csr_cmd <= 3'h5;
        end else begin
          exe_csr_cmd <= InstDecoder_io_cinfo_csr_cmd;
        end
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_illegal <= InstDecoder_io_cinfo_illegal;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_pc <= io_front_pc;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_inst <= InstDecoder_io_inst;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        if (_T_187) begin
          exe_rs2_data <= exe_wbdata;
        end else begin
          if (_T_189) begin
            if (_T_360) begin
              exe_rs2_data <= io_mem_resp_bits_data;
            end else begin
              if (_T_361) begin
                exe_rs2_data <= csr_io_rw_rdata;
              end else begin
                exe_rs2_data <= mem_exe_out;
              end
            end
          end else begin
            if (_T_191) begin
              exe_rs2_data <= wb_wbdata;
            end else begin
              exe_rs2_data <= rf_rs2_data;
            end
          end
        end
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_wb_sel <= InstDecoder_io_cinfo_wb_sel;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_mem_fcn <= InstDecoder_io_cinfo_mem_fcn;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_mem_typ <= InstDecoder_io_cinfo_mem_typ;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_fencei <= InstDecoder_io_cinfo_fencei;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_br_type <= InstDecoder_io_cinfo_br_type;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_branch <= InstDecoder_io_cinfo_is_branch;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_push <= InstDecoder_io_cinfo_push;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_pop <= InstDecoder_io_cinfo_pop;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_pred <= io_front_pred;
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        if (_T_195) begin
          exe_op1_data <= InstDecoder_io_dinfo_imm_z;
        end else begin
          if (_T_196) begin
            exe_op1_data <= io_front_pc;
          end else begin
            if (_T_178) begin
              exe_op1_data <= exe_wbdata;
            end else begin
              if (_T_180) begin
                if (_T_360) begin
                  exe_op1_data <= io_mem_resp_bits_data;
                end else begin
                  if (_T_361) begin
                    exe_op1_data <= csr_io_rw_rdata;
                  end else begin
                    exe_op1_data <= mem_exe_out;
                  end
                end
              end else begin
                if (_T_182) begin
                  exe_op1_data <= wb_wbdata;
                end else begin
                  exe_op1_data <= rf_rs1_data;
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        if (_T_199) begin
          exe_op2_data <= InstDecoder_io_dinfo_imm_i;
        end else begin
          if (_T_200) begin
            exe_op2_data <= InstDecoder_io_dinfo_imm_s;
          end else begin
            if (_T_201) begin
              exe_op2_data <= InstDecoder_io_dinfo_imm_sb;
            end else begin
              if (_T_202) begin
                exe_op2_data <= InstDecoder_io_dinfo_imm_u;
              end else begin
                if (_T_203) begin
                  exe_op2_data <= InstDecoder_io_dinfo_imm_uj;
                end else begin
                  if (_T_187) begin
                    exe_op2_data <= exe_wbdata;
                  end else begin
                    if (_T_189) begin
                      if (_T_360) begin
                        exe_op2_data <= io_mem_resp_bits_data;
                      end else begin
                        if (_T_361) begin
                          exe_op2_data <= csr_io_rw_rdata;
                        end else begin
                          exe_op2_data <= mem_exe_out;
                        end
                      end
                    end else begin
                      if (_T_191) begin
                        exe_op2_data <= wb_wbdata;
                      end else begin
                        exe_op2_data <= rf_rs2_data;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (!(_T_215)) begin
      if (_T_213) begin
        exe_alu_fun <= InstDecoder_io_cinfo_alu_fun;
      end
    end
    if (reset) begin
      exe_valid <= 1'h0;
    end else begin
      if (_T_215) begin
        exe_valid <= 1'h0;
      end else begin
        if (_T_213) begin
          exe_valid <= _T_224;
        end
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_rf_wen <= exe_rf_wen;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_wbaddr <= exe_wbaddr;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_mem_en <= exe_mem_en;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_csr_cmd <= exe_csr_cmd;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_illegal <= exe_illegal;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_pc <= exe_pc;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_inst <= exe_inst;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_wb_sel <= exe_wb_sel;
      end
    end
    if (reset) begin
      mem_valid <= 1'h0;
    end else begin
      if (_T_312) begin
        mem_valid <= 1'h0;
      end else begin
        if (_T_213) begin
          mem_valid <= exe_valid;
        end
      end
    end
    if (!(_T_312)) begin
      wb_rf_wen <= mem_rf_wen;
    end
    if (!(_T_312)) begin
      wb_wbaddr <= mem_wbaddr;
    end
    if (reset) begin
      wb_valid <= 1'h0;
    end else begin
      if (_T_312) begin
        wb_valid <= 1'h0;
      end else begin
        wb_valid <= mem_valid;
      end
    end
    if (!(_T_312)) begin
      if (_T_360) begin
        wb_wbdata <= io_mem_resp_bits_data;
      end else begin
        if (_T_361) begin
          wb_wbdata <= csr_io_rw_rdata;
        end else begin
          wb_wbdata <= mem_exe_out;
        end
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_exe_out <= exe_wbdata;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_ma_load <= exe_wire_ma_load;
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_ma_store <= exe_wire_ma_store;
      end
    end
    if (reset) begin
      _T_248 <= 1'h1;
    end else begin
      if (_T_213) begin
        _T_248 <= 1'h1;
      end else begin
        if (exe_wire_pop) begin
          _T_248 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_256 <= 1'h1;
    end else begin
      if (_T_213) begin
        _T_256 <= 1'h1;
      end else begin
        if (exe_wire_push) begin
          _T_256 <= 1'h0;
        end
      end
    end
    if (reset) begin
      _T_273 <= 1'h1;
    end else begin
      if (_T_213) begin
        _T_273 <= 1'h1;
      end else begin
        if (_T_268) begin
          _T_273 <= 1'h0;
        end
      end
    end
    if (!(_T_312)) begin
      if (_T_213) begin
        mem_jpnpc <= _T_328;
      end
    end
    if (reset) begin
      _T_459 <= 1'h1;
    end else begin
      if (_T_213) begin
        _T_459 <= 1'h1;
      end else begin
        if (mispredict) begin
          _T_459 <= 1'h0;
        end
      end
    end
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (_T_500) begin
          $fwrite(32'h80000002,"Core: Cyc= %d (%x, %x, %x) %c %c %c ExeInst: DASM(%x)\n",io_cyc,io_front_pc,exe_pc,mem_pc,_T_473,_T_490,_T_493,_T_497); // @[BackEnd.scala 339:9:@5598.6]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (wb_valid & _T_500) begin
          $fwrite(32'h80000002,"Core: Cyc= %d WB[ %x %x %x]\n",io_cyc,wb_wire_rf_wen,wb_wbaddr,wb_wbdata); // @[BackEnd.scala 354:11:@5604.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
    `ifndef SYNTHESIS
    `ifdef PRINTF_COND
      if (`PRINTF_COND) begin
    `endif
        if (io_front_feedBack_valid & _T_500) begin
          $fwrite(32'h80000002,"BranchJump: Cyc= %d kill %x pc %x tgt %x actual %x expect %x inst DASM(%x)\n",io_cyc,mispredict,exe_pc,next_pc,io_front_feedBack_bits_redirect,_T_504,exe_inst); // @[BackEnd.scala 362:11:@5612.8]
        end
    `ifdef PRINTF_COND
      end
    `endif
    `endif // SYNTHESIS
  end
endmodule
module rv32_toy( // @[:@5616.2]
  input         clock, // @[:@5617.4]
  input         reset, // @[:@5618.4]
  output        io_imem_req_valid, // @[:@5619.4]
  output [31:0] io_imem_req_bits_addr, // @[:@5619.4]
  input         io_imem_resp_valid, // @[:@5619.4]
  input  [31:0] io_imem_resp_bits_data, // @[:@5619.4]
  output        io_dmem_req_valid, // @[:@5619.4]
  output [31:0] io_dmem_req_bits_addr, // @[:@5619.4]
  output [31:0] io_dmem_req_bits_data, // @[:@5619.4]
  output        io_dmem_req_bits_fcn, // @[:@5619.4]
  output [2:0]  io_dmem_req_bits_typ, // @[:@5619.4]
  input         io_dmem_resp_valid, // @[:@5619.4]
  input  [31:0] io_dmem_resp_bits_data // @[:@5619.4]
);
  wire  frontEnd_clock; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_reset; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_cyc; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_mem_req_valid; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_mem_req_bits_addr; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_mem_resp_valid; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_mem_resp_bits_data; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_xcpt_valid; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_xcpt_bits; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_kill; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_fence; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_forward; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_ras_pop; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_ras_push_valid; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_ras_push_bits; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_fb_pc; // @[Core.scala 30:24:@5621.4]
  wire [1:0] frontEnd_io_back_fb_type; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_feedBack_valid; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_feedBack_bits_redirect; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_feedBack_bits_tgt; // @[Core.scala 30:24:@5621.4]
  wire  frontEnd_io_back_inst_valid; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_inst_bits; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_pc; // @[Core.scala 30:24:@5621.4]
  wire [31:0] frontEnd_io_back_pred; // @[Core.scala 30:24:@5621.4]
  wire  backEnd_clock; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_reset; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_mem_req_valid; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_mem_req_bits_addr; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_mem_req_bits_data; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_mem_req_bits_fcn; // @[Core.scala 31:24:@5624.4]
  wire [2:0] backEnd_io_mem_req_bits_typ; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_mem_resp_valid; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_mem_resp_bits_data; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_cyc; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_xcpt_valid; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_xcpt_bits; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_kill; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_fence; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_forward; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_ras_pop; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_ras_push_valid; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_ras_push_bits; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_fb_pc; // @[Core.scala 31:24:@5624.4]
  wire [1:0] backEnd_io_front_fb_type; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_feedBack_valid; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_feedBack_bits_redirect; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_feedBack_bits_tgt; // @[Core.scala 31:24:@5624.4]
  wire  backEnd_io_front_inst_valid; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_inst_bits; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_pc; // @[Core.scala 31:24:@5624.4]
  wire [31:0] backEnd_io_front_pred; // @[Core.scala 31:24:@5624.4]
  FrontEnd frontEnd ( // @[Core.scala 30:24:@5621.4]
    .clock(frontEnd_clock),
    .reset(frontEnd_reset),
    .io_cyc(frontEnd_io_cyc),
    .io_mem_req_valid(frontEnd_io_mem_req_valid),
    .io_mem_req_bits_addr(frontEnd_io_mem_req_bits_addr),
    .io_mem_resp_valid(frontEnd_io_mem_resp_valid),
    .io_mem_resp_bits_data(frontEnd_io_mem_resp_bits_data),
    .io_back_xcpt_valid(frontEnd_io_back_xcpt_valid),
    .io_back_xcpt_bits(frontEnd_io_back_xcpt_bits),
    .io_back_kill(frontEnd_io_back_kill),
    .io_back_fence(frontEnd_io_back_fence),
    .io_back_forward(frontEnd_io_back_forward),
    .io_back_ras_pop(frontEnd_io_back_ras_pop),
    .io_back_ras_push_valid(frontEnd_io_back_ras_push_valid),
    .io_back_ras_push_bits(frontEnd_io_back_ras_push_bits),
    .io_back_fb_pc(frontEnd_io_back_fb_pc),
    .io_back_fb_type(frontEnd_io_back_fb_type),
    .io_back_feedBack_valid(frontEnd_io_back_feedBack_valid),
    .io_back_feedBack_bits_redirect(frontEnd_io_back_feedBack_bits_redirect),
    .io_back_feedBack_bits_tgt(frontEnd_io_back_feedBack_bits_tgt),
    .io_back_inst_valid(frontEnd_io_back_inst_valid),
    .io_back_inst_bits(frontEnd_io_back_inst_bits),
    .io_back_pc(frontEnd_io_back_pc),
    .io_back_pred(frontEnd_io_back_pred)
  );
  BackEnd backEnd ( // @[Core.scala 31:24:@5624.4]
    .clock(backEnd_clock),
    .reset(backEnd_reset),
    .io_mem_req_valid(backEnd_io_mem_req_valid),
    .io_mem_req_bits_addr(backEnd_io_mem_req_bits_addr),
    .io_mem_req_bits_data(backEnd_io_mem_req_bits_data),
    .io_mem_req_bits_fcn(backEnd_io_mem_req_bits_fcn),
    .io_mem_req_bits_typ(backEnd_io_mem_req_bits_typ),
    .io_mem_resp_valid(backEnd_io_mem_resp_valid),
    .io_mem_resp_bits_data(backEnd_io_mem_resp_bits_data),
    .io_cyc(backEnd_io_cyc),
    .io_front_xcpt_valid(backEnd_io_front_xcpt_valid),
    .io_front_xcpt_bits(backEnd_io_front_xcpt_bits),
    .io_front_kill(backEnd_io_front_kill),
    .io_front_fence(backEnd_io_front_fence),
    .io_front_forward(backEnd_io_front_forward),
    .io_front_ras_pop(backEnd_io_front_ras_pop),
    .io_front_ras_push_valid(backEnd_io_front_ras_push_valid),
    .io_front_ras_push_bits(backEnd_io_front_ras_push_bits),
    .io_front_fb_pc(backEnd_io_front_fb_pc),
    .io_front_fb_type(backEnd_io_front_fb_type),
    .io_front_feedBack_valid(backEnd_io_front_feedBack_valid),
    .io_front_feedBack_bits_redirect(backEnd_io_front_feedBack_bits_redirect),
    .io_front_feedBack_bits_tgt(backEnd_io_front_feedBack_bits_tgt),
    .io_front_inst_valid(backEnd_io_front_inst_valid),
    .io_front_inst_bits(backEnd_io_front_inst_bits),
    .io_front_pc(backEnd_io_front_pc),
    .io_front_pred(backEnd_io_front_pred)
  );
  assign io_imem_req_valid = frontEnd_io_mem_req_valid; // @[Core.scala 32:20:@5633.4]
  assign io_imem_req_bits_addr = frontEnd_io_mem_req_bits_addr; // @[Core.scala 32:20:@5632.4]
  assign io_dmem_req_valid = backEnd_io_mem_req_valid; // @[Core.scala 33:20:@5641.4]
  assign io_dmem_req_bits_addr = backEnd_io_mem_req_bits_addr; // @[Core.scala 33:20:@5640.4]
  assign io_dmem_req_bits_data = backEnd_io_mem_req_bits_data; // @[Core.scala 33:20:@5639.4]
  assign io_dmem_req_bits_fcn = backEnd_io_mem_req_bits_fcn; // @[Core.scala 33:20:@5638.4]
  assign io_dmem_req_bits_typ = backEnd_io_mem_req_bits_typ; // @[Core.scala 33:20:@5637.4]
  assign frontEnd_clock = clock; // @[:@5622.4]
  assign frontEnd_reset = reset; // @[:@5623.4]
  assign frontEnd_io_cyc = backEnd_io_cyc; // @[Core.scala 35:20:@5660.4]
  assign frontEnd_io_mem_resp_valid = io_imem_resp_valid; // @[Core.scala 32:20:@5628.4]
  assign frontEnd_io_mem_resp_bits_data = io_imem_resp_bits_data; // @[Core.scala 32:20:@5627.4]
  assign frontEnd_io_back_xcpt_valid = backEnd_io_front_xcpt_valid; // @[Core.scala 34:20:@5659.4]
  assign frontEnd_io_back_xcpt_bits = backEnd_io_front_xcpt_bits; // @[Core.scala 34:20:@5658.4]
  assign frontEnd_io_back_kill = backEnd_io_front_kill; // @[Core.scala 34:20:@5657.4]
  assign frontEnd_io_back_fence = backEnd_io_front_fence; // @[Core.scala 34:20:@5656.4]
  assign frontEnd_io_back_forward = backEnd_io_front_forward; // @[Core.scala 34:20:@5655.4]
  assign frontEnd_io_back_ras_pop = backEnd_io_front_ras_pop; // @[Core.scala 34:20:@5654.4]
  assign frontEnd_io_back_ras_push_valid = backEnd_io_front_ras_push_valid; // @[Core.scala 34:20:@5653.4]
  assign frontEnd_io_back_ras_push_bits = backEnd_io_front_ras_push_bits; // @[Core.scala 34:20:@5652.4]
  assign frontEnd_io_back_fb_pc = backEnd_io_front_fb_pc; // @[Core.scala 34:20:@5651.4]
  assign frontEnd_io_back_fb_type = backEnd_io_front_fb_type; // @[Core.scala 34:20:@5650.4]
  assign frontEnd_io_back_feedBack_valid = backEnd_io_front_feedBack_valid; // @[Core.scala 34:20:@5649.4]
  assign frontEnd_io_back_feedBack_bits_redirect = backEnd_io_front_feedBack_bits_redirect; // @[Core.scala 34:20:@5648.4]
  assign frontEnd_io_back_feedBack_bits_tgt = backEnd_io_front_feedBack_bits_tgt; // @[Core.scala 34:20:@5647.4]
  assign backEnd_clock = clock; // @[:@5625.4]
  assign backEnd_reset = reset; // @[:@5626.4]
  assign backEnd_io_mem_resp_valid = io_dmem_resp_valid; // @[Core.scala 33:20:@5636.4]
  assign backEnd_io_mem_resp_bits_data = io_dmem_resp_bits_data; // @[Core.scala 33:20:@5635.4]
  assign backEnd_io_front_inst_valid = frontEnd_io_back_inst_valid; // @[Core.scala 34:20:@5646.4]
  assign backEnd_io_front_inst_bits = frontEnd_io_back_inst_bits; // @[Core.scala 34:20:@5645.4]
  assign backEnd_io_front_pc = frontEnd_io_back_pc; // @[Core.scala 34:20:@5644.4]
  assign backEnd_io_front_pred = frontEnd_io_back_pred; // @[Core.scala 34:20:@5643.4]
endmodule
